// Generator : SpinalHDL v1.4.1    git head : d1b4746673438bc5f242515335278fa39a666c38
// Component : FFT2d
// Git hash  : 5f24b07ffbfeb9934f5bea4487f4e9b5769de5ba



module FFT2d (
  input               io_line_in_valid,
  input      [17:0]   io_line_in_payload_0_real,
  input      [17:0]   io_line_in_payload_0_imag,
  input      [17:0]   io_line_in_payload_1_real,
  input      [17:0]   io_line_in_payload_1_imag,
  input      [17:0]   io_line_in_payload_2_real,
  input      [17:0]   io_line_in_payload_2_imag,
  input      [17:0]   io_line_in_payload_3_real,
  input      [17:0]   io_line_in_payload_3_imag,
  input      [17:0]   io_line_in_payload_4_real,
  input      [17:0]   io_line_in_payload_4_imag,
  input      [17:0]   io_line_in_payload_5_real,
  input      [17:0]   io_line_in_payload_5_imag,
  input      [17:0]   io_line_in_payload_6_real,
  input      [17:0]   io_line_in_payload_6_imag,
  input      [17:0]   io_line_in_payload_7_real,
  input      [17:0]   io_line_in_payload_7_imag,
  input      [17:0]   io_line_in_payload_8_real,
  input      [17:0]   io_line_in_payload_8_imag,
  input      [17:0]   io_line_in_payload_9_real,
  input      [17:0]   io_line_in_payload_9_imag,
  input      [17:0]   io_line_in_payload_10_real,
  input      [17:0]   io_line_in_payload_10_imag,
  input      [17:0]   io_line_in_payload_11_real,
  input      [17:0]   io_line_in_payload_11_imag,
  input      [17:0]   io_line_in_payload_12_real,
  input      [17:0]   io_line_in_payload_12_imag,
  input      [17:0]   io_line_in_payload_13_real,
  input      [17:0]   io_line_in_payload_13_imag,
  input      [17:0]   io_line_in_payload_14_real,
  input      [17:0]   io_line_in_payload_14_imag,
  input      [17:0]   io_line_in_payload_15_real,
  input      [17:0]   io_line_in_payload_15_imag,
  input      [17:0]   io_line_in_payload_16_real,
  input      [17:0]   io_line_in_payload_16_imag,
  input      [17:0]   io_line_in_payload_17_real,
  input      [17:0]   io_line_in_payload_17_imag,
  input      [17:0]   io_line_in_payload_18_real,
  input      [17:0]   io_line_in_payload_18_imag,
  input      [17:0]   io_line_in_payload_19_real,
  input      [17:0]   io_line_in_payload_19_imag,
  input      [17:0]   io_line_in_payload_20_real,
  input      [17:0]   io_line_in_payload_20_imag,
  input      [17:0]   io_line_in_payload_21_real,
  input      [17:0]   io_line_in_payload_21_imag,
  input      [17:0]   io_line_in_payload_22_real,
  input      [17:0]   io_line_in_payload_22_imag,
  input      [17:0]   io_line_in_payload_23_real,
  input      [17:0]   io_line_in_payload_23_imag,
  input      [17:0]   io_line_in_payload_24_real,
  input      [17:0]   io_line_in_payload_24_imag,
  input      [17:0]   io_line_in_payload_25_real,
  input      [17:0]   io_line_in_payload_25_imag,
  input      [17:0]   io_line_in_payload_26_real,
  input      [17:0]   io_line_in_payload_26_imag,
  input      [17:0]   io_line_in_payload_27_real,
  input      [17:0]   io_line_in_payload_27_imag,
  input      [17:0]   io_line_in_payload_28_real,
  input      [17:0]   io_line_in_payload_28_imag,
  input      [17:0]   io_line_in_payload_29_real,
  input      [17:0]   io_line_in_payload_29_imag,
  input      [17:0]   io_line_in_payload_30_real,
  input      [17:0]   io_line_in_payload_30_imag,
  input      [17:0]   io_line_in_payload_31_real,
  input      [17:0]   io_line_in_payload_31_imag,
  input      [17:0]   io_line_in_payload_32_real,
  input      [17:0]   io_line_in_payload_32_imag,
  input      [17:0]   io_line_in_payload_33_real,
  input      [17:0]   io_line_in_payload_33_imag,
  input      [17:0]   io_line_in_payload_34_real,
  input      [17:0]   io_line_in_payload_34_imag,
  input      [17:0]   io_line_in_payload_35_real,
  input      [17:0]   io_line_in_payload_35_imag,
  input      [17:0]   io_line_in_payload_36_real,
  input      [17:0]   io_line_in_payload_36_imag,
  input      [17:0]   io_line_in_payload_37_real,
  input      [17:0]   io_line_in_payload_37_imag,
  input      [17:0]   io_line_in_payload_38_real,
  input      [17:0]   io_line_in_payload_38_imag,
  input      [17:0]   io_line_in_payload_39_real,
  input      [17:0]   io_line_in_payload_39_imag,
  input      [17:0]   io_line_in_payload_40_real,
  input      [17:0]   io_line_in_payload_40_imag,
  input      [17:0]   io_line_in_payload_41_real,
  input      [17:0]   io_line_in_payload_41_imag,
  input      [17:0]   io_line_in_payload_42_real,
  input      [17:0]   io_line_in_payload_42_imag,
  input      [17:0]   io_line_in_payload_43_real,
  input      [17:0]   io_line_in_payload_43_imag,
  input      [17:0]   io_line_in_payload_44_real,
  input      [17:0]   io_line_in_payload_44_imag,
  input      [17:0]   io_line_in_payload_45_real,
  input      [17:0]   io_line_in_payload_45_imag,
  input      [17:0]   io_line_in_payload_46_real,
  input      [17:0]   io_line_in_payload_46_imag,
  input      [17:0]   io_line_in_payload_47_real,
  input      [17:0]   io_line_in_payload_47_imag,
  input      [17:0]   io_line_in_payload_48_real,
  input      [17:0]   io_line_in_payload_48_imag,
  input      [17:0]   io_line_in_payload_49_real,
  input      [17:0]   io_line_in_payload_49_imag,
  input      [17:0]   io_line_in_payload_50_real,
  input      [17:0]   io_line_in_payload_50_imag,
  input      [17:0]   io_line_in_payload_51_real,
  input      [17:0]   io_line_in_payload_51_imag,
  input      [17:0]   io_line_in_payload_52_real,
  input      [17:0]   io_line_in_payload_52_imag,
  input      [17:0]   io_line_in_payload_53_real,
  input      [17:0]   io_line_in_payload_53_imag,
  input      [17:0]   io_line_in_payload_54_real,
  input      [17:0]   io_line_in_payload_54_imag,
  input      [17:0]   io_line_in_payload_55_real,
  input      [17:0]   io_line_in_payload_55_imag,
  input      [17:0]   io_line_in_payload_56_real,
  input      [17:0]   io_line_in_payload_56_imag,
  input      [17:0]   io_line_in_payload_57_real,
  input      [17:0]   io_line_in_payload_57_imag,
  input      [17:0]   io_line_in_payload_58_real,
  input      [17:0]   io_line_in_payload_58_imag,
  input      [17:0]   io_line_in_payload_59_real,
  input      [17:0]   io_line_in_payload_59_imag,
  input      [17:0]   io_line_in_payload_60_real,
  input      [17:0]   io_line_in_payload_60_imag,
  input      [17:0]   io_line_in_payload_61_real,
  input      [17:0]   io_line_in_payload_61_imag,
  input      [17:0]   io_line_in_payload_62_real,
  input      [17:0]   io_line_in_payload_62_imag,
  input      [17:0]   io_line_in_payload_63_real,
  input      [17:0]   io_line_in_payload_63_imag,
  output              io_line_out_valid,
  output     [17:0]   io_line_out_payload_0_real,
  output     [17:0]   io_line_out_payload_0_imag,
  output     [17:0]   io_line_out_payload_1_real,
  output     [17:0]   io_line_out_payload_1_imag,
  output     [17:0]   io_line_out_payload_2_real,
  output     [17:0]   io_line_out_payload_2_imag,
  output     [17:0]   io_line_out_payload_3_real,
  output     [17:0]   io_line_out_payload_3_imag,
  output     [17:0]   io_line_out_payload_4_real,
  output     [17:0]   io_line_out_payload_4_imag,
  output     [17:0]   io_line_out_payload_5_real,
  output     [17:0]   io_line_out_payload_5_imag,
  output     [17:0]   io_line_out_payload_6_real,
  output     [17:0]   io_line_out_payload_6_imag,
  output     [17:0]   io_line_out_payload_7_real,
  output     [17:0]   io_line_out_payload_7_imag,
  output     [17:0]   io_line_out_payload_8_real,
  output     [17:0]   io_line_out_payload_8_imag,
  output     [17:0]   io_line_out_payload_9_real,
  output     [17:0]   io_line_out_payload_9_imag,
  output     [17:0]   io_line_out_payload_10_real,
  output     [17:0]   io_line_out_payload_10_imag,
  output     [17:0]   io_line_out_payload_11_real,
  output     [17:0]   io_line_out_payload_11_imag,
  output     [17:0]   io_line_out_payload_12_real,
  output     [17:0]   io_line_out_payload_12_imag,
  output     [17:0]   io_line_out_payload_13_real,
  output     [17:0]   io_line_out_payload_13_imag,
  output     [17:0]   io_line_out_payload_14_real,
  output     [17:0]   io_line_out_payload_14_imag,
  output     [17:0]   io_line_out_payload_15_real,
  output     [17:0]   io_line_out_payload_15_imag,
  output     [17:0]   io_line_out_payload_16_real,
  output     [17:0]   io_line_out_payload_16_imag,
  output     [17:0]   io_line_out_payload_17_real,
  output     [17:0]   io_line_out_payload_17_imag,
  output     [17:0]   io_line_out_payload_18_real,
  output     [17:0]   io_line_out_payload_18_imag,
  output     [17:0]   io_line_out_payload_19_real,
  output     [17:0]   io_line_out_payload_19_imag,
  output     [17:0]   io_line_out_payload_20_real,
  output     [17:0]   io_line_out_payload_20_imag,
  output     [17:0]   io_line_out_payload_21_real,
  output     [17:0]   io_line_out_payload_21_imag,
  output     [17:0]   io_line_out_payload_22_real,
  output     [17:0]   io_line_out_payload_22_imag,
  output     [17:0]   io_line_out_payload_23_real,
  output     [17:0]   io_line_out_payload_23_imag,
  output     [17:0]   io_line_out_payload_24_real,
  output     [17:0]   io_line_out_payload_24_imag,
  output     [17:0]   io_line_out_payload_25_real,
  output     [17:0]   io_line_out_payload_25_imag,
  output     [17:0]   io_line_out_payload_26_real,
  output     [17:0]   io_line_out_payload_26_imag,
  output     [17:0]   io_line_out_payload_27_real,
  output     [17:0]   io_line_out_payload_27_imag,
  output     [17:0]   io_line_out_payload_28_real,
  output     [17:0]   io_line_out_payload_28_imag,
  output     [17:0]   io_line_out_payload_29_real,
  output     [17:0]   io_line_out_payload_29_imag,
  output     [17:0]   io_line_out_payload_30_real,
  output     [17:0]   io_line_out_payload_30_imag,
  output     [17:0]   io_line_out_payload_31_real,
  output     [17:0]   io_line_out_payload_31_imag,
  output     [17:0]   io_line_out_payload_32_real,
  output     [17:0]   io_line_out_payload_32_imag,
  output     [17:0]   io_line_out_payload_33_real,
  output     [17:0]   io_line_out_payload_33_imag,
  output     [17:0]   io_line_out_payload_34_real,
  output     [17:0]   io_line_out_payload_34_imag,
  output     [17:0]   io_line_out_payload_35_real,
  output     [17:0]   io_line_out_payload_35_imag,
  output     [17:0]   io_line_out_payload_36_real,
  output     [17:0]   io_line_out_payload_36_imag,
  output     [17:0]   io_line_out_payload_37_real,
  output     [17:0]   io_line_out_payload_37_imag,
  output     [17:0]   io_line_out_payload_38_real,
  output     [17:0]   io_line_out_payload_38_imag,
  output     [17:0]   io_line_out_payload_39_real,
  output     [17:0]   io_line_out_payload_39_imag,
  output     [17:0]   io_line_out_payload_40_real,
  output     [17:0]   io_line_out_payload_40_imag,
  output     [17:0]   io_line_out_payload_41_real,
  output     [17:0]   io_line_out_payload_41_imag,
  output     [17:0]   io_line_out_payload_42_real,
  output     [17:0]   io_line_out_payload_42_imag,
  output     [17:0]   io_line_out_payload_43_real,
  output     [17:0]   io_line_out_payload_43_imag,
  output     [17:0]   io_line_out_payload_44_real,
  output     [17:0]   io_line_out_payload_44_imag,
  output     [17:0]   io_line_out_payload_45_real,
  output     [17:0]   io_line_out_payload_45_imag,
  output     [17:0]   io_line_out_payload_46_real,
  output     [17:0]   io_line_out_payload_46_imag,
  output     [17:0]   io_line_out_payload_47_real,
  output     [17:0]   io_line_out_payload_47_imag,
  output     [17:0]   io_line_out_payload_48_real,
  output     [17:0]   io_line_out_payload_48_imag,
  output     [17:0]   io_line_out_payload_49_real,
  output     [17:0]   io_line_out_payload_49_imag,
  output     [17:0]   io_line_out_payload_50_real,
  output     [17:0]   io_line_out_payload_50_imag,
  output     [17:0]   io_line_out_payload_51_real,
  output     [17:0]   io_line_out_payload_51_imag,
  output     [17:0]   io_line_out_payload_52_real,
  output     [17:0]   io_line_out_payload_52_imag,
  output     [17:0]   io_line_out_payload_53_real,
  output     [17:0]   io_line_out_payload_53_imag,
  output     [17:0]   io_line_out_payload_54_real,
  output     [17:0]   io_line_out_payload_54_imag,
  output     [17:0]   io_line_out_payload_55_real,
  output     [17:0]   io_line_out_payload_55_imag,
  output     [17:0]   io_line_out_payload_56_real,
  output     [17:0]   io_line_out_payload_56_imag,
  output     [17:0]   io_line_out_payload_57_real,
  output     [17:0]   io_line_out_payload_57_imag,
  output     [17:0]   io_line_out_payload_58_real,
  output     [17:0]   io_line_out_payload_58_imag,
  output     [17:0]   io_line_out_payload_59_real,
  output     [17:0]   io_line_out_payload_59_imag,
  output     [17:0]   io_line_out_payload_60_real,
  output     [17:0]   io_line_out_payload_60_imag,
  output     [17:0]   io_line_out_payload_61_real,
  output     [17:0]   io_line_out_payload_61_imag,
  output     [17:0]   io_line_out_payload_62_real,
  output     [17:0]   io_line_out_payload_62_imag,
  output     [17:0]   io_line_out_payload_63_real,
  output     [17:0]   io_line_out_payload_63_imag,
  input               clk,
  input               reset
);
  reg        [17:0]   _zz_194;
  reg        [17:0]   _zz_195;
  reg        [17:0]   _zz_196;
  reg        [17:0]   _zz_197;
  reg        [17:0]   _zz_198;
  reg        [17:0]   _zz_199;
  reg        [17:0]   _zz_200;
  reg        [17:0]   _zz_201;
  reg        [17:0]   _zz_202;
  reg        [17:0]   _zz_203;
  reg        [17:0]   _zz_204;
  reg        [17:0]   _zz_205;
  reg        [17:0]   _zz_206;
  reg        [17:0]   _zz_207;
  reg        [17:0]   _zz_208;
  reg        [17:0]   _zz_209;
  reg        [17:0]   _zz_210;
  reg        [17:0]   _zz_211;
  reg        [17:0]   _zz_212;
  reg        [17:0]   _zz_213;
  reg        [17:0]   _zz_214;
  reg        [17:0]   _zz_215;
  reg        [17:0]   _zz_216;
  reg        [17:0]   _zz_217;
  reg        [17:0]   _zz_218;
  reg        [17:0]   _zz_219;
  reg        [17:0]   _zz_220;
  reg        [17:0]   _zz_221;
  reg        [17:0]   _zz_222;
  reg        [17:0]   _zz_223;
  reg        [17:0]   _zz_224;
  reg        [17:0]   _zz_225;
  reg        [17:0]   _zz_226;
  reg        [17:0]   _zz_227;
  reg        [17:0]   _zz_228;
  reg        [17:0]   _zz_229;
  reg        [17:0]   _zz_230;
  reg        [17:0]   _zz_231;
  reg        [17:0]   _zz_232;
  reg        [17:0]   _zz_233;
  reg        [17:0]   _zz_234;
  reg        [17:0]   _zz_235;
  reg        [17:0]   _zz_236;
  reg        [17:0]   _zz_237;
  reg        [17:0]   _zz_238;
  reg        [17:0]   _zz_239;
  reg        [17:0]   _zz_240;
  reg        [17:0]   _zz_241;
  reg        [17:0]   _zz_242;
  reg        [17:0]   _zz_243;
  reg        [17:0]   _zz_244;
  reg        [17:0]   _zz_245;
  reg        [17:0]   _zz_246;
  reg        [17:0]   _zz_247;
  reg        [17:0]   _zz_248;
  reg        [17:0]   _zz_249;
  reg        [17:0]   _zz_250;
  reg        [17:0]   _zz_251;
  reg        [17:0]   _zz_252;
  reg        [17:0]   _zz_253;
  reg        [17:0]   _zz_254;
  reg        [17:0]   _zz_255;
  reg        [17:0]   _zz_256;
  reg        [17:0]   _zz_257;
  reg        [17:0]   _zz_258;
  reg        [17:0]   _zz_259;
  reg        [17:0]   _zz_260;
  reg        [17:0]   _zz_261;
  reg        [17:0]   _zz_262;
  reg        [17:0]   _zz_263;
  reg        [17:0]   _zz_264;
  reg        [17:0]   _zz_265;
  reg        [17:0]   _zz_266;
  reg        [17:0]   _zz_267;
  reg        [17:0]   _zz_268;
  reg        [17:0]   _zz_269;
  reg        [17:0]   _zz_270;
  reg        [17:0]   _zz_271;
  reg        [17:0]   _zz_272;
  reg        [17:0]   _zz_273;
  reg        [17:0]   _zz_274;
  reg        [17:0]   _zz_275;
  reg        [17:0]   _zz_276;
  reg        [17:0]   _zz_277;
  reg        [17:0]   _zz_278;
  reg        [17:0]   _zz_279;
  reg        [17:0]   _zz_280;
  reg        [17:0]   _zz_281;
  reg        [17:0]   _zz_282;
  reg        [17:0]   _zz_283;
  reg        [17:0]   _zz_284;
  reg        [17:0]   _zz_285;
  reg        [17:0]   _zz_286;
  reg        [17:0]   _zz_287;
  reg        [17:0]   _zz_288;
  reg        [17:0]   _zz_289;
  reg        [17:0]   _zz_290;
  reg        [17:0]   _zz_291;
  reg        [17:0]   _zz_292;
  reg        [17:0]   _zz_293;
  reg        [17:0]   _zz_294;
  reg        [17:0]   _zz_295;
  reg        [17:0]   _zz_296;
  reg        [17:0]   _zz_297;
  reg        [17:0]   _zz_298;
  reg        [17:0]   _zz_299;
  reg        [17:0]   _zz_300;
  reg        [17:0]   _zz_301;
  reg        [17:0]   _zz_302;
  reg        [17:0]   _zz_303;
  reg        [17:0]   _zz_304;
  reg        [17:0]   _zz_305;
  reg        [17:0]   _zz_306;
  reg        [17:0]   _zz_307;
  reg        [17:0]   _zz_308;
  reg        [17:0]   _zz_309;
  reg        [17:0]   _zz_310;
  reg        [17:0]   _zz_311;
  reg        [17:0]   _zz_312;
  reg        [17:0]   _zz_313;
  reg        [17:0]   _zz_314;
  reg        [17:0]   _zz_315;
  reg        [17:0]   _zz_316;
  reg        [17:0]   _zz_317;
  reg        [17:0]   _zz_318;
  reg        [17:0]   _zz_319;
  reg        [17:0]   _zz_320;
  reg        [17:0]   _zz_321;
  wire                myFFT_2_fft_row_valid;
  wire       [17:0]   myFFT_2_fft_row_payload_0_real;
  wire       [17:0]   myFFT_2_fft_row_payload_0_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_1_real;
  wire       [17:0]   myFFT_2_fft_row_payload_1_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_2_real;
  wire       [17:0]   myFFT_2_fft_row_payload_2_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_3_real;
  wire       [17:0]   myFFT_2_fft_row_payload_3_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_4_real;
  wire       [17:0]   myFFT_2_fft_row_payload_4_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_5_real;
  wire       [17:0]   myFFT_2_fft_row_payload_5_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_6_real;
  wire       [17:0]   myFFT_2_fft_row_payload_6_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_7_real;
  wire       [17:0]   myFFT_2_fft_row_payload_7_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_8_real;
  wire       [17:0]   myFFT_2_fft_row_payload_8_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_9_real;
  wire       [17:0]   myFFT_2_fft_row_payload_9_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_10_real;
  wire       [17:0]   myFFT_2_fft_row_payload_10_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_11_real;
  wire       [17:0]   myFFT_2_fft_row_payload_11_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_12_real;
  wire       [17:0]   myFFT_2_fft_row_payload_12_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_13_real;
  wire       [17:0]   myFFT_2_fft_row_payload_13_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_14_real;
  wire       [17:0]   myFFT_2_fft_row_payload_14_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_15_real;
  wire       [17:0]   myFFT_2_fft_row_payload_15_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_16_real;
  wire       [17:0]   myFFT_2_fft_row_payload_16_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_17_real;
  wire       [17:0]   myFFT_2_fft_row_payload_17_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_18_real;
  wire       [17:0]   myFFT_2_fft_row_payload_18_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_19_real;
  wire       [17:0]   myFFT_2_fft_row_payload_19_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_20_real;
  wire       [17:0]   myFFT_2_fft_row_payload_20_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_21_real;
  wire       [17:0]   myFFT_2_fft_row_payload_21_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_22_real;
  wire       [17:0]   myFFT_2_fft_row_payload_22_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_23_real;
  wire       [17:0]   myFFT_2_fft_row_payload_23_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_24_real;
  wire       [17:0]   myFFT_2_fft_row_payload_24_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_25_real;
  wire       [17:0]   myFFT_2_fft_row_payload_25_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_26_real;
  wire       [17:0]   myFFT_2_fft_row_payload_26_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_27_real;
  wire       [17:0]   myFFT_2_fft_row_payload_27_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_28_real;
  wire       [17:0]   myFFT_2_fft_row_payload_28_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_29_real;
  wire       [17:0]   myFFT_2_fft_row_payload_29_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_30_real;
  wire       [17:0]   myFFT_2_fft_row_payload_30_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_31_real;
  wire       [17:0]   myFFT_2_fft_row_payload_31_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_32_real;
  wire       [17:0]   myFFT_2_fft_row_payload_32_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_33_real;
  wire       [17:0]   myFFT_2_fft_row_payload_33_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_34_real;
  wire       [17:0]   myFFT_2_fft_row_payload_34_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_35_real;
  wire       [17:0]   myFFT_2_fft_row_payload_35_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_36_real;
  wire       [17:0]   myFFT_2_fft_row_payload_36_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_37_real;
  wire       [17:0]   myFFT_2_fft_row_payload_37_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_38_real;
  wire       [17:0]   myFFT_2_fft_row_payload_38_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_39_real;
  wire       [17:0]   myFFT_2_fft_row_payload_39_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_40_real;
  wire       [17:0]   myFFT_2_fft_row_payload_40_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_41_real;
  wire       [17:0]   myFFT_2_fft_row_payload_41_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_42_real;
  wire       [17:0]   myFFT_2_fft_row_payload_42_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_43_real;
  wire       [17:0]   myFFT_2_fft_row_payload_43_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_44_real;
  wire       [17:0]   myFFT_2_fft_row_payload_44_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_45_real;
  wire       [17:0]   myFFT_2_fft_row_payload_45_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_46_real;
  wire       [17:0]   myFFT_2_fft_row_payload_46_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_47_real;
  wire       [17:0]   myFFT_2_fft_row_payload_47_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_48_real;
  wire       [17:0]   myFFT_2_fft_row_payload_48_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_49_real;
  wire       [17:0]   myFFT_2_fft_row_payload_49_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_50_real;
  wire       [17:0]   myFFT_2_fft_row_payload_50_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_51_real;
  wire       [17:0]   myFFT_2_fft_row_payload_51_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_52_real;
  wire       [17:0]   myFFT_2_fft_row_payload_52_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_53_real;
  wire       [17:0]   myFFT_2_fft_row_payload_53_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_54_real;
  wire       [17:0]   myFFT_2_fft_row_payload_54_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_55_real;
  wire       [17:0]   myFFT_2_fft_row_payload_55_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_56_real;
  wire       [17:0]   myFFT_2_fft_row_payload_56_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_57_real;
  wire       [17:0]   myFFT_2_fft_row_payload_57_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_58_real;
  wire       [17:0]   myFFT_2_fft_row_payload_58_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_59_real;
  wire       [17:0]   myFFT_2_fft_row_payload_59_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_60_real;
  wire       [17:0]   myFFT_2_fft_row_payload_60_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_61_real;
  wire       [17:0]   myFFT_2_fft_row_payload_61_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_62_real;
  wire       [17:0]   myFFT_2_fft_row_payload_62_imag;
  wire       [17:0]   myFFT_2_fft_row_payload_63_real;
  wire       [17:0]   myFFT_2_fft_row_payload_63_imag;
  wire                myFFT_3_fft_col_out_valid;
  wire       [17:0]   myFFT_3_fft_col_out_payload_0_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_0_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_1_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_1_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_2_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_2_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_3_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_3_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_4_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_4_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_5_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_5_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_6_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_6_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_7_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_7_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_8_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_8_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_9_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_9_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_10_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_10_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_11_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_11_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_12_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_12_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_13_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_13_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_14_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_14_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_15_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_15_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_16_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_16_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_17_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_17_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_18_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_18_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_19_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_19_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_20_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_20_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_21_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_21_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_22_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_22_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_23_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_23_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_24_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_24_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_25_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_25_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_26_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_26_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_27_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_27_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_28_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_28_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_29_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_29_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_30_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_30_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_31_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_31_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_32_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_32_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_33_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_33_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_34_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_34_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_35_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_35_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_36_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_36_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_37_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_37_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_38_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_38_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_39_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_39_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_40_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_40_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_41_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_41_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_42_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_42_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_43_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_43_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_44_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_44_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_45_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_45_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_46_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_46_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_47_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_47_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_48_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_48_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_49_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_49_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_50_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_50_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_51_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_51_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_52_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_52_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_53_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_53_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_54_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_54_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_55_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_55_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_56_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_56_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_57_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_57_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_58_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_58_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_59_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_59_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_60_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_60_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_61_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_61_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_62_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_62_imag;
  wire       [17:0]   myFFT_3_fft_col_out_payload_63_real;
  wire       [17:0]   myFFT_3_fft_col_out_payload_63_imag;
  wire       [0:0]    _zz_322;
  wire       [5:0]    _zz_323;
  wire       [0:0]    _zz_324;
  wire       [5:0]    _zz_325;
  reg        [17:0]   img_reg_array_0_0_real;
  reg        [17:0]   img_reg_array_0_0_imag;
  reg        [17:0]   img_reg_array_0_1_real;
  reg        [17:0]   img_reg_array_0_1_imag;
  reg        [17:0]   img_reg_array_0_2_real;
  reg        [17:0]   img_reg_array_0_2_imag;
  reg        [17:0]   img_reg_array_0_3_real;
  reg        [17:0]   img_reg_array_0_3_imag;
  reg        [17:0]   img_reg_array_0_4_real;
  reg        [17:0]   img_reg_array_0_4_imag;
  reg        [17:0]   img_reg_array_0_5_real;
  reg        [17:0]   img_reg_array_0_5_imag;
  reg        [17:0]   img_reg_array_0_6_real;
  reg        [17:0]   img_reg_array_0_6_imag;
  reg        [17:0]   img_reg_array_0_7_real;
  reg        [17:0]   img_reg_array_0_7_imag;
  reg        [17:0]   img_reg_array_0_8_real;
  reg        [17:0]   img_reg_array_0_8_imag;
  reg        [17:0]   img_reg_array_0_9_real;
  reg        [17:0]   img_reg_array_0_9_imag;
  reg        [17:0]   img_reg_array_0_10_real;
  reg        [17:0]   img_reg_array_0_10_imag;
  reg        [17:0]   img_reg_array_0_11_real;
  reg        [17:0]   img_reg_array_0_11_imag;
  reg        [17:0]   img_reg_array_0_12_real;
  reg        [17:0]   img_reg_array_0_12_imag;
  reg        [17:0]   img_reg_array_0_13_real;
  reg        [17:0]   img_reg_array_0_13_imag;
  reg        [17:0]   img_reg_array_0_14_real;
  reg        [17:0]   img_reg_array_0_14_imag;
  reg        [17:0]   img_reg_array_0_15_real;
  reg        [17:0]   img_reg_array_0_15_imag;
  reg        [17:0]   img_reg_array_0_16_real;
  reg        [17:0]   img_reg_array_0_16_imag;
  reg        [17:0]   img_reg_array_0_17_real;
  reg        [17:0]   img_reg_array_0_17_imag;
  reg        [17:0]   img_reg_array_0_18_real;
  reg        [17:0]   img_reg_array_0_18_imag;
  reg        [17:0]   img_reg_array_0_19_real;
  reg        [17:0]   img_reg_array_0_19_imag;
  reg        [17:0]   img_reg_array_0_20_real;
  reg        [17:0]   img_reg_array_0_20_imag;
  reg        [17:0]   img_reg_array_0_21_real;
  reg        [17:0]   img_reg_array_0_21_imag;
  reg        [17:0]   img_reg_array_0_22_real;
  reg        [17:0]   img_reg_array_0_22_imag;
  reg        [17:0]   img_reg_array_0_23_real;
  reg        [17:0]   img_reg_array_0_23_imag;
  reg        [17:0]   img_reg_array_0_24_real;
  reg        [17:0]   img_reg_array_0_24_imag;
  reg        [17:0]   img_reg_array_0_25_real;
  reg        [17:0]   img_reg_array_0_25_imag;
  reg        [17:0]   img_reg_array_0_26_real;
  reg        [17:0]   img_reg_array_0_26_imag;
  reg        [17:0]   img_reg_array_0_27_real;
  reg        [17:0]   img_reg_array_0_27_imag;
  reg        [17:0]   img_reg_array_0_28_real;
  reg        [17:0]   img_reg_array_0_28_imag;
  reg        [17:0]   img_reg_array_0_29_real;
  reg        [17:0]   img_reg_array_0_29_imag;
  reg        [17:0]   img_reg_array_0_30_real;
  reg        [17:0]   img_reg_array_0_30_imag;
  reg        [17:0]   img_reg_array_0_31_real;
  reg        [17:0]   img_reg_array_0_31_imag;
  reg        [17:0]   img_reg_array_0_32_real;
  reg        [17:0]   img_reg_array_0_32_imag;
  reg        [17:0]   img_reg_array_0_33_real;
  reg        [17:0]   img_reg_array_0_33_imag;
  reg        [17:0]   img_reg_array_0_34_real;
  reg        [17:0]   img_reg_array_0_34_imag;
  reg        [17:0]   img_reg_array_0_35_real;
  reg        [17:0]   img_reg_array_0_35_imag;
  reg        [17:0]   img_reg_array_0_36_real;
  reg        [17:0]   img_reg_array_0_36_imag;
  reg        [17:0]   img_reg_array_0_37_real;
  reg        [17:0]   img_reg_array_0_37_imag;
  reg        [17:0]   img_reg_array_0_38_real;
  reg        [17:0]   img_reg_array_0_38_imag;
  reg        [17:0]   img_reg_array_0_39_real;
  reg        [17:0]   img_reg_array_0_39_imag;
  reg        [17:0]   img_reg_array_0_40_real;
  reg        [17:0]   img_reg_array_0_40_imag;
  reg        [17:0]   img_reg_array_0_41_real;
  reg        [17:0]   img_reg_array_0_41_imag;
  reg        [17:0]   img_reg_array_0_42_real;
  reg        [17:0]   img_reg_array_0_42_imag;
  reg        [17:0]   img_reg_array_0_43_real;
  reg        [17:0]   img_reg_array_0_43_imag;
  reg        [17:0]   img_reg_array_0_44_real;
  reg        [17:0]   img_reg_array_0_44_imag;
  reg        [17:0]   img_reg_array_0_45_real;
  reg        [17:0]   img_reg_array_0_45_imag;
  reg        [17:0]   img_reg_array_0_46_real;
  reg        [17:0]   img_reg_array_0_46_imag;
  reg        [17:0]   img_reg_array_0_47_real;
  reg        [17:0]   img_reg_array_0_47_imag;
  reg        [17:0]   img_reg_array_0_48_real;
  reg        [17:0]   img_reg_array_0_48_imag;
  reg        [17:0]   img_reg_array_0_49_real;
  reg        [17:0]   img_reg_array_0_49_imag;
  reg        [17:0]   img_reg_array_0_50_real;
  reg        [17:0]   img_reg_array_0_50_imag;
  reg        [17:0]   img_reg_array_0_51_real;
  reg        [17:0]   img_reg_array_0_51_imag;
  reg        [17:0]   img_reg_array_0_52_real;
  reg        [17:0]   img_reg_array_0_52_imag;
  reg        [17:0]   img_reg_array_0_53_real;
  reg        [17:0]   img_reg_array_0_53_imag;
  reg        [17:0]   img_reg_array_0_54_real;
  reg        [17:0]   img_reg_array_0_54_imag;
  reg        [17:0]   img_reg_array_0_55_real;
  reg        [17:0]   img_reg_array_0_55_imag;
  reg        [17:0]   img_reg_array_0_56_real;
  reg        [17:0]   img_reg_array_0_56_imag;
  reg        [17:0]   img_reg_array_0_57_real;
  reg        [17:0]   img_reg_array_0_57_imag;
  reg        [17:0]   img_reg_array_0_58_real;
  reg        [17:0]   img_reg_array_0_58_imag;
  reg        [17:0]   img_reg_array_0_59_real;
  reg        [17:0]   img_reg_array_0_59_imag;
  reg        [17:0]   img_reg_array_0_60_real;
  reg        [17:0]   img_reg_array_0_60_imag;
  reg        [17:0]   img_reg_array_0_61_real;
  reg        [17:0]   img_reg_array_0_61_imag;
  reg        [17:0]   img_reg_array_0_62_real;
  reg        [17:0]   img_reg_array_0_62_imag;
  reg        [17:0]   img_reg_array_0_63_real;
  reg        [17:0]   img_reg_array_0_63_imag;
  reg        [17:0]   img_reg_array_1_0_real;
  reg        [17:0]   img_reg_array_1_0_imag;
  reg        [17:0]   img_reg_array_1_1_real;
  reg        [17:0]   img_reg_array_1_1_imag;
  reg        [17:0]   img_reg_array_1_2_real;
  reg        [17:0]   img_reg_array_1_2_imag;
  reg        [17:0]   img_reg_array_1_3_real;
  reg        [17:0]   img_reg_array_1_3_imag;
  reg        [17:0]   img_reg_array_1_4_real;
  reg        [17:0]   img_reg_array_1_4_imag;
  reg        [17:0]   img_reg_array_1_5_real;
  reg        [17:0]   img_reg_array_1_5_imag;
  reg        [17:0]   img_reg_array_1_6_real;
  reg        [17:0]   img_reg_array_1_6_imag;
  reg        [17:0]   img_reg_array_1_7_real;
  reg        [17:0]   img_reg_array_1_7_imag;
  reg        [17:0]   img_reg_array_1_8_real;
  reg        [17:0]   img_reg_array_1_8_imag;
  reg        [17:0]   img_reg_array_1_9_real;
  reg        [17:0]   img_reg_array_1_9_imag;
  reg        [17:0]   img_reg_array_1_10_real;
  reg        [17:0]   img_reg_array_1_10_imag;
  reg        [17:0]   img_reg_array_1_11_real;
  reg        [17:0]   img_reg_array_1_11_imag;
  reg        [17:0]   img_reg_array_1_12_real;
  reg        [17:0]   img_reg_array_1_12_imag;
  reg        [17:0]   img_reg_array_1_13_real;
  reg        [17:0]   img_reg_array_1_13_imag;
  reg        [17:0]   img_reg_array_1_14_real;
  reg        [17:0]   img_reg_array_1_14_imag;
  reg        [17:0]   img_reg_array_1_15_real;
  reg        [17:0]   img_reg_array_1_15_imag;
  reg        [17:0]   img_reg_array_1_16_real;
  reg        [17:0]   img_reg_array_1_16_imag;
  reg        [17:0]   img_reg_array_1_17_real;
  reg        [17:0]   img_reg_array_1_17_imag;
  reg        [17:0]   img_reg_array_1_18_real;
  reg        [17:0]   img_reg_array_1_18_imag;
  reg        [17:0]   img_reg_array_1_19_real;
  reg        [17:0]   img_reg_array_1_19_imag;
  reg        [17:0]   img_reg_array_1_20_real;
  reg        [17:0]   img_reg_array_1_20_imag;
  reg        [17:0]   img_reg_array_1_21_real;
  reg        [17:0]   img_reg_array_1_21_imag;
  reg        [17:0]   img_reg_array_1_22_real;
  reg        [17:0]   img_reg_array_1_22_imag;
  reg        [17:0]   img_reg_array_1_23_real;
  reg        [17:0]   img_reg_array_1_23_imag;
  reg        [17:0]   img_reg_array_1_24_real;
  reg        [17:0]   img_reg_array_1_24_imag;
  reg        [17:0]   img_reg_array_1_25_real;
  reg        [17:0]   img_reg_array_1_25_imag;
  reg        [17:0]   img_reg_array_1_26_real;
  reg        [17:0]   img_reg_array_1_26_imag;
  reg        [17:0]   img_reg_array_1_27_real;
  reg        [17:0]   img_reg_array_1_27_imag;
  reg        [17:0]   img_reg_array_1_28_real;
  reg        [17:0]   img_reg_array_1_28_imag;
  reg        [17:0]   img_reg_array_1_29_real;
  reg        [17:0]   img_reg_array_1_29_imag;
  reg        [17:0]   img_reg_array_1_30_real;
  reg        [17:0]   img_reg_array_1_30_imag;
  reg        [17:0]   img_reg_array_1_31_real;
  reg        [17:0]   img_reg_array_1_31_imag;
  reg        [17:0]   img_reg_array_1_32_real;
  reg        [17:0]   img_reg_array_1_32_imag;
  reg        [17:0]   img_reg_array_1_33_real;
  reg        [17:0]   img_reg_array_1_33_imag;
  reg        [17:0]   img_reg_array_1_34_real;
  reg        [17:0]   img_reg_array_1_34_imag;
  reg        [17:0]   img_reg_array_1_35_real;
  reg        [17:0]   img_reg_array_1_35_imag;
  reg        [17:0]   img_reg_array_1_36_real;
  reg        [17:0]   img_reg_array_1_36_imag;
  reg        [17:0]   img_reg_array_1_37_real;
  reg        [17:0]   img_reg_array_1_37_imag;
  reg        [17:0]   img_reg_array_1_38_real;
  reg        [17:0]   img_reg_array_1_38_imag;
  reg        [17:0]   img_reg_array_1_39_real;
  reg        [17:0]   img_reg_array_1_39_imag;
  reg        [17:0]   img_reg_array_1_40_real;
  reg        [17:0]   img_reg_array_1_40_imag;
  reg        [17:0]   img_reg_array_1_41_real;
  reg        [17:0]   img_reg_array_1_41_imag;
  reg        [17:0]   img_reg_array_1_42_real;
  reg        [17:0]   img_reg_array_1_42_imag;
  reg        [17:0]   img_reg_array_1_43_real;
  reg        [17:0]   img_reg_array_1_43_imag;
  reg        [17:0]   img_reg_array_1_44_real;
  reg        [17:0]   img_reg_array_1_44_imag;
  reg        [17:0]   img_reg_array_1_45_real;
  reg        [17:0]   img_reg_array_1_45_imag;
  reg        [17:0]   img_reg_array_1_46_real;
  reg        [17:0]   img_reg_array_1_46_imag;
  reg        [17:0]   img_reg_array_1_47_real;
  reg        [17:0]   img_reg_array_1_47_imag;
  reg        [17:0]   img_reg_array_1_48_real;
  reg        [17:0]   img_reg_array_1_48_imag;
  reg        [17:0]   img_reg_array_1_49_real;
  reg        [17:0]   img_reg_array_1_49_imag;
  reg        [17:0]   img_reg_array_1_50_real;
  reg        [17:0]   img_reg_array_1_50_imag;
  reg        [17:0]   img_reg_array_1_51_real;
  reg        [17:0]   img_reg_array_1_51_imag;
  reg        [17:0]   img_reg_array_1_52_real;
  reg        [17:0]   img_reg_array_1_52_imag;
  reg        [17:0]   img_reg_array_1_53_real;
  reg        [17:0]   img_reg_array_1_53_imag;
  reg        [17:0]   img_reg_array_1_54_real;
  reg        [17:0]   img_reg_array_1_54_imag;
  reg        [17:0]   img_reg_array_1_55_real;
  reg        [17:0]   img_reg_array_1_55_imag;
  reg        [17:0]   img_reg_array_1_56_real;
  reg        [17:0]   img_reg_array_1_56_imag;
  reg        [17:0]   img_reg_array_1_57_real;
  reg        [17:0]   img_reg_array_1_57_imag;
  reg        [17:0]   img_reg_array_1_58_real;
  reg        [17:0]   img_reg_array_1_58_imag;
  reg        [17:0]   img_reg_array_1_59_real;
  reg        [17:0]   img_reg_array_1_59_imag;
  reg        [17:0]   img_reg_array_1_60_real;
  reg        [17:0]   img_reg_array_1_60_imag;
  reg        [17:0]   img_reg_array_1_61_real;
  reg        [17:0]   img_reg_array_1_61_imag;
  reg        [17:0]   img_reg_array_1_62_real;
  reg        [17:0]   img_reg_array_1_62_imag;
  reg        [17:0]   img_reg_array_1_63_real;
  reg        [17:0]   img_reg_array_1_63_imag;
  reg        [17:0]   img_reg_array_2_0_real;
  reg        [17:0]   img_reg_array_2_0_imag;
  reg        [17:0]   img_reg_array_2_1_real;
  reg        [17:0]   img_reg_array_2_1_imag;
  reg        [17:0]   img_reg_array_2_2_real;
  reg        [17:0]   img_reg_array_2_2_imag;
  reg        [17:0]   img_reg_array_2_3_real;
  reg        [17:0]   img_reg_array_2_3_imag;
  reg        [17:0]   img_reg_array_2_4_real;
  reg        [17:0]   img_reg_array_2_4_imag;
  reg        [17:0]   img_reg_array_2_5_real;
  reg        [17:0]   img_reg_array_2_5_imag;
  reg        [17:0]   img_reg_array_2_6_real;
  reg        [17:0]   img_reg_array_2_6_imag;
  reg        [17:0]   img_reg_array_2_7_real;
  reg        [17:0]   img_reg_array_2_7_imag;
  reg        [17:0]   img_reg_array_2_8_real;
  reg        [17:0]   img_reg_array_2_8_imag;
  reg        [17:0]   img_reg_array_2_9_real;
  reg        [17:0]   img_reg_array_2_9_imag;
  reg        [17:0]   img_reg_array_2_10_real;
  reg        [17:0]   img_reg_array_2_10_imag;
  reg        [17:0]   img_reg_array_2_11_real;
  reg        [17:0]   img_reg_array_2_11_imag;
  reg        [17:0]   img_reg_array_2_12_real;
  reg        [17:0]   img_reg_array_2_12_imag;
  reg        [17:0]   img_reg_array_2_13_real;
  reg        [17:0]   img_reg_array_2_13_imag;
  reg        [17:0]   img_reg_array_2_14_real;
  reg        [17:0]   img_reg_array_2_14_imag;
  reg        [17:0]   img_reg_array_2_15_real;
  reg        [17:0]   img_reg_array_2_15_imag;
  reg        [17:0]   img_reg_array_2_16_real;
  reg        [17:0]   img_reg_array_2_16_imag;
  reg        [17:0]   img_reg_array_2_17_real;
  reg        [17:0]   img_reg_array_2_17_imag;
  reg        [17:0]   img_reg_array_2_18_real;
  reg        [17:0]   img_reg_array_2_18_imag;
  reg        [17:0]   img_reg_array_2_19_real;
  reg        [17:0]   img_reg_array_2_19_imag;
  reg        [17:0]   img_reg_array_2_20_real;
  reg        [17:0]   img_reg_array_2_20_imag;
  reg        [17:0]   img_reg_array_2_21_real;
  reg        [17:0]   img_reg_array_2_21_imag;
  reg        [17:0]   img_reg_array_2_22_real;
  reg        [17:0]   img_reg_array_2_22_imag;
  reg        [17:0]   img_reg_array_2_23_real;
  reg        [17:0]   img_reg_array_2_23_imag;
  reg        [17:0]   img_reg_array_2_24_real;
  reg        [17:0]   img_reg_array_2_24_imag;
  reg        [17:0]   img_reg_array_2_25_real;
  reg        [17:0]   img_reg_array_2_25_imag;
  reg        [17:0]   img_reg_array_2_26_real;
  reg        [17:0]   img_reg_array_2_26_imag;
  reg        [17:0]   img_reg_array_2_27_real;
  reg        [17:0]   img_reg_array_2_27_imag;
  reg        [17:0]   img_reg_array_2_28_real;
  reg        [17:0]   img_reg_array_2_28_imag;
  reg        [17:0]   img_reg_array_2_29_real;
  reg        [17:0]   img_reg_array_2_29_imag;
  reg        [17:0]   img_reg_array_2_30_real;
  reg        [17:0]   img_reg_array_2_30_imag;
  reg        [17:0]   img_reg_array_2_31_real;
  reg        [17:0]   img_reg_array_2_31_imag;
  reg        [17:0]   img_reg_array_2_32_real;
  reg        [17:0]   img_reg_array_2_32_imag;
  reg        [17:0]   img_reg_array_2_33_real;
  reg        [17:0]   img_reg_array_2_33_imag;
  reg        [17:0]   img_reg_array_2_34_real;
  reg        [17:0]   img_reg_array_2_34_imag;
  reg        [17:0]   img_reg_array_2_35_real;
  reg        [17:0]   img_reg_array_2_35_imag;
  reg        [17:0]   img_reg_array_2_36_real;
  reg        [17:0]   img_reg_array_2_36_imag;
  reg        [17:0]   img_reg_array_2_37_real;
  reg        [17:0]   img_reg_array_2_37_imag;
  reg        [17:0]   img_reg_array_2_38_real;
  reg        [17:0]   img_reg_array_2_38_imag;
  reg        [17:0]   img_reg_array_2_39_real;
  reg        [17:0]   img_reg_array_2_39_imag;
  reg        [17:0]   img_reg_array_2_40_real;
  reg        [17:0]   img_reg_array_2_40_imag;
  reg        [17:0]   img_reg_array_2_41_real;
  reg        [17:0]   img_reg_array_2_41_imag;
  reg        [17:0]   img_reg_array_2_42_real;
  reg        [17:0]   img_reg_array_2_42_imag;
  reg        [17:0]   img_reg_array_2_43_real;
  reg        [17:0]   img_reg_array_2_43_imag;
  reg        [17:0]   img_reg_array_2_44_real;
  reg        [17:0]   img_reg_array_2_44_imag;
  reg        [17:0]   img_reg_array_2_45_real;
  reg        [17:0]   img_reg_array_2_45_imag;
  reg        [17:0]   img_reg_array_2_46_real;
  reg        [17:0]   img_reg_array_2_46_imag;
  reg        [17:0]   img_reg_array_2_47_real;
  reg        [17:0]   img_reg_array_2_47_imag;
  reg        [17:0]   img_reg_array_2_48_real;
  reg        [17:0]   img_reg_array_2_48_imag;
  reg        [17:0]   img_reg_array_2_49_real;
  reg        [17:0]   img_reg_array_2_49_imag;
  reg        [17:0]   img_reg_array_2_50_real;
  reg        [17:0]   img_reg_array_2_50_imag;
  reg        [17:0]   img_reg_array_2_51_real;
  reg        [17:0]   img_reg_array_2_51_imag;
  reg        [17:0]   img_reg_array_2_52_real;
  reg        [17:0]   img_reg_array_2_52_imag;
  reg        [17:0]   img_reg_array_2_53_real;
  reg        [17:0]   img_reg_array_2_53_imag;
  reg        [17:0]   img_reg_array_2_54_real;
  reg        [17:0]   img_reg_array_2_54_imag;
  reg        [17:0]   img_reg_array_2_55_real;
  reg        [17:0]   img_reg_array_2_55_imag;
  reg        [17:0]   img_reg_array_2_56_real;
  reg        [17:0]   img_reg_array_2_56_imag;
  reg        [17:0]   img_reg_array_2_57_real;
  reg        [17:0]   img_reg_array_2_57_imag;
  reg        [17:0]   img_reg_array_2_58_real;
  reg        [17:0]   img_reg_array_2_58_imag;
  reg        [17:0]   img_reg_array_2_59_real;
  reg        [17:0]   img_reg_array_2_59_imag;
  reg        [17:0]   img_reg_array_2_60_real;
  reg        [17:0]   img_reg_array_2_60_imag;
  reg        [17:0]   img_reg_array_2_61_real;
  reg        [17:0]   img_reg_array_2_61_imag;
  reg        [17:0]   img_reg_array_2_62_real;
  reg        [17:0]   img_reg_array_2_62_imag;
  reg        [17:0]   img_reg_array_2_63_real;
  reg        [17:0]   img_reg_array_2_63_imag;
  reg        [17:0]   img_reg_array_3_0_real;
  reg        [17:0]   img_reg_array_3_0_imag;
  reg        [17:0]   img_reg_array_3_1_real;
  reg        [17:0]   img_reg_array_3_1_imag;
  reg        [17:0]   img_reg_array_3_2_real;
  reg        [17:0]   img_reg_array_3_2_imag;
  reg        [17:0]   img_reg_array_3_3_real;
  reg        [17:0]   img_reg_array_3_3_imag;
  reg        [17:0]   img_reg_array_3_4_real;
  reg        [17:0]   img_reg_array_3_4_imag;
  reg        [17:0]   img_reg_array_3_5_real;
  reg        [17:0]   img_reg_array_3_5_imag;
  reg        [17:0]   img_reg_array_3_6_real;
  reg        [17:0]   img_reg_array_3_6_imag;
  reg        [17:0]   img_reg_array_3_7_real;
  reg        [17:0]   img_reg_array_3_7_imag;
  reg        [17:0]   img_reg_array_3_8_real;
  reg        [17:0]   img_reg_array_3_8_imag;
  reg        [17:0]   img_reg_array_3_9_real;
  reg        [17:0]   img_reg_array_3_9_imag;
  reg        [17:0]   img_reg_array_3_10_real;
  reg        [17:0]   img_reg_array_3_10_imag;
  reg        [17:0]   img_reg_array_3_11_real;
  reg        [17:0]   img_reg_array_3_11_imag;
  reg        [17:0]   img_reg_array_3_12_real;
  reg        [17:0]   img_reg_array_3_12_imag;
  reg        [17:0]   img_reg_array_3_13_real;
  reg        [17:0]   img_reg_array_3_13_imag;
  reg        [17:0]   img_reg_array_3_14_real;
  reg        [17:0]   img_reg_array_3_14_imag;
  reg        [17:0]   img_reg_array_3_15_real;
  reg        [17:0]   img_reg_array_3_15_imag;
  reg        [17:0]   img_reg_array_3_16_real;
  reg        [17:0]   img_reg_array_3_16_imag;
  reg        [17:0]   img_reg_array_3_17_real;
  reg        [17:0]   img_reg_array_3_17_imag;
  reg        [17:0]   img_reg_array_3_18_real;
  reg        [17:0]   img_reg_array_3_18_imag;
  reg        [17:0]   img_reg_array_3_19_real;
  reg        [17:0]   img_reg_array_3_19_imag;
  reg        [17:0]   img_reg_array_3_20_real;
  reg        [17:0]   img_reg_array_3_20_imag;
  reg        [17:0]   img_reg_array_3_21_real;
  reg        [17:0]   img_reg_array_3_21_imag;
  reg        [17:0]   img_reg_array_3_22_real;
  reg        [17:0]   img_reg_array_3_22_imag;
  reg        [17:0]   img_reg_array_3_23_real;
  reg        [17:0]   img_reg_array_3_23_imag;
  reg        [17:0]   img_reg_array_3_24_real;
  reg        [17:0]   img_reg_array_3_24_imag;
  reg        [17:0]   img_reg_array_3_25_real;
  reg        [17:0]   img_reg_array_3_25_imag;
  reg        [17:0]   img_reg_array_3_26_real;
  reg        [17:0]   img_reg_array_3_26_imag;
  reg        [17:0]   img_reg_array_3_27_real;
  reg        [17:0]   img_reg_array_3_27_imag;
  reg        [17:0]   img_reg_array_3_28_real;
  reg        [17:0]   img_reg_array_3_28_imag;
  reg        [17:0]   img_reg_array_3_29_real;
  reg        [17:0]   img_reg_array_3_29_imag;
  reg        [17:0]   img_reg_array_3_30_real;
  reg        [17:0]   img_reg_array_3_30_imag;
  reg        [17:0]   img_reg_array_3_31_real;
  reg        [17:0]   img_reg_array_3_31_imag;
  reg        [17:0]   img_reg_array_3_32_real;
  reg        [17:0]   img_reg_array_3_32_imag;
  reg        [17:0]   img_reg_array_3_33_real;
  reg        [17:0]   img_reg_array_3_33_imag;
  reg        [17:0]   img_reg_array_3_34_real;
  reg        [17:0]   img_reg_array_3_34_imag;
  reg        [17:0]   img_reg_array_3_35_real;
  reg        [17:0]   img_reg_array_3_35_imag;
  reg        [17:0]   img_reg_array_3_36_real;
  reg        [17:0]   img_reg_array_3_36_imag;
  reg        [17:0]   img_reg_array_3_37_real;
  reg        [17:0]   img_reg_array_3_37_imag;
  reg        [17:0]   img_reg_array_3_38_real;
  reg        [17:0]   img_reg_array_3_38_imag;
  reg        [17:0]   img_reg_array_3_39_real;
  reg        [17:0]   img_reg_array_3_39_imag;
  reg        [17:0]   img_reg_array_3_40_real;
  reg        [17:0]   img_reg_array_3_40_imag;
  reg        [17:0]   img_reg_array_3_41_real;
  reg        [17:0]   img_reg_array_3_41_imag;
  reg        [17:0]   img_reg_array_3_42_real;
  reg        [17:0]   img_reg_array_3_42_imag;
  reg        [17:0]   img_reg_array_3_43_real;
  reg        [17:0]   img_reg_array_3_43_imag;
  reg        [17:0]   img_reg_array_3_44_real;
  reg        [17:0]   img_reg_array_3_44_imag;
  reg        [17:0]   img_reg_array_3_45_real;
  reg        [17:0]   img_reg_array_3_45_imag;
  reg        [17:0]   img_reg_array_3_46_real;
  reg        [17:0]   img_reg_array_3_46_imag;
  reg        [17:0]   img_reg_array_3_47_real;
  reg        [17:0]   img_reg_array_3_47_imag;
  reg        [17:0]   img_reg_array_3_48_real;
  reg        [17:0]   img_reg_array_3_48_imag;
  reg        [17:0]   img_reg_array_3_49_real;
  reg        [17:0]   img_reg_array_3_49_imag;
  reg        [17:0]   img_reg_array_3_50_real;
  reg        [17:0]   img_reg_array_3_50_imag;
  reg        [17:0]   img_reg_array_3_51_real;
  reg        [17:0]   img_reg_array_3_51_imag;
  reg        [17:0]   img_reg_array_3_52_real;
  reg        [17:0]   img_reg_array_3_52_imag;
  reg        [17:0]   img_reg_array_3_53_real;
  reg        [17:0]   img_reg_array_3_53_imag;
  reg        [17:0]   img_reg_array_3_54_real;
  reg        [17:0]   img_reg_array_3_54_imag;
  reg        [17:0]   img_reg_array_3_55_real;
  reg        [17:0]   img_reg_array_3_55_imag;
  reg        [17:0]   img_reg_array_3_56_real;
  reg        [17:0]   img_reg_array_3_56_imag;
  reg        [17:0]   img_reg_array_3_57_real;
  reg        [17:0]   img_reg_array_3_57_imag;
  reg        [17:0]   img_reg_array_3_58_real;
  reg        [17:0]   img_reg_array_3_58_imag;
  reg        [17:0]   img_reg_array_3_59_real;
  reg        [17:0]   img_reg_array_3_59_imag;
  reg        [17:0]   img_reg_array_3_60_real;
  reg        [17:0]   img_reg_array_3_60_imag;
  reg        [17:0]   img_reg_array_3_61_real;
  reg        [17:0]   img_reg_array_3_61_imag;
  reg        [17:0]   img_reg_array_3_62_real;
  reg        [17:0]   img_reg_array_3_62_imag;
  reg        [17:0]   img_reg_array_3_63_real;
  reg        [17:0]   img_reg_array_3_63_imag;
  reg        [17:0]   img_reg_array_4_0_real;
  reg        [17:0]   img_reg_array_4_0_imag;
  reg        [17:0]   img_reg_array_4_1_real;
  reg        [17:0]   img_reg_array_4_1_imag;
  reg        [17:0]   img_reg_array_4_2_real;
  reg        [17:0]   img_reg_array_4_2_imag;
  reg        [17:0]   img_reg_array_4_3_real;
  reg        [17:0]   img_reg_array_4_3_imag;
  reg        [17:0]   img_reg_array_4_4_real;
  reg        [17:0]   img_reg_array_4_4_imag;
  reg        [17:0]   img_reg_array_4_5_real;
  reg        [17:0]   img_reg_array_4_5_imag;
  reg        [17:0]   img_reg_array_4_6_real;
  reg        [17:0]   img_reg_array_4_6_imag;
  reg        [17:0]   img_reg_array_4_7_real;
  reg        [17:0]   img_reg_array_4_7_imag;
  reg        [17:0]   img_reg_array_4_8_real;
  reg        [17:0]   img_reg_array_4_8_imag;
  reg        [17:0]   img_reg_array_4_9_real;
  reg        [17:0]   img_reg_array_4_9_imag;
  reg        [17:0]   img_reg_array_4_10_real;
  reg        [17:0]   img_reg_array_4_10_imag;
  reg        [17:0]   img_reg_array_4_11_real;
  reg        [17:0]   img_reg_array_4_11_imag;
  reg        [17:0]   img_reg_array_4_12_real;
  reg        [17:0]   img_reg_array_4_12_imag;
  reg        [17:0]   img_reg_array_4_13_real;
  reg        [17:0]   img_reg_array_4_13_imag;
  reg        [17:0]   img_reg_array_4_14_real;
  reg        [17:0]   img_reg_array_4_14_imag;
  reg        [17:0]   img_reg_array_4_15_real;
  reg        [17:0]   img_reg_array_4_15_imag;
  reg        [17:0]   img_reg_array_4_16_real;
  reg        [17:0]   img_reg_array_4_16_imag;
  reg        [17:0]   img_reg_array_4_17_real;
  reg        [17:0]   img_reg_array_4_17_imag;
  reg        [17:0]   img_reg_array_4_18_real;
  reg        [17:0]   img_reg_array_4_18_imag;
  reg        [17:0]   img_reg_array_4_19_real;
  reg        [17:0]   img_reg_array_4_19_imag;
  reg        [17:0]   img_reg_array_4_20_real;
  reg        [17:0]   img_reg_array_4_20_imag;
  reg        [17:0]   img_reg_array_4_21_real;
  reg        [17:0]   img_reg_array_4_21_imag;
  reg        [17:0]   img_reg_array_4_22_real;
  reg        [17:0]   img_reg_array_4_22_imag;
  reg        [17:0]   img_reg_array_4_23_real;
  reg        [17:0]   img_reg_array_4_23_imag;
  reg        [17:0]   img_reg_array_4_24_real;
  reg        [17:0]   img_reg_array_4_24_imag;
  reg        [17:0]   img_reg_array_4_25_real;
  reg        [17:0]   img_reg_array_4_25_imag;
  reg        [17:0]   img_reg_array_4_26_real;
  reg        [17:0]   img_reg_array_4_26_imag;
  reg        [17:0]   img_reg_array_4_27_real;
  reg        [17:0]   img_reg_array_4_27_imag;
  reg        [17:0]   img_reg_array_4_28_real;
  reg        [17:0]   img_reg_array_4_28_imag;
  reg        [17:0]   img_reg_array_4_29_real;
  reg        [17:0]   img_reg_array_4_29_imag;
  reg        [17:0]   img_reg_array_4_30_real;
  reg        [17:0]   img_reg_array_4_30_imag;
  reg        [17:0]   img_reg_array_4_31_real;
  reg        [17:0]   img_reg_array_4_31_imag;
  reg        [17:0]   img_reg_array_4_32_real;
  reg        [17:0]   img_reg_array_4_32_imag;
  reg        [17:0]   img_reg_array_4_33_real;
  reg        [17:0]   img_reg_array_4_33_imag;
  reg        [17:0]   img_reg_array_4_34_real;
  reg        [17:0]   img_reg_array_4_34_imag;
  reg        [17:0]   img_reg_array_4_35_real;
  reg        [17:0]   img_reg_array_4_35_imag;
  reg        [17:0]   img_reg_array_4_36_real;
  reg        [17:0]   img_reg_array_4_36_imag;
  reg        [17:0]   img_reg_array_4_37_real;
  reg        [17:0]   img_reg_array_4_37_imag;
  reg        [17:0]   img_reg_array_4_38_real;
  reg        [17:0]   img_reg_array_4_38_imag;
  reg        [17:0]   img_reg_array_4_39_real;
  reg        [17:0]   img_reg_array_4_39_imag;
  reg        [17:0]   img_reg_array_4_40_real;
  reg        [17:0]   img_reg_array_4_40_imag;
  reg        [17:0]   img_reg_array_4_41_real;
  reg        [17:0]   img_reg_array_4_41_imag;
  reg        [17:0]   img_reg_array_4_42_real;
  reg        [17:0]   img_reg_array_4_42_imag;
  reg        [17:0]   img_reg_array_4_43_real;
  reg        [17:0]   img_reg_array_4_43_imag;
  reg        [17:0]   img_reg_array_4_44_real;
  reg        [17:0]   img_reg_array_4_44_imag;
  reg        [17:0]   img_reg_array_4_45_real;
  reg        [17:0]   img_reg_array_4_45_imag;
  reg        [17:0]   img_reg_array_4_46_real;
  reg        [17:0]   img_reg_array_4_46_imag;
  reg        [17:0]   img_reg_array_4_47_real;
  reg        [17:0]   img_reg_array_4_47_imag;
  reg        [17:0]   img_reg_array_4_48_real;
  reg        [17:0]   img_reg_array_4_48_imag;
  reg        [17:0]   img_reg_array_4_49_real;
  reg        [17:0]   img_reg_array_4_49_imag;
  reg        [17:0]   img_reg_array_4_50_real;
  reg        [17:0]   img_reg_array_4_50_imag;
  reg        [17:0]   img_reg_array_4_51_real;
  reg        [17:0]   img_reg_array_4_51_imag;
  reg        [17:0]   img_reg_array_4_52_real;
  reg        [17:0]   img_reg_array_4_52_imag;
  reg        [17:0]   img_reg_array_4_53_real;
  reg        [17:0]   img_reg_array_4_53_imag;
  reg        [17:0]   img_reg_array_4_54_real;
  reg        [17:0]   img_reg_array_4_54_imag;
  reg        [17:0]   img_reg_array_4_55_real;
  reg        [17:0]   img_reg_array_4_55_imag;
  reg        [17:0]   img_reg_array_4_56_real;
  reg        [17:0]   img_reg_array_4_56_imag;
  reg        [17:0]   img_reg_array_4_57_real;
  reg        [17:0]   img_reg_array_4_57_imag;
  reg        [17:0]   img_reg_array_4_58_real;
  reg        [17:0]   img_reg_array_4_58_imag;
  reg        [17:0]   img_reg_array_4_59_real;
  reg        [17:0]   img_reg_array_4_59_imag;
  reg        [17:0]   img_reg_array_4_60_real;
  reg        [17:0]   img_reg_array_4_60_imag;
  reg        [17:0]   img_reg_array_4_61_real;
  reg        [17:0]   img_reg_array_4_61_imag;
  reg        [17:0]   img_reg_array_4_62_real;
  reg        [17:0]   img_reg_array_4_62_imag;
  reg        [17:0]   img_reg_array_4_63_real;
  reg        [17:0]   img_reg_array_4_63_imag;
  reg        [17:0]   img_reg_array_5_0_real;
  reg        [17:0]   img_reg_array_5_0_imag;
  reg        [17:0]   img_reg_array_5_1_real;
  reg        [17:0]   img_reg_array_5_1_imag;
  reg        [17:0]   img_reg_array_5_2_real;
  reg        [17:0]   img_reg_array_5_2_imag;
  reg        [17:0]   img_reg_array_5_3_real;
  reg        [17:0]   img_reg_array_5_3_imag;
  reg        [17:0]   img_reg_array_5_4_real;
  reg        [17:0]   img_reg_array_5_4_imag;
  reg        [17:0]   img_reg_array_5_5_real;
  reg        [17:0]   img_reg_array_5_5_imag;
  reg        [17:0]   img_reg_array_5_6_real;
  reg        [17:0]   img_reg_array_5_6_imag;
  reg        [17:0]   img_reg_array_5_7_real;
  reg        [17:0]   img_reg_array_5_7_imag;
  reg        [17:0]   img_reg_array_5_8_real;
  reg        [17:0]   img_reg_array_5_8_imag;
  reg        [17:0]   img_reg_array_5_9_real;
  reg        [17:0]   img_reg_array_5_9_imag;
  reg        [17:0]   img_reg_array_5_10_real;
  reg        [17:0]   img_reg_array_5_10_imag;
  reg        [17:0]   img_reg_array_5_11_real;
  reg        [17:0]   img_reg_array_5_11_imag;
  reg        [17:0]   img_reg_array_5_12_real;
  reg        [17:0]   img_reg_array_5_12_imag;
  reg        [17:0]   img_reg_array_5_13_real;
  reg        [17:0]   img_reg_array_5_13_imag;
  reg        [17:0]   img_reg_array_5_14_real;
  reg        [17:0]   img_reg_array_5_14_imag;
  reg        [17:0]   img_reg_array_5_15_real;
  reg        [17:0]   img_reg_array_5_15_imag;
  reg        [17:0]   img_reg_array_5_16_real;
  reg        [17:0]   img_reg_array_5_16_imag;
  reg        [17:0]   img_reg_array_5_17_real;
  reg        [17:0]   img_reg_array_5_17_imag;
  reg        [17:0]   img_reg_array_5_18_real;
  reg        [17:0]   img_reg_array_5_18_imag;
  reg        [17:0]   img_reg_array_5_19_real;
  reg        [17:0]   img_reg_array_5_19_imag;
  reg        [17:0]   img_reg_array_5_20_real;
  reg        [17:0]   img_reg_array_5_20_imag;
  reg        [17:0]   img_reg_array_5_21_real;
  reg        [17:0]   img_reg_array_5_21_imag;
  reg        [17:0]   img_reg_array_5_22_real;
  reg        [17:0]   img_reg_array_5_22_imag;
  reg        [17:0]   img_reg_array_5_23_real;
  reg        [17:0]   img_reg_array_5_23_imag;
  reg        [17:0]   img_reg_array_5_24_real;
  reg        [17:0]   img_reg_array_5_24_imag;
  reg        [17:0]   img_reg_array_5_25_real;
  reg        [17:0]   img_reg_array_5_25_imag;
  reg        [17:0]   img_reg_array_5_26_real;
  reg        [17:0]   img_reg_array_5_26_imag;
  reg        [17:0]   img_reg_array_5_27_real;
  reg        [17:0]   img_reg_array_5_27_imag;
  reg        [17:0]   img_reg_array_5_28_real;
  reg        [17:0]   img_reg_array_5_28_imag;
  reg        [17:0]   img_reg_array_5_29_real;
  reg        [17:0]   img_reg_array_5_29_imag;
  reg        [17:0]   img_reg_array_5_30_real;
  reg        [17:0]   img_reg_array_5_30_imag;
  reg        [17:0]   img_reg_array_5_31_real;
  reg        [17:0]   img_reg_array_5_31_imag;
  reg        [17:0]   img_reg_array_5_32_real;
  reg        [17:0]   img_reg_array_5_32_imag;
  reg        [17:0]   img_reg_array_5_33_real;
  reg        [17:0]   img_reg_array_5_33_imag;
  reg        [17:0]   img_reg_array_5_34_real;
  reg        [17:0]   img_reg_array_5_34_imag;
  reg        [17:0]   img_reg_array_5_35_real;
  reg        [17:0]   img_reg_array_5_35_imag;
  reg        [17:0]   img_reg_array_5_36_real;
  reg        [17:0]   img_reg_array_5_36_imag;
  reg        [17:0]   img_reg_array_5_37_real;
  reg        [17:0]   img_reg_array_5_37_imag;
  reg        [17:0]   img_reg_array_5_38_real;
  reg        [17:0]   img_reg_array_5_38_imag;
  reg        [17:0]   img_reg_array_5_39_real;
  reg        [17:0]   img_reg_array_5_39_imag;
  reg        [17:0]   img_reg_array_5_40_real;
  reg        [17:0]   img_reg_array_5_40_imag;
  reg        [17:0]   img_reg_array_5_41_real;
  reg        [17:0]   img_reg_array_5_41_imag;
  reg        [17:0]   img_reg_array_5_42_real;
  reg        [17:0]   img_reg_array_5_42_imag;
  reg        [17:0]   img_reg_array_5_43_real;
  reg        [17:0]   img_reg_array_5_43_imag;
  reg        [17:0]   img_reg_array_5_44_real;
  reg        [17:0]   img_reg_array_5_44_imag;
  reg        [17:0]   img_reg_array_5_45_real;
  reg        [17:0]   img_reg_array_5_45_imag;
  reg        [17:0]   img_reg_array_5_46_real;
  reg        [17:0]   img_reg_array_5_46_imag;
  reg        [17:0]   img_reg_array_5_47_real;
  reg        [17:0]   img_reg_array_5_47_imag;
  reg        [17:0]   img_reg_array_5_48_real;
  reg        [17:0]   img_reg_array_5_48_imag;
  reg        [17:0]   img_reg_array_5_49_real;
  reg        [17:0]   img_reg_array_5_49_imag;
  reg        [17:0]   img_reg_array_5_50_real;
  reg        [17:0]   img_reg_array_5_50_imag;
  reg        [17:0]   img_reg_array_5_51_real;
  reg        [17:0]   img_reg_array_5_51_imag;
  reg        [17:0]   img_reg_array_5_52_real;
  reg        [17:0]   img_reg_array_5_52_imag;
  reg        [17:0]   img_reg_array_5_53_real;
  reg        [17:0]   img_reg_array_5_53_imag;
  reg        [17:0]   img_reg_array_5_54_real;
  reg        [17:0]   img_reg_array_5_54_imag;
  reg        [17:0]   img_reg_array_5_55_real;
  reg        [17:0]   img_reg_array_5_55_imag;
  reg        [17:0]   img_reg_array_5_56_real;
  reg        [17:0]   img_reg_array_5_56_imag;
  reg        [17:0]   img_reg_array_5_57_real;
  reg        [17:0]   img_reg_array_5_57_imag;
  reg        [17:0]   img_reg_array_5_58_real;
  reg        [17:0]   img_reg_array_5_58_imag;
  reg        [17:0]   img_reg_array_5_59_real;
  reg        [17:0]   img_reg_array_5_59_imag;
  reg        [17:0]   img_reg_array_5_60_real;
  reg        [17:0]   img_reg_array_5_60_imag;
  reg        [17:0]   img_reg_array_5_61_real;
  reg        [17:0]   img_reg_array_5_61_imag;
  reg        [17:0]   img_reg_array_5_62_real;
  reg        [17:0]   img_reg_array_5_62_imag;
  reg        [17:0]   img_reg_array_5_63_real;
  reg        [17:0]   img_reg_array_5_63_imag;
  reg        [17:0]   img_reg_array_6_0_real;
  reg        [17:0]   img_reg_array_6_0_imag;
  reg        [17:0]   img_reg_array_6_1_real;
  reg        [17:0]   img_reg_array_6_1_imag;
  reg        [17:0]   img_reg_array_6_2_real;
  reg        [17:0]   img_reg_array_6_2_imag;
  reg        [17:0]   img_reg_array_6_3_real;
  reg        [17:0]   img_reg_array_6_3_imag;
  reg        [17:0]   img_reg_array_6_4_real;
  reg        [17:0]   img_reg_array_6_4_imag;
  reg        [17:0]   img_reg_array_6_5_real;
  reg        [17:0]   img_reg_array_6_5_imag;
  reg        [17:0]   img_reg_array_6_6_real;
  reg        [17:0]   img_reg_array_6_6_imag;
  reg        [17:0]   img_reg_array_6_7_real;
  reg        [17:0]   img_reg_array_6_7_imag;
  reg        [17:0]   img_reg_array_6_8_real;
  reg        [17:0]   img_reg_array_6_8_imag;
  reg        [17:0]   img_reg_array_6_9_real;
  reg        [17:0]   img_reg_array_6_9_imag;
  reg        [17:0]   img_reg_array_6_10_real;
  reg        [17:0]   img_reg_array_6_10_imag;
  reg        [17:0]   img_reg_array_6_11_real;
  reg        [17:0]   img_reg_array_6_11_imag;
  reg        [17:0]   img_reg_array_6_12_real;
  reg        [17:0]   img_reg_array_6_12_imag;
  reg        [17:0]   img_reg_array_6_13_real;
  reg        [17:0]   img_reg_array_6_13_imag;
  reg        [17:0]   img_reg_array_6_14_real;
  reg        [17:0]   img_reg_array_6_14_imag;
  reg        [17:0]   img_reg_array_6_15_real;
  reg        [17:0]   img_reg_array_6_15_imag;
  reg        [17:0]   img_reg_array_6_16_real;
  reg        [17:0]   img_reg_array_6_16_imag;
  reg        [17:0]   img_reg_array_6_17_real;
  reg        [17:0]   img_reg_array_6_17_imag;
  reg        [17:0]   img_reg_array_6_18_real;
  reg        [17:0]   img_reg_array_6_18_imag;
  reg        [17:0]   img_reg_array_6_19_real;
  reg        [17:0]   img_reg_array_6_19_imag;
  reg        [17:0]   img_reg_array_6_20_real;
  reg        [17:0]   img_reg_array_6_20_imag;
  reg        [17:0]   img_reg_array_6_21_real;
  reg        [17:0]   img_reg_array_6_21_imag;
  reg        [17:0]   img_reg_array_6_22_real;
  reg        [17:0]   img_reg_array_6_22_imag;
  reg        [17:0]   img_reg_array_6_23_real;
  reg        [17:0]   img_reg_array_6_23_imag;
  reg        [17:0]   img_reg_array_6_24_real;
  reg        [17:0]   img_reg_array_6_24_imag;
  reg        [17:0]   img_reg_array_6_25_real;
  reg        [17:0]   img_reg_array_6_25_imag;
  reg        [17:0]   img_reg_array_6_26_real;
  reg        [17:0]   img_reg_array_6_26_imag;
  reg        [17:0]   img_reg_array_6_27_real;
  reg        [17:0]   img_reg_array_6_27_imag;
  reg        [17:0]   img_reg_array_6_28_real;
  reg        [17:0]   img_reg_array_6_28_imag;
  reg        [17:0]   img_reg_array_6_29_real;
  reg        [17:0]   img_reg_array_6_29_imag;
  reg        [17:0]   img_reg_array_6_30_real;
  reg        [17:0]   img_reg_array_6_30_imag;
  reg        [17:0]   img_reg_array_6_31_real;
  reg        [17:0]   img_reg_array_6_31_imag;
  reg        [17:0]   img_reg_array_6_32_real;
  reg        [17:0]   img_reg_array_6_32_imag;
  reg        [17:0]   img_reg_array_6_33_real;
  reg        [17:0]   img_reg_array_6_33_imag;
  reg        [17:0]   img_reg_array_6_34_real;
  reg        [17:0]   img_reg_array_6_34_imag;
  reg        [17:0]   img_reg_array_6_35_real;
  reg        [17:0]   img_reg_array_6_35_imag;
  reg        [17:0]   img_reg_array_6_36_real;
  reg        [17:0]   img_reg_array_6_36_imag;
  reg        [17:0]   img_reg_array_6_37_real;
  reg        [17:0]   img_reg_array_6_37_imag;
  reg        [17:0]   img_reg_array_6_38_real;
  reg        [17:0]   img_reg_array_6_38_imag;
  reg        [17:0]   img_reg_array_6_39_real;
  reg        [17:0]   img_reg_array_6_39_imag;
  reg        [17:0]   img_reg_array_6_40_real;
  reg        [17:0]   img_reg_array_6_40_imag;
  reg        [17:0]   img_reg_array_6_41_real;
  reg        [17:0]   img_reg_array_6_41_imag;
  reg        [17:0]   img_reg_array_6_42_real;
  reg        [17:0]   img_reg_array_6_42_imag;
  reg        [17:0]   img_reg_array_6_43_real;
  reg        [17:0]   img_reg_array_6_43_imag;
  reg        [17:0]   img_reg_array_6_44_real;
  reg        [17:0]   img_reg_array_6_44_imag;
  reg        [17:0]   img_reg_array_6_45_real;
  reg        [17:0]   img_reg_array_6_45_imag;
  reg        [17:0]   img_reg_array_6_46_real;
  reg        [17:0]   img_reg_array_6_46_imag;
  reg        [17:0]   img_reg_array_6_47_real;
  reg        [17:0]   img_reg_array_6_47_imag;
  reg        [17:0]   img_reg_array_6_48_real;
  reg        [17:0]   img_reg_array_6_48_imag;
  reg        [17:0]   img_reg_array_6_49_real;
  reg        [17:0]   img_reg_array_6_49_imag;
  reg        [17:0]   img_reg_array_6_50_real;
  reg        [17:0]   img_reg_array_6_50_imag;
  reg        [17:0]   img_reg_array_6_51_real;
  reg        [17:0]   img_reg_array_6_51_imag;
  reg        [17:0]   img_reg_array_6_52_real;
  reg        [17:0]   img_reg_array_6_52_imag;
  reg        [17:0]   img_reg_array_6_53_real;
  reg        [17:0]   img_reg_array_6_53_imag;
  reg        [17:0]   img_reg_array_6_54_real;
  reg        [17:0]   img_reg_array_6_54_imag;
  reg        [17:0]   img_reg_array_6_55_real;
  reg        [17:0]   img_reg_array_6_55_imag;
  reg        [17:0]   img_reg_array_6_56_real;
  reg        [17:0]   img_reg_array_6_56_imag;
  reg        [17:0]   img_reg_array_6_57_real;
  reg        [17:0]   img_reg_array_6_57_imag;
  reg        [17:0]   img_reg_array_6_58_real;
  reg        [17:0]   img_reg_array_6_58_imag;
  reg        [17:0]   img_reg_array_6_59_real;
  reg        [17:0]   img_reg_array_6_59_imag;
  reg        [17:0]   img_reg_array_6_60_real;
  reg        [17:0]   img_reg_array_6_60_imag;
  reg        [17:0]   img_reg_array_6_61_real;
  reg        [17:0]   img_reg_array_6_61_imag;
  reg        [17:0]   img_reg_array_6_62_real;
  reg        [17:0]   img_reg_array_6_62_imag;
  reg        [17:0]   img_reg_array_6_63_real;
  reg        [17:0]   img_reg_array_6_63_imag;
  reg        [17:0]   img_reg_array_7_0_real;
  reg        [17:0]   img_reg_array_7_0_imag;
  reg        [17:0]   img_reg_array_7_1_real;
  reg        [17:0]   img_reg_array_7_1_imag;
  reg        [17:0]   img_reg_array_7_2_real;
  reg        [17:0]   img_reg_array_7_2_imag;
  reg        [17:0]   img_reg_array_7_3_real;
  reg        [17:0]   img_reg_array_7_3_imag;
  reg        [17:0]   img_reg_array_7_4_real;
  reg        [17:0]   img_reg_array_7_4_imag;
  reg        [17:0]   img_reg_array_7_5_real;
  reg        [17:0]   img_reg_array_7_5_imag;
  reg        [17:0]   img_reg_array_7_6_real;
  reg        [17:0]   img_reg_array_7_6_imag;
  reg        [17:0]   img_reg_array_7_7_real;
  reg        [17:0]   img_reg_array_7_7_imag;
  reg        [17:0]   img_reg_array_7_8_real;
  reg        [17:0]   img_reg_array_7_8_imag;
  reg        [17:0]   img_reg_array_7_9_real;
  reg        [17:0]   img_reg_array_7_9_imag;
  reg        [17:0]   img_reg_array_7_10_real;
  reg        [17:0]   img_reg_array_7_10_imag;
  reg        [17:0]   img_reg_array_7_11_real;
  reg        [17:0]   img_reg_array_7_11_imag;
  reg        [17:0]   img_reg_array_7_12_real;
  reg        [17:0]   img_reg_array_7_12_imag;
  reg        [17:0]   img_reg_array_7_13_real;
  reg        [17:0]   img_reg_array_7_13_imag;
  reg        [17:0]   img_reg_array_7_14_real;
  reg        [17:0]   img_reg_array_7_14_imag;
  reg        [17:0]   img_reg_array_7_15_real;
  reg        [17:0]   img_reg_array_7_15_imag;
  reg        [17:0]   img_reg_array_7_16_real;
  reg        [17:0]   img_reg_array_7_16_imag;
  reg        [17:0]   img_reg_array_7_17_real;
  reg        [17:0]   img_reg_array_7_17_imag;
  reg        [17:0]   img_reg_array_7_18_real;
  reg        [17:0]   img_reg_array_7_18_imag;
  reg        [17:0]   img_reg_array_7_19_real;
  reg        [17:0]   img_reg_array_7_19_imag;
  reg        [17:0]   img_reg_array_7_20_real;
  reg        [17:0]   img_reg_array_7_20_imag;
  reg        [17:0]   img_reg_array_7_21_real;
  reg        [17:0]   img_reg_array_7_21_imag;
  reg        [17:0]   img_reg_array_7_22_real;
  reg        [17:0]   img_reg_array_7_22_imag;
  reg        [17:0]   img_reg_array_7_23_real;
  reg        [17:0]   img_reg_array_7_23_imag;
  reg        [17:0]   img_reg_array_7_24_real;
  reg        [17:0]   img_reg_array_7_24_imag;
  reg        [17:0]   img_reg_array_7_25_real;
  reg        [17:0]   img_reg_array_7_25_imag;
  reg        [17:0]   img_reg_array_7_26_real;
  reg        [17:0]   img_reg_array_7_26_imag;
  reg        [17:0]   img_reg_array_7_27_real;
  reg        [17:0]   img_reg_array_7_27_imag;
  reg        [17:0]   img_reg_array_7_28_real;
  reg        [17:0]   img_reg_array_7_28_imag;
  reg        [17:0]   img_reg_array_7_29_real;
  reg        [17:0]   img_reg_array_7_29_imag;
  reg        [17:0]   img_reg_array_7_30_real;
  reg        [17:0]   img_reg_array_7_30_imag;
  reg        [17:0]   img_reg_array_7_31_real;
  reg        [17:0]   img_reg_array_7_31_imag;
  reg        [17:0]   img_reg_array_7_32_real;
  reg        [17:0]   img_reg_array_7_32_imag;
  reg        [17:0]   img_reg_array_7_33_real;
  reg        [17:0]   img_reg_array_7_33_imag;
  reg        [17:0]   img_reg_array_7_34_real;
  reg        [17:0]   img_reg_array_7_34_imag;
  reg        [17:0]   img_reg_array_7_35_real;
  reg        [17:0]   img_reg_array_7_35_imag;
  reg        [17:0]   img_reg_array_7_36_real;
  reg        [17:0]   img_reg_array_7_36_imag;
  reg        [17:0]   img_reg_array_7_37_real;
  reg        [17:0]   img_reg_array_7_37_imag;
  reg        [17:0]   img_reg_array_7_38_real;
  reg        [17:0]   img_reg_array_7_38_imag;
  reg        [17:0]   img_reg_array_7_39_real;
  reg        [17:0]   img_reg_array_7_39_imag;
  reg        [17:0]   img_reg_array_7_40_real;
  reg        [17:0]   img_reg_array_7_40_imag;
  reg        [17:0]   img_reg_array_7_41_real;
  reg        [17:0]   img_reg_array_7_41_imag;
  reg        [17:0]   img_reg_array_7_42_real;
  reg        [17:0]   img_reg_array_7_42_imag;
  reg        [17:0]   img_reg_array_7_43_real;
  reg        [17:0]   img_reg_array_7_43_imag;
  reg        [17:0]   img_reg_array_7_44_real;
  reg        [17:0]   img_reg_array_7_44_imag;
  reg        [17:0]   img_reg_array_7_45_real;
  reg        [17:0]   img_reg_array_7_45_imag;
  reg        [17:0]   img_reg_array_7_46_real;
  reg        [17:0]   img_reg_array_7_46_imag;
  reg        [17:0]   img_reg_array_7_47_real;
  reg        [17:0]   img_reg_array_7_47_imag;
  reg        [17:0]   img_reg_array_7_48_real;
  reg        [17:0]   img_reg_array_7_48_imag;
  reg        [17:0]   img_reg_array_7_49_real;
  reg        [17:0]   img_reg_array_7_49_imag;
  reg        [17:0]   img_reg_array_7_50_real;
  reg        [17:0]   img_reg_array_7_50_imag;
  reg        [17:0]   img_reg_array_7_51_real;
  reg        [17:0]   img_reg_array_7_51_imag;
  reg        [17:0]   img_reg_array_7_52_real;
  reg        [17:0]   img_reg_array_7_52_imag;
  reg        [17:0]   img_reg_array_7_53_real;
  reg        [17:0]   img_reg_array_7_53_imag;
  reg        [17:0]   img_reg_array_7_54_real;
  reg        [17:0]   img_reg_array_7_54_imag;
  reg        [17:0]   img_reg_array_7_55_real;
  reg        [17:0]   img_reg_array_7_55_imag;
  reg        [17:0]   img_reg_array_7_56_real;
  reg        [17:0]   img_reg_array_7_56_imag;
  reg        [17:0]   img_reg_array_7_57_real;
  reg        [17:0]   img_reg_array_7_57_imag;
  reg        [17:0]   img_reg_array_7_58_real;
  reg        [17:0]   img_reg_array_7_58_imag;
  reg        [17:0]   img_reg_array_7_59_real;
  reg        [17:0]   img_reg_array_7_59_imag;
  reg        [17:0]   img_reg_array_7_60_real;
  reg        [17:0]   img_reg_array_7_60_imag;
  reg        [17:0]   img_reg_array_7_61_real;
  reg        [17:0]   img_reg_array_7_61_imag;
  reg        [17:0]   img_reg_array_7_62_real;
  reg        [17:0]   img_reg_array_7_62_imag;
  reg        [17:0]   img_reg_array_7_63_real;
  reg        [17:0]   img_reg_array_7_63_imag;
  reg        [17:0]   img_reg_array_8_0_real;
  reg        [17:0]   img_reg_array_8_0_imag;
  reg        [17:0]   img_reg_array_8_1_real;
  reg        [17:0]   img_reg_array_8_1_imag;
  reg        [17:0]   img_reg_array_8_2_real;
  reg        [17:0]   img_reg_array_8_2_imag;
  reg        [17:0]   img_reg_array_8_3_real;
  reg        [17:0]   img_reg_array_8_3_imag;
  reg        [17:0]   img_reg_array_8_4_real;
  reg        [17:0]   img_reg_array_8_4_imag;
  reg        [17:0]   img_reg_array_8_5_real;
  reg        [17:0]   img_reg_array_8_5_imag;
  reg        [17:0]   img_reg_array_8_6_real;
  reg        [17:0]   img_reg_array_8_6_imag;
  reg        [17:0]   img_reg_array_8_7_real;
  reg        [17:0]   img_reg_array_8_7_imag;
  reg        [17:0]   img_reg_array_8_8_real;
  reg        [17:0]   img_reg_array_8_8_imag;
  reg        [17:0]   img_reg_array_8_9_real;
  reg        [17:0]   img_reg_array_8_9_imag;
  reg        [17:0]   img_reg_array_8_10_real;
  reg        [17:0]   img_reg_array_8_10_imag;
  reg        [17:0]   img_reg_array_8_11_real;
  reg        [17:0]   img_reg_array_8_11_imag;
  reg        [17:0]   img_reg_array_8_12_real;
  reg        [17:0]   img_reg_array_8_12_imag;
  reg        [17:0]   img_reg_array_8_13_real;
  reg        [17:0]   img_reg_array_8_13_imag;
  reg        [17:0]   img_reg_array_8_14_real;
  reg        [17:0]   img_reg_array_8_14_imag;
  reg        [17:0]   img_reg_array_8_15_real;
  reg        [17:0]   img_reg_array_8_15_imag;
  reg        [17:0]   img_reg_array_8_16_real;
  reg        [17:0]   img_reg_array_8_16_imag;
  reg        [17:0]   img_reg_array_8_17_real;
  reg        [17:0]   img_reg_array_8_17_imag;
  reg        [17:0]   img_reg_array_8_18_real;
  reg        [17:0]   img_reg_array_8_18_imag;
  reg        [17:0]   img_reg_array_8_19_real;
  reg        [17:0]   img_reg_array_8_19_imag;
  reg        [17:0]   img_reg_array_8_20_real;
  reg        [17:0]   img_reg_array_8_20_imag;
  reg        [17:0]   img_reg_array_8_21_real;
  reg        [17:0]   img_reg_array_8_21_imag;
  reg        [17:0]   img_reg_array_8_22_real;
  reg        [17:0]   img_reg_array_8_22_imag;
  reg        [17:0]   img_reg_array_8_23_real;
  reg        [17:0]   img_reg_array_8_23_imag;
  reg        [17:0]   img_reg_array_8_24_real;
  reg        [17:0]   img_reg_array_8_24_imag;
  reg        [17:0]   img_reg_array_8_25_real;
  reg        [17:0]   img_reg_array_8_25_imag;
  reg        [17:0]   img_reg_array_8_26_real;
  reg        [17:0]   img_reg_array_8_26_imag;
  reg        [17:0]   img_reg_array_8_27_real;
  reg        [17:0]   img_reg_array_8_27_imag;
  reg        [17:0]   img_reg_array_8_28_real;
  reg        [17:0]   img_reg_array_8_28_imag;
  reg        [17:0]   img_reg_array_8_29_real;
  reg        [17:0]   img_reg_array_8_29_imag;
  reg        [17:0]   img_reg_array_8_30_real;
  reg        [17:0]   img_reg_array_8_30_imag;
  reg        [17:0]   img_reg_array_8_31_real;
  reg        [17:0]   img_reg_array_8_31_imag;
  reg        [17:0]   img_reg_array_8_32_real;
  reg        [17:0]   img_reg_array_8_32_imag;
  reg        [17:0]   img_reg_array_8_33_real;
  reg        [17:0]   img_reg_array_8_33_imag;
  reg        [17:0]   img_reg_array_8_34_real;
  reg        [17:0]   img_reg_array_8_34_imag;
  reg        [17:0]   img_reg_array_8_35_real;
  reg        [17:0]   img_reg_array_8_35_imag;
  reg        [17:0]   img_reg_array_8_36_real;
  reg        [17:0]   img_reg_array_8_36_imag;
  reg        [17:0]   img_reg_array_8_37_real;
  reg        [17:0]   img_reg_array_8_37_imag;
  reg        [17:0]   img_reg_array_8_38_real;
  reg        [17:0]   img_reg_array_8_38_imag;
  reg        [17:0]   img_reg_array_8_39_real;
  reg        [17:0]   img_reg_array_8_39_imag;
  reg        [17:0]   img_reg_array_8_40_real;
  reg        [17:0]   img_reg_array_8_40_imag;
  reg        [17:0]   img_reg_array_8_41_real;
  reg        [17:0]   img_reg_array_8_41_imag;
  reg        [17:0]   img_reg_array_8_42_real;
  reg        [17:0]   img_reg_array_8_42_imag;
  reg        [17:0]   img_reg_array_8_43_real;
  reg        [17:0]   img_reg_array_8_43_imag;
  reg        [17:0]   img_reg_array_8_44_real;
  reg        [17:0]   img_reg_array_8_44_imag;
  reg        [17:0]   img_reg_array_8_45_real;
  reg        [17:0]   img_reg_array_8_45_imag;
  reg        [17:0]   img_reg_array_8_46_real;
  reg        [17:0]   img_reg_array_8_46_imag;
  reg        [17:0]   img_reg_array_8_47_real;
  reg        [17:0]   img_reg_array_8_47_imag;
  reg        [17:0]   img_reg_array_8_48_real;
  reg        [17:0]   img_reg_array_8_48_imag;
  reg        [17:0]   img_reg_array_8_49_real;
  reg        [17:0]   img_reg_array_8_49_imag;
  reg        [17:0]   img_reg_array_8_50_real;
  reg        [17:0]   img_reg_array_8_50_imag;
  reg        [17:0]   img_reg_array_8_51_real;
  reg        [17:0]   img_reg_array_8_51_imag;
  reg        [17:0]   img_reg_array_8_52_real;
  reg        [17:0]   img_reg_array_8_52_imag;
  reg        [17:0]   img_reg_array_8_53_real;
  reg        [17:0]   img_reg_array_8_53_imag;
  reg        [17:0]   img_reg_array_8_54_real;
  reg        [17:0]   img_reg_array_8_54_imag;
  reg        [17:0]   img_reg_array_8_55_real;
  reg        [17:0]   img_reg_array_8_55_imag;
  reg        [17:0]   img_reg_array_8_56_real;
  reg        [17:0]   img_reg_array_8_56_imag;
  reg        [17:0]   img_reg_array_8_57_real;
  reg        [17:0]   img_reg_array_8_57_imag;
  reg        [17:0]   img_reg_array_8_58_real;
  reg        [17:0]   img_reg_array_8_58_imag;
  reg        [17:0]   img_reg_array_8_59_real;
  reg        [17:0]   img_reg_array_8_59_imag;
  reg        [17:0]   img_reg_array_8_60_real;
  reg        [17:0]   img_reg_array_8_60_imag;
  reg        [17:0]   img_reg_array_8_61_real;
  reg        [17:0]   img_reg_array_8_61_imag;
  reg        [17:0]   img_reg_array_8_62_real;
  reg        [17:0]   img_reg_array_8_62_imag;
  reg        [17:0]   img_reg_array_8_63_real;
  reg        [17:0]   img_reg_array_8_63_imag;
  reg        [17:0]   img_reg_array_9_0_real;
  reg        [17:0]   img_reg_array_9_0_imag;
  reg        [17:0]   img_reg_array_9_1_real;
  reg        [17:0]   img_reg_array_9_1_imag;
  reg        [17:0]   img_reg_array_9_2_real;
  reg        [17:0]   img_reg_array_9_2_imag;
  reg        [17:0]   img_reg_array_9_3_real;
  reg        [17:0]   img_reg_array_9_3_imag;
  reg        [17:0]   img_reg_array_9_4_real;
  reg        [17:0]   img_reg_array_9_4_imag;
  reg        [17:0]   img_reg_array_9_5_real;
  reg        [17:0]   img_reg_array_9_5_imag;
  reg        [17:0]   img_reg_array_9_6_real;
  reg        [17:0]   img_reg_array_9_6_imag;
  reg        [17:0]   img_reg_array_9_7_real;
  reg        [17:0]   img_reg_array_9_7_imag;
  reg        [17:0]   img_reg_array_9_8_real;
  reg        [17:0]   img_reg_array_9_8_imag;
  reg        [17:0]   img_reg_array_9_9_real;
  reg        [17:0]   img_reg_array_9_9_imag;
  reg        [17:0]   img_reg_array_9_10_real;
  reg        [17:0]   img_reg_array_9_10_imag;
  reg        [17:0]   img_reg_array_9_11_real;
  reg        [17:0]   img_reg_array_9_11_imag;
  reg        [17:0]   img_reg_array_9_12_real;
  reg        [17:0]   img_reg_array_9_12_imag;
  reg        [17:0]   img_reg_array_9_13_real;
  reg        [17:0]   img_reg_array_9_13_imag;
  reg        [17:0]   img_reg_array_9_14_real;
  reg        [17:0]   img_reg_array_9_14_imag;
  reg        [17:0]   img_reg_array_9_15_real;
  reg        [17:0]   img_reg_array_9_15_imag;
  reg        [17:0]   img_reg_array_9_16_real;
  reg        [17:0]   img_reg_array_9_16_imag;
  reg        [17:0]   img_reg_array_9_17_real;
  reg        [17:0]   img_reg_array_9_17_imag;
  reg        [17:0]   img_reg_array_9_18_real;
  reg        [17:0]   img_reg_array_9_18_imag;
  reg        [17:0]   img_reg_array_9_19_real;
  reg        [17:0]   img_reg_array_9_19_imag;
  reg        [17:0]   img_reg_array_9_20_real;
  reg        [17:0]   img_reg_array_9_20_imag;
  reg        [17:0]   img_reg_array_9_21_real;
  reg        [17:0]   img_reg_array_9_21_imag;
  reg        [17:0]   img_reg_array_9_22_real;
  reg        [17:0]   img_reg_array_9_22_imag;
  reg        [17:0]   img_reg_array_9_23_real;
  reg        [17:0]   img_reg_array_9_23_imag;
  reg        [17:0]   img_reg_array_9_24_real;
  reg        [17:0]   img_reg_array_9_24_imag;
  reg        [17:0]   img_reg_array_9_25_real;
  reg        [17:0]   img_reg_array_9_25_imag;
  reg        [17:0]   img_reg_array_9_26_real;
  reg        [17:0]   img_reg_array_9_26_imag;
  reg        [17:0]   img_reg_array_9_27_real;
  reg        [17:0]   img_reg_array_9_27_imag;
  reg        [17:0]   img_reg_array_9_28_real;
  reg        [17:0]   img_reg_array_9_28_imag;
  reg        [17:0]   img_reg_array_9_29_real;
  reg        [17:0]   img_reg_array_9_29_imag;
  reg        [17:0]   img_reg_array_9_30_real;
  reg        [17:0]   img_reg_array_9_30_imag;
  reg        [17:0]   img_reg_array_9_31_real;
  reg        [17:0]   img_reg_array_9_31_imag;
  reg        [17:0]   img_reg_array_9_32_real;
  reg        [17:0]   img_reg_array_9_32_imag;
  reg        [17:0]   img_reg_array_9_33_real;
  reg        [17:0]   img_reg_array_9_33_imag;
  reg        [17:0]   img_reg_array_9_34_real;
  reg        [17:0]   img_reg_array_9_34_imag;
  reg        [17:0]   img_reg_array_9_35_real;
  reg        [17:0]   img_reg_array_9_35_imag;
  reg        [17:0]   img_reg_array_9_36_real;
  reg        [17:0]   img_reg_array_9_36_imag;
  reg        [17:0]   img_reg_array_9_37_real;
  reg        [17:0]   img_reg_array_9_37_imag;
  reg        [17:0]   img_reg_array_9_38_real;
  reg        [17:0]   img_reg_array_9_38_imag;
  reg        [17:0]   img_reg_array_9_39_real;
  reg        [17:0]   img_reg_array_9_39_imag;
  reg        [17:0]   img_reg_array_9_40_real;
  reg        [17:0]   img_reg_array_9_40_imag;
  reg        [17:0]   img_reg_array_9_41_real;
  reg        [17:0]   img_reg_array_9_41_imag;
  reg        [17:0]   img_reg_array_9_42_real;
  reg        [17:0]   img_reg_array_9_42_imag;
  reg        [17:0]   img_reg_array_9_43_real;
  reg        [17:0]   img_reg_array_9_43_imag;
  reg        [17:0]   img_reg_array_9_44_real;
  reg        [17:0]   img_reg_array_9_44_imag;
  reg        [17:0]   img_reg_array_9_45_real;
  reg        [17:0]   img_reg_array_9_45_imag;
  reg        [17:0]   img_reg_array_9_46_real;
  reg        [17:0]   img_reg_array_9_46_imag;
  reg        [17:0]   img_reg_array_9_47_real;
  reg        [17:0]   img_reg_array_9_47_imag;
  reg        [17:0]   img_reg_array_9_48_real;
  reg        [17:0]   img_reg_array_9_48_imag;
  reg        [17:0]   img_reg_array_9_49_real;
  reg        [17:0]   img_reg_array_9_49_imag;
  reg        [17:0]   img_reg_array_9_50_real;
  reg        [17:0]   img_reg_array_9_50_imag;
  reg        [17:0]   img_reg_array_9_51_real;
  reg        [17:0]   img_reg_array_9_51_imag;
  reg        [17:0]   img_reg_array_9_52_real;
  reg        [17:0]   img_reg_array_9_52_imag;
  reg        [17:0]   img_reg_array_9_53_real;
  reg        [17:0]   img_reg_array_9_53_imag;
  reg        [17:0]   img_reg_array_9_54_real;
  reg        [17:0]   img_reg_array_9_54_imag;
  reg        [17:0]   img_reg_array_9_55_real;
  reg        [17:0]   img_reg_array_9_55_imag;
  reg        [17:0]   img_reg_array_9_56_real;
  reg        [17:0]   img_reg_array_9_56_imag;
  reg        [17:0]   img_reg_array_9_57_real;
  reg        [17:0]   img_reg_array_9_57_imag;
  reg        [17:0]   img_reg_array_9_58_real;
  reg        [17:0]   img_reg_array_9_58_imag;
  reg        [17:0]   img_reg_array_9_59_real;
  reg        [17:0]   img_reg_array_9_59_imag;
  reg        [17:0]   img_reg_array_9_60_real;
  reg        [17:0]   img_reg_array_9_60_imag;
  reg        [17:0]   img_reg_array_9_61_real;
  reg        [17:0]   img_reg_array_9_61_imag;
  reg        [17:0]   img_reg_array_9_62_real;
  reg        [17:0]   img_reg_array_9_62_imag;
  reg        [17:0]   img_reg_array_9_63_real;
  reg        [17:0]   img_reg_array_9_63_imag;
  reg        [17:0]   img_reg_array_10_0_real;
  reg        [17:0]   img_reg_array_10_0_imag;
  reg        [17:0]   img_reg_array_10_1_real;
  reg        [17:0]   img_reg_array_10_1_imag;
  reg        [17:0]   img_reg_array_10_2_real;
  reg        [17:0]   img_reg_array_10_2_imag;
  reg        [17:0]   img_reg_array_10_3_real;
  reg        [17:0]   img_reg_array_10_3_imag;
  reg        [17:0]   img_reg_array_10_4_real;
  reg        [17:0]   img_reg_array_10_4_imag;
  reg        [17:0]   img_reg_array_10_5_real;
  reg        [17:0]   img_reg_array_10_5_imag;
  reg        [17:0]   img_reg_array_10_6_real;
  reg        [17:0]   img_reg_array_10_6_imag;
  reg        [17:0]   img_reg_array_10_7_real;
  reg        [17:0]   img_reg_array_10_7_imag;
  reg        [17:0]   img_reg_array_10_8_real;
  reg        [17:0]   img_reg_array_10_8_imag;
  reg        [17:0]   img_reg_array_10_9_real;
  reg        [17:0]   img_reg_array_10_9_imag;
  reg        [17:0]   img_reg_array_10_10_real;
  reg        [17:0]   img_reg_array_10_10_imag;
  reg        [17:0]   img_reg_array_10_11_real;
  reg        [17:0]   img_reg_array_10_11_imag;
  reg        [17:0]   img_reg_array_10_12_real;
  reg        [17:0]   img_reg_array_10_12_imag;
  reg        [17:0]   img_reg_array_10_13_real;
  reg        [17:0]   img_reg_array_10_13_imag;
  reg        [17:0]   img_reg_array_10_14_real;
  reg        [17:0]   img_reg_array_10_14_imag;
  reg        [17:0]   img_reg_array_10_15_real;
  reg        [17:0]   img_reg_array_10_15_imag;
  reg        [17:0]   img_reg_array_10_16_real;
  reg        [17:0]   img_reg_array_10_16_imag;
  reg        [17:0]   img_reg_array_10_17_real;
  reg        [17:0]   img_reg_array_10_17_imag;
  reg        [17:0]   img_reg_array_10_18_real;
  reg        [17:0]   img_reg_array_10_18_imag;
  reg        [17:0]   img_reg_array_10_19_real;
  reg        [17:0]   img_reg_array_10_19_imag;
  reg        [17:0]   img_reg_array_10_20_real;
  reg        [17:0]   img_reg_array_10_20_imag;
  reg        [17:0]   img_reg_array_10_21_real;
  reg        [17:0]   img_reg_array_10_21_imag;
  reg        [17:0]   img_reg_array_10_22_real;
  reg        [17:0]   img_reg_array_10_22_imag;
  reg        [17:0]   img_reg_array_10_23_real;
  reg        [17:0]   img_reg_array_10_23_imag;
  reg        [17:0]   img_reg_array_10_24_real;
  reg        [17:0]   img_reg_array_10_24_imag;
  reg        [17:0]   img_reg_array_10_25_real;
  reg        [17:0]   img_reg_array_10_25_imag;
  reg        [17:0]   img_reg_array_10_26_real;
  reg        [17:0]   img_reg_array_10_26_imag;
  reg        [17:0]   img_reg_array_10_27_real;
  reg        [17:0]   img_reg_array_10_27_imag;
  reg        [17:0]   img_reg_array_10_28_real;
  reg        [17:0]   img_reg_array_10_28_imag;
  reg        [17:0]   img_reg_array_10_29_real;
  reg        [17:0]   img_reg_array_10_29_imag;
  reg        [17:0]   img_reg_array_10_30_real;
  reg        [17:0]   img_reg_array_10_30_imag;
  reg        [17:0]   img_reg_array_10_31_real;
  reg        [17:0]   img_reg_array_10_31_imag;
  reg        [17:0]   img_reg_array_10_32_real;
  reg        [17:0]   img_reg_array_10_32_imag;
  reg        [17:0]   img_reg_array_10_33_real;
  reg        [17:0]   img_reg_array_10_33_imag;
  reg        [17:0]   img_reg_array_10_34_real;
  reg        [17:0]   img_reg_array_10_34_imag;
  reg        [17:0]   img_reg_array_10_35_real;
  reg        [17:0]   img_reg_array_10_35_imag;
  reg        [17:0]   img_reg_array_10_36_real;
  reg        [17:0]   img_reg_array_10_36_imag;
  reg        [17:0]   img_reg_array_10_37_real;
  reg        [17:0]   img_reg_array_10_37_imag;
  reg        [17:0]   img_reg_array_10_38_real;
  reg        [17:0]   img_reg_array_10_38_imag;
  reg        [17:0]   img_reg_array_10_39_real;
  reg        [17:0]   img_reg_array_10_39_imag;
  reg        [17:0]   img_reg_array_10_40_real;
  reg        [17:0]   img_reg_array_10_40_imag;
  reg        [17:0]   img_reg_array_10_41_real;
  reg        [17:0]   img_reg_array_10_41_imag;
  reg        [17:0]   img_reg_array_10_42_real;
  reg        [17:0]   img_reg_array_10_42_imag;
  reg        [17:0]   img_reg_array_10_43_real;
  reg        [17:0]   img_reg_array_10_43_imag;
  reg        [17:0]   img_reg_array_10_44_real;
  reg        [17:0]   img_reg_array_10_44_imag;
  reg        [17:0]   img_reg_array_10_45_real;
  reg        [17:0]   img_reg_array_10_45_imag;
  reg        [17:0]   img_reg_array_10_46_real;
  reg        [17:0]   img_reg_array_10_46_imag;
  reg        [17:0]   img_reg_array_10_47_real;
  reg        [17:0]   img_reg_array_10_47_imag;
  reg        [17:0]   img_reg_array_10_48_real;
  reg        [17:0]   img_reg_array_10_48_imag;
  reg        [17:0]   img_reg_array_10_49_real;
  reg        [17:0]   img_reg_array_10_49_imag;
  reg        [17:0]   img_reg_array_10_50_real;
  reg        [17:0]   img_reg_array_10_50_imag;
  reg        [17:0]   img_reg_array_10_51_real;
  reg        [17:0]   img_reg_array_10_51_imag;
  reg        [17:0]   img_reg_array_10_52_real;
  reg        [17:0]   img_reg_array_10_52_imag;
  reg        [17:0]   img_reg_array_10_53_real;
  reg        [17:0]   img_reg_array_10_53_imag;
  reg        [17:0]   img_reg_array_10_54_real;
  reg        [17:0]   img_reg_array_10_54_imag;
  reg        [17:0]   img_reg_array_10_55_real;
  reg        [17:0]   img_reg_array_10_55_imag;
  reg        [17:0]   img_reg_array_10_56_real;
  reg        [17:0]   img_reg_array_10_56_imag;
  reg        [17:0]   img_reg_array_10_57_real;
  reg        [17:0]   img_reg_array_10_57_imag;
  reg        [17:0]   img_reg_array_10_58_real;
  reg        [17:0]   img_reg_array_10_58_imag;
  reg        [17:0]   img_reg_array_10_59_real;
  reg        [17:0]   img_reg_array_10_59_imag;
  reg        [17:0]   img_reg_array_10_60_real;
  reg        [17:0]   img_reg_array_10_60_imag;
  reg        [17:0]   img_reg_array_10_61_real;
  reg        [17:0]   img_reg_array_10_61_imag;
  reg        [17:0]   img_reg_array_10_62_real;
  reg        [17:0]   img_reg_array_10_62_imag;
  reg        [17:0]   img_reg_array_10_63_real;
  reg        [17:0]   img_reg_array_10_63_imag;
  reg        [17:0]   img_reg_array_11_0_real;
  reg        [17:0]   img_reg_array_11_0_imag;
  reg        [17:0]   img_reg_array_11_1_real;
  reg        [17:0]   img_reg_array_11_1_imag;
  reg        [17:0]   img_reg_array_11_2_real;
  reg        [17:0]   img_reg_array_11_2_imag;
  reg        [17:0]   img_reg_array_11_3_real;
  reg        [17:0]   img_reg_array_11_3_imag;
  reg        [17:0]   img_reg_array_11_4_real;
  reg        [17:0]   img_reg_array_11_4_imag;
  reg        [17:0]   img_reg_array_11_5_real;
  reg        [17:0]   img_reg_array_11_5_imag;
  reg        [17:0]   img_reg_array_11_6_real;
  reg        [17:0]   img_reg_array_11_6_imag;
  reg        [17:0]   img_reg_array_11_7_real;
  reg        [17:0]   img_reg_array_11_7_imag;
  reg        [17:0]   img_reg_array_11_8_real;
  reg        [17:0]   img_reg_array_11_8_imag;
  reg        [17:0]   img_reg_array_11_9_real;
  reg        [17:0]   img_reg_array_11_9_imag;
  reg        [17:0]   img_reg_array_11_10_real;
  reg        [17:0]   img_reg_array_11_10_imag;
  reg        [17:0]   img_reg_array_11_11_real;
  reg        [17:0]   img_reg_array_11_11_imag;
  reg        [17:0]   img_reg_array_11_12_real;
  reg        [17:0]   img_reg_array_11_12_imag;
  reg        [17:0]   img_reg_array_11_13_real;
  reg        [17:0]   img_reg_array_11_13_imag;
  reg        [17:0]   img_reg_array_11_14_real;
  reg        [17:0]   img_reg_array_11_14_imag;
  reg        [17:0]   img_reg_array_11_15_real;
  reg        [17:0]   img_reg_array_11_15_imag;
  reg        [17:0]   img_reg_array_11_16_real;
  reg        [17:0]   img_reg_array_11_16_imag;
  reg        [17:0]   img_reg_array_11_17_real;
  reg        [17:0]   img_reg_array_11_17_imag;
  reg        [17:0]   img_reg_array_11_18_real;
  reg        [17:0]   img_reg_array_11_18_imag;
  reg        [17:0]   img_reg_array_11_19_real;
  reg        [17:0]   img_reg_array_11_19_imag;
  reg        [17:0]   img_reg_array_11_20_real;
  reg        [17:0]   img_reg_array_11_20_imag;
  reg        [17:0]   img_reg_array_11_21_real;
  reg        [17:0]   img_reg_array_11_21_imag;
  reg        [17:0]   img_reg_array_11_22_real;
  reg        [17:0]   img_reg_array_11_22_imag;
  reg        [17:0]   img_reg_array_11_23_real;
  reg        [17:0]   img_reg_array_11_23_imag;
  reg        [17:0]   img_reg_array_11_24_real;
  reg        [17:0]   img_reg_array_11_24_imag;
  reg        [17:0]   img_reg_array_11_25_real;
  reg        [17:0]   img_reg_array_11_25_imag;
  reg        [17:0]   img_reg_array_11_26_real;
  reg        [17:0]   img_reg_array_11_26_imag;
  reg        [17:0]   img_reg_array_11_27_real;
  reg        [17:0]   img_reg_array_11_27_imag;
  reg        [17:0]   img_reg_array_11_28_real;
  reg        [17:0]   img_reg_array_11_28_imag;
  reg        [17:0]   img_reg_array_11_29_real;
  reg        [17:0]   img_reg_array_11_29_imag;
  reg        [17:0]   img_reg_array_11_30_real;
  reg        [17:0]   img_reg_array_11_30_imag;
  reg        [17:0]   img_reg_array_11_31_real;
  reg        [17:0]   img_reg_array_11_31_imag;
  reg        [17:0]   img_reg_array_11_32_real;
  reg        [17:0]   img_reg_array_11_32_imag;
  reg        [17:0]   img_reg_array_11_33_real;
  reg        [17:0]   img_reg_array_11_33_imag;
  reg        [17:0]   img_reg_array_11_34_real;
  reg        [17:0]   img_reg_array_11_34_imag;
  reg        [17:0]   img_reg_array_11_35_real;
  reg        [17:0]   img_reg_array_11_35_imag;
  reg        [17:0]   img_reg_array_11_36_real;
  reg        [17:0]   img_reg_array_11_36_imag;
  reg        [17:0]   img_reg_array_11_37_real;
  reg        [17:0]   img_reg_array_11_37_imag;
  reg        [17:0]   img_reg_array_11_38_real;
  reg        [17:0]   img_reg_array_11_38_imag;
  reg        [17:0]   img_reg_array_11_39_real;
  reg        [17:0]   img_reg_array_11_39_imag;
  reg        [17:0]   img_reg_array_11_40_real;
  reg        [17:0]   img_reg_array_11_40_imag;
  reg        [17:0]   img_reg_array_11_41_real;
  reg        [17:0]   img_reg_array_11_41_imag;
  reg        [17:0]   img_reg_array_11_42_real;
  reg        [17:0]   img_reg_array_11_42_imag;
  reg        [17:0]   img_reg_array_11_43_real;
  reg        [17:0]   img_reg_array_11_43_imag;
  reg        [17:0]   img_reg_array_11_44_real;
  reg        [17:0]   img_reg_array_11_44_imag;
  reg        [17:0]   img_reg_array_11_45_real;
  reg        [17:0]   img_reg_array_11_45_imag;
  reg        [17:0]   img_reg_array_11_46_real;
  reg        [17:0]   img_reg_array_11_46_imag;
  reg        [17:0]   img_reg_array_11_47_real;
  reg        [17:0]   img_reg_array_11_47_imag;
  reg        [17:0]   img_reg_array_11_48_real;
  reg        [17:0]   img_reg_array_11_48_imag;
  reg        [17:0]   img_reg_array_11_49_real;
  reg        [17:0]   img_reg_array_11_49_imag;
  reg        [17:0]   img_reg_array_11_50_real;
  reg        [17:0]   img_reg_array_11_50_imag;
  reg        [17:0]   img_reg_array_11_51_real;
  reg        [17:0]   img_reg_array_11_51_imag;
  reg        [17:0]   img_reg_array_11_52_real;
  reg        [17:0]   img_reg_array_11_52_imag;
  reg        [17:0]   img_reg_array_11_53_real;
  reg        [17:0]   img_reg_array_11_53_imag;
  reg        [17:0]   img_reg_array_11_54_real;
  reg        [17:0]   img_reg_array_11_54_imag;
  reg        [17:0]   img_reg_array_11_55_real;
  reg        [17:0]   img_reg_array_11_55_imag;
  reg        [17:0]   img_reg_array_11_56_real;
  reg        [17:0]   img_reg_array_11_56_imag;
  reg        [17:0]   img_reg_array_11_57_real;
  reg        [17:0]   img_reg_array_11_57_imag;
  reg        [17:0]   img_reg_array_11_58_real;
  reg        [17:0]   img_reg_array_11_58_imag;
  reg        [17:0]   img_reg_array_11_59_real;
  reg        [17:0]   img_reg_array_11_59_imag;
  reg        [17:0]   img_reg_array_11_60_real;
  reg        [17:0]   img_reg_array_11_60_imag;
  reg        [17:0]   img_reg_array_11_61_real;
  reg        [17:0]   img_reg_array_11_61_imag;
  reg        [17:0]   img_reg_array_11_62_real;
  reg        [17:0]   img_reg_array_11_62_imag;
  reg        [17:0]   img_reg_array_11_63_real;
  reg        [17:0]   img_reg_array_11_63_imag;
  reg        [17:0]   img_reg_array_12_0_real;
  reg        [17:0]   img_reg_array_12_0_imag;
  reg        [17:0]   img_reg_array_12_1_real;
  reg        [17:0]   img_reg_array_12_1_imag;
  reg        [17:0]   img_reg_array_12_2_real;
  reg        [17:0]   img_reg_array_12_2_imag;
  reg        [17:0]   img_reg_array_12_3_real;
  reg        [17:0]   img_reg_array_12_3_imag;
  reg        [17:0]   img_reg_array_12_4_real;
  reg        [17:0]   img_reg_array_12_4_imag;
  reg        [17:0]   img_reg_array_12_5_real;
  reg        [17:0]   img_reg_array_12_5_imag;
  reg        [17:0]   img_reg_array_12_6_real;
  reg        [17:0]   img_reg_array_12_6_imag;
  reg        [17:0]   img_reg_array_12_7_real;
  reg        [17:0]   img_reg_array_12_7_imag;
  reg        [17:0]   img_reg_array_12_8_real;
  reg        [17:0]   img_reg_array_12_8_imag;
  reg        [17:0]   img_reg_array_12_9_real;
  reg        [17:0]   img_reg_array_12_9_imag;
  reg        [17:0]   img_reg_array_12_10_real;
  reg        [17:0]   img_reg_array_12_10_imag;
  reg        [17:0]   img_reg_array_12_11_real;
  reg        [17:0]   img_reg_array_12_11_imag;
  reg        [17:0]   img_reg_array_12_12_real;
  reg        [17:0]   img_reg_array_12_12_imag;
  reg        [17:0]   img_reg_array_12_13_real;
  reg        [17:0]   img_reg_array_12_13_imag;
  reg        [17:0]   img_reg_array_12_14_real;
  reg        [17:0]   img_reg_array_12_14_imag;
  reg        [17:0]   img_reg_array_12_15_real;
  reg        [17:0]   img_reg_array_12_15_imag;
  reg        [17:0]   img_reg_array_12_16_real;
  reg        [17:0]   img_reg_array_12_16_imag;
  reg        [17:0]   img_reg_array_12_17_real;
  reg        [17:0]   img_reg_array_12_17_imag;
  reg        [17:0]   img_reg_array_12_18_real;
  reg        [17:0]   img_reg_array_12_18_imag;
  reg        [17:0]   img_reg_array_12_19_real;
  reg        [17:0]   img_reg_array_12_19_imag;
  reg        [17:0]   img_reg_array_12_20_real;
  reg        [17:0]   img_reg_array_12_20_imag;
  reg        [17:0]   img_reg_array_12_21_real;
  reg        [17:0]   img_reg_array_12_21_imag;
  reg        [17:0]   img_reg_array_12_22_real;
  reg        [17:0]   img_reg_array_12_22_imag;
  reg        [17:0]   img_reg_array_12_23_real;
  reg        [17:0]   img_reg_array_12_23_imag;
  reg        [17:0]   img_reg_array_12_24_real;
  reg        [17:0]   img_reg_array_12_24_imag;
  reg        [17:0]   img_reg_array_12_25_real;
  reg        [17:0]   img_reg_array_12_25_imag;
  reg        [17:0]   img_reg_array_12_26_real;
  reg        [17:0]   img_reg_array_12_26_imag;
  reg        [17:0]   img_reg_array_12_27_real;
  reg        [17:0]   img_reg_array_12_27_imag;
  reg        [17:0]   img_reg_array_12_28_real;
  reg        [17:0]   img_reg_array_12_28_imag;
  reg        [17:0]   img_reg_array_12_29_real;
  reg        [17:0]   img_reg_array_12_29_imag;
  reg        [17:0]   img_reg_array_12_30_real;
  reg        [17:0]   img_reg_array_12_30_imag;
  reg        [17:0]   img_reg_array_12_31_real;
  reg        [17:0]   img_reg_array_12_31_imag;
  reg        [17:0]   img_reg_array_12_32_real;
  reg        [17:0]   img_reg_array_12_32_imag;
  reg        [17:0]   img_reg_array_12_33_real;
  reg        [17:0]   img_reg_array_12_33_imag;
  reg        [17:0]   img_reg_array_12_34_real;
  reg        [17:0]   img_reg_array_12_34_imag;
  reg        [17:0]   img_reg_array_12_35_real;
  reg        [17:0]   img_reg_array_12_35_imag;
  reg        [17:0]   img_reg_array_12_36_real;
  reg        [17:0]   img_reg_array_12_36_imag;
  reg        [17:0]   img_reg_array_12_37_real;
  reg        [17:0]   img_reg_array_12_37_imag;
  reg        [17:0]   img_reg_array_12_38_real;
  reg        [17:0]   img_reg_array_12_38_imag;
  reg        [17:0]   img_reg_array_12_39_real;
  reg        [17:0]   img_reg_array_12_39_imag;
  reg        [17:0]   img_reg_array_12_40_real;
  reg        [17:0]   img_reg_array_12_40_imag;
  reg        [17:0]   img_reg_array_12_41_real;
  reg        [17:0]   img_reg_array_12_41_imag;
  reg        [17:0]   img_reg_array_12_42_real;
  reg        [17:0]   img_reg_array_12_42_imag;
  reg        [17:0]   img_reg_array_12_43_real;
  reg        [17:0]   img_reg_array_12_43_imag;
  reg        [17:0]   img_reg_array_12_44_real;
  reg        [17:0]   img_reg_array_12_44_imag;
  reg        [17:0]   img_reg_array_12_45_real;
  reg        [17:0]   img_reg_array_12_45_imag;
  reg        [17:0]   img_reg_array_12_46_real;
  reg        [17:0]   img_reg_array_12_46_imag;
  reg        [17:0]   img_reg_array_12_47_real;
  reg        [17:0]   img_reg_array_12_47_imag;
  reg        [17:0]   img_reg_array_12_48_real;
  reg        [17:0]   img_reg_array_12_48_imag;
  reg        [17:0]   img_reg_array_12_49_real;
  reg        [17:0]   img_reg_array_12_49_imag;
  reg        [17:0]   img_reg_array_12_50_real;
  reg        [17:0]   img_reg_array_12_50_imag;
  reg        [17:0]   img_reg_array_12_51_real;
  reg        [17:0]   img_reg_array_12_51_imag;
  reg        [17:0]   img_reg_array_12_52_real;
  reg        [17:0]   img_reg_array_12_52_imag;
  reg        [17:0]   img_reg_array_12_53_real;
  reg        [17:0]   img_reg_array_12_53_imag;
  reg        [17:0]   img_reg_array_12_54_real;
  reg        [17:0]   img_reg_array_12_54_imag;
  reg        [17:0]   img_reg_array_12_55_real;
  reg        [17:0]   img_reg_array_12_55_imag;
  reg        [17:0]   img_reg_array_12_56_real;
  reg        [17:0]   img_reg_array_12_56_imag;
  reg        [17:0]   img_reg_array_12_57_real;
  reg        [17:0]   img_reg_array_12_57_imag;
  reg        [17:0]   img_reg_array_12_58_real;
  reg        [17:0]   img_reg_array_12_58_imag;
  reg        [17:0]   img_reg_array_12_59_real;
  reg        [17:0]   img_reg_array_12_59_imag;
  reg        [17:0]   img_reg_array_12_60_real;
  reg        [17:0]   img_reg_array_12_60_imag;
  reg        [17:0]   img_reg_array_12_61_real;
  reg        [17:0]   img_reg_array_12_61_imag;
  reg        [17:0]   img_reg_array_12_62_real;
  reg        [17:0]   img_reg_array_12_62_imag;
  reg        [17:0]   img_reg_array_12_63_real;
  reg        [17:0]   img_reg_array_12_63_imag;
  reg        [17:0]   img_reg_array_13_0_real;
  reg        [17:0]   img_reg_array_13_0_imag;
  reg        [17:0]   img_reg_array_13_1_real;
  reg        [17:0]   img_reg_array_13_1_imag;
  reg        [17:0]   img_reg_array_13_2_real;
  reg        [17:0]   img_reg_array_13_2_imag;
  reg        [17:0]   img_reg_array_13_3_real;
  reg        [17:0]   img_reg_array_13_3_imag;
  reg        [17:0]   img_reg_array_13_4_real;
  reg        [17:0]   img_reg_array_13_4_imag;
  reg        [17:0]   img_reg_array_13_5_real;
  reg        [17:0]   img_reg_array_13_5_imag;
  reg        [17:0]   img_reg_array_13_6_real;
  reg        [17:0]   img_reg_array_13_6_imag;
  reg        [17:0]   img_reg_array_13_7_real;
  reg        [17:0]   img_reg_array_13_7_imag;
  reg        [17:0]   img_reg_array_13_8_real;
  reg        [17:0]   img_reg_array_13_8_imag;
  reg        [17:0]   img_reg_array_13_9_real;
  reg        [17:0]   img_reg_array_13_9_imag;
  reg        [17:0]   img_reg_array_13_10_real;
  reg        [17:0]   img_reg_array_13_10_imag;
  reg        [17:0]   img_reg_array_13_11_real;
  reg        [17:0]   img_reg_array_13_11_imag;
  reg        [17:0]   img_reg_array_13_12_real;
  reg        [17:0]   img_reg_array_13_12_imag;
  reg        [17:0]   img_reg_array_13_13_real;
  reg        [17:0]   img_reg_array_13_13_imag;
  reg        [17:0]   img_reg_array_13_14_real;
  reg        [17:0]   img_reg_array_13_14_imag;
  reg        [17:0]   img_reg_array_13_15_real;
  reg        [17:0]   img_reg_array_13_15_imag;
  reg        [17:0]   img_reg_array_13_16_real;
  reg        [17:0]   img_reg_array_13_16_imag;
  reg        [17:0]   img_reg_array_13_17_real;
  reg        [17:0]   img_reg_array_13_17_imag;
  reg        [17:0]   img_reg_array_13_18_real;
  reg        [17:0]   img_reg_array_13_18_imag;
  reg        [17:0]   img_reg_array_13_19_real;
  reg        [17:0]   img_reg_array_13_19_imag;
  reg        [17:0]   img_reg_array_13_20_real;
  reg        [17:0]   img_reg_array_13_20_imag;
  reg        [17:0]   img_reg_array_13_21_real;
  reg        [17:0]   img_reg_array_13_21_imag;
  reg        [17:0]   img_reg_array_13_22_real;
  reg        [17:0]   img_reg_array_13_22_imag;
  reg        [17:0]   img_reg_array_13_23_real;
  reg        [17:0]   img_reg_array_13_23_imag;
  reg        [17:0]   img_reg_array_13_24_real;
  reg        [17:0]   img_reg_array_13_24_imag;
  reg        [17:0]   img_reg_array_13_25_real;
  reg        [17:0]   img_reg_array_13_25_imag;
  reg        [17:0]   img_reg_array_13_26_real;
  reg        [17:0]   img_reg_array_13_26_imag;
  reg        [17:0]   img_reg_array_13_27_real;
  reg        [17:0]   img_reg_array_13_27_imag;
  reg        [17:0]   img_reg_array_13_28_real;
  reg        [17:0]   img_reg_array_13_28_imag;
  reg        [17:0]   img_reg_array_13_29_real;
  reg        [17:0]   img_reg_array_13_29_imag;
  reg        [17:0]   img_reg_array_13_30_real;
  reg        [17:0]   img_reg_array_13_30_imag;
  reg        [17:0]   img_reg_array_13_31_real;
  reg        [17:0]   img_reg_array_13_31_imag;
  reg        [17:0]   img_reg_array_13_32_real;
  reg        [17:0]   img_reg_array_13_32_imag;
  reg        [17:0]   img_reg_array_13_33_real;
  reg        [17:0]   img_reg_array_13_33_imag;
  reg        [17:0]   img_reg_array_13_34_real;
  reg        [17:0]   img_reg_array_13_34_imag;
  reg        [17:0]   img_reg_array_13_35_real;
  reg        [17:0]   img_reg_array_13_35_imag;
  reg        [17:0]   img_reg_array_13_36_real;
  reg        [17:0]   img_reg_array_13_36_imag;
  reg        [17:0]   img_reg_array_13_37_real;
  reg        [17:0]   img_reg_array_13_37_imag;
  reg        [17:0]   img_reg_array_13_38_real;
  reg        [17:0]   img_reg_array_13_38_imag;
  reg        [17:0]   img_reg_array_13_39_real;
  reg        [17:0]   img_reg_array_13_39_imag;
  reg        [17:0]   img_reg_array_13_40_real;
  reg        [17:0]   img_reg_array_13_40_imag;
  reg        [17:0]   img_reg_array_13_41_real;
  reg        [17:0]   img_reg_array_13_41_imag;
  reg        [17:0]   img_reg_array_13_42_real;
  reg        [17:0]   img_reg_array_13_42_imag;
  reg        [17:0]   img_reg_array_13_43_real;
  reg        [17:0]   img_reg_array_13_43_imag;
  reg        [17:0]   img_reg_array_13_44_real;
  reg        [17:0]   img_reg_array_13_44_imag;
  reg        [17:0]   img_reg_array_13_45_real;
  reg        [17:0]   img_reg_array_13_45_imag;
  reg        [17:0]   img_reg_array_13_46_real;
  reg        [17:0]   img_reg_array_13_46_imag;
  reg        [17:0]   img_reg_array_13_47_real;
  reg        [17:0]   img_reg_array_13_47_imag;
  reg        [17:0]   img_reg_array_13_48_real;
  reg        [17:0]   img_reg_array_13_48_imag;
  reg        [17:0]   img_reg_array_13_49_real;
  reg        [17:0]   img_reg_array_13_49_imag;
  reg        [17:0]   img_reg_array_13_50_real;
  reg        [17:0]   img_reg_array_13_50_imag;
  reg        [17:0]   img_reg_array_13_51_real;
  reg        [17:0]   img_reg_array_13_51_imag;
  reg        [17:0]   img_reg_array_13_52_real;
  reg        [17:0]   img_reg_array_13_52_imag;
  reg        [17:0]   img_reg_array_13_53_real;
  reg        [17:0]   img_reg_array_13_53_imag;
  reg        [17:0]   img_reg_array_13_54_real;
  reg        [17:0]   img_reg_array_13_54_imag;
  reg        [17:0]   img_reg_array_13_55_real;
  reg        [17:0]   img_reg_array_13_55_imag;
  reg        [17:0]   img_reg_array_13_56_real;
  reg        [17:0]   img_reg_array_13_56_imag;
  reg        [17:0]   img_reg_array_13_57_real;
  reg        [17:0]   img_reg_array_13_57_imag;
  reg        [17:0]   img_reg_array_13_58_real;
  reg        [17:0]   img_reg_array_13_58_imag;
  reg        [17:0]   img_reg_array_13_59_real;
  reg        [17:0]   img_reg_array_13_59_imag;
  reg        [17:0]   img_reg_array_13_60_real;
  reg        [17:0]   img_reg_array_13_60_imag;
  reg        [17:0]   img_reg_array_13_61_real;
  reg        [17:0]   img_reg_array_13_61_imag;
  reg        [17:0]   img_reg_array_13_62_real;
  reg        [17:0]   img_reg_array_13_62_imag;
  reg        [17:0]   img_reg_array_13_63_real;
  reg        [17:0]   img_reg_array_13_63_imag;
  reg        [17:0]   img_reg_array_14_0_real;
  reg        [17:0]   img_reg_array_14_0_imag;
  reg        [17:0]   img_reg_array_14_1_real;
  reg        [17:0]   img_reg_array_14_1_imag;
  reg        [17:0]   img_reg_array_14_2_real;
  reg        [17:0]   img_reg_array_14_2_imag;
  reg        [17:0]   img_reg_array_14_3_real;
  reg        [17:0]   img_reg_array_14_3_imag;
  reg        [17:0]   img_reg_array_14_4_real;
  reg        [17:0]   img_reg_array_14_4_imag;
  reg        [17:0]   img_reg_array_14_5_real;
  reg        [17:0]   img_reg_array_14_5_imag;
  reg        [17:0]   img_reg_array_14_6_real;
  reg        [17:0]   img_reg_array_14_6_imag;
  reg        [17:0]   img_reg_array_14_7_real;
  reg        [17:0]   img_reg_array_14_7_imag;
  reg        [17:0]   img_reg_array_14_8_real;
  reg        [17:0]   img_reg_array_14_8_imag;
  reg        [17:0]   img_reg_array_14_9_real;
  reg        [17:0]   img_reg_array_14_9_imag;
  reg        [17:0]   img_reg_array_14_10_real;
  reg        [17:0]   img_reg_array_14_10_imag;
  reg        [17:0]   img_reg_array_14_11_real;
  reg        [17:0]   img_reg_array_14_11_imag;
  reg        [17:0]   img_reg_array_14_12_real;
  reg        [17:0]   img_reg_array_14_12_imag;
  reg        [17:0]   img_reg_array_14_13_real;
  reg        [17:0]   img_reg_array_14_13_imag;
  reg        [17:0]   img_reg_array_14_14_real;
  reg        [17:0]   img_reg_array_14_14_imag;
  reg        [17:0]   img_reg_array_14_15_real;
  reg        [17:0]   img_reg_array_14_15_imag;
  reg        [17:0]   img_reg_array_14_16_real;
  reg        [17:0]   img_reg_array_14_16_imag;
  reg        [17:0]   img_reg_array_14_17_real;
  reg        [17:0]   img_reg_array_14_17_imag;
  reg        [17:0]   img_reg_array_14_18_real;
  reg        [17:0]   img_reg_array_14_18_imag;
  reg        [17:0]   img_reg_array_14_19_real;
  reg        [17:0]   img_reg_array_14_19_imag;
  reg        [17:0]   img_reg_array_14_20_real;
  reg        [17:0]   img_reg_array_14_20_imag;
  reg        [17:0]   img_reg_array_14_21_real;
  reg        [17:0]   img_reg_array_14_21_imag;
  reg        [17:0]   img_reg_array_14_22_real;
  reg        [17:0]   img_reg_array_14_22_imag;
  reg        [17:0]   img_reg_array_14_23_real;
  reg        [17:0]   img_reg_array_14_23_imag;
  reg        [17:0]   img_reg_array_14_24_real;
  reg        [17:0]   img_reg_array_14_24_imag;
  reg        [17:0]   img_reg_array_14_25_real;
  reg        [17:0]   img_reg_array_14_25_imag;
  reg        [17:0]   img_reg_array_14_26_real;
  reg        [17:0]   img_reg_array_14_26_imag;
  reg        [17:0]   img_reg_array_14_27_real;
  reg        [17:0]   img_reg_array_14_27_imag;
  reg        [17:0]   img_reg_array_14_28_real;
  reg        [17:0]   img_reg_array_14_28_imag;
  reg        [17:0]   img_reg_array_14_29_real;
  reg        [17:0]   img_reg_array_14_29_imag;
  reg        [17:0]   img_reg_array_14_30_real;
  reg        [17:0]   img_reg_array_14_30_imag;
  reg        [17:0]   img_reg_array_14_31_real;
  reg        [17:0]   img_reg_array_14_31_imag;
  reg        [17:0]   img_reg_array_14_32_real;
  reg        [17:0]   img_reg_array_14_32_imag;
  reg        [17:0]   img_reg_array_14_33_real;
  reg        [17:0]   img_reg_array_14_33_imag;
  reg        [17:0]   img_reg_array_14_34_real;
  reg        [17:0]   img_reg_array_14_34_imag;
  reg        [17:0]   img_reg_array_14_35_real;
  reg        [17:0]   img_reg_array_14_35_imag;
  reg        [17:0]   img_reg_array_14_36_real;
  reg        [17:0]   img_reg_array_14_36_imag;
  reg        [17:0]   img_reg_array_14_37_real;
  reg        [17:0]   img_reg_array_14_37_imag;
  reg        [17:0]   img_reg_array_14_38_real;
  reg        [17:0]   img_reg_array_14_38_imag;
  reg        [17:0]   img_reg_array_14_39_real;
  reg        [17:0]   img_reg_array_14_39_imag;
  reg        [17:0]   img_reg_array_14_40_real;
  reg        [17:0]   img_reg_array_14_40_imag;
  reg        [17:0]   img_reg_array_14_41_real;
  reg        [17:0]   img_reg_array_14_41_imag;
  reg        [17:0]   img_reg_array_14_42_real;
  reg        [17:0]   img_reg_array_14_42_imag;
  reg        [17:0]   img_reg_array_14_43_real;
  reg        [17:0]   img_reg_array_14_43_imag;
  reg        [17:0]   img_reg_array_14_44_real;
  reg        [17:0]   img_reg_array_14_44_imag;
  reg        [17:0]   img_reg_array_14_45_real;
  reg        [17:0]   img_reg_array_14_45_imag;
  reg        [17:0]   img_reg_array_14_46_real;
  reg        [17:0]   img_reg_array_14_46_imag;
  reg        [17:0]   img_reg_array_14_47_real;
  reg        [17:0]   img_reg_array_14_47_imag;
  reg        [17:0]   img_reg_array_14_48_real;
  reg        [17:0]   img_reg_array_14_48_imag;
  reg        [17:0]   img_reg_array_14_49_real;
  reg        [17:0]   img_reg_array_14_49_imag;
  reg        [17:0]   img_reg_array_14_50_real;
  reg        [17:0]   img_reg_array_14_50_imag;
  reg        [17:0]   img_reg_array_14_51_real;
  reg        [17:0]   img_reg_array_14_51_imag;
  reg        [17:0]   img_reg_array_14_52_real;
  reg        [17:0]   img_reg_array_14_52_imag;
  reg        [17:0]   img_reg_array_14_53_real;
  reg        [17:0]   img_reg_array_14_53_imag;
  reg        [17:0]   img_reg_array_14_54_real;
  reg        [17:0]   img_reg_array_14_54_imag;
  reg        [17:0]   img_reg_array_14_55_real;
  reg        [17:0]   img_reg_array_14_55_imag;
  reg        [17:0]   img_reg_array_14_56_real;
  reg        [17:0]   img_reg_array_14_56_imag;
  reg        [17:0]   img_reg_array_14_57_real;
  reg        [17:0]   img_reg_array_14_57_imag;
  reg        [17:0]   img_reg_array_14_58_real;
  reg        [17:0]   img_reg_array_14_58_imag;
  reg        [17:0]   img_reg_array_14_59_real;
  reg        [17:0]   img_reg_array_14_59_imag;
  reg        [17:0]   img_reg_array_14_60_real;
  reg        [17:0]   img_reg_array_14_60_imag;
  reg        [17:0]   img_reg_array_14_61_real;
  reg        [17:0]   img_reg_array_14_61_imag;
  reg        [17:0]   img_reg_array_14_62_real;
  reg        [17:0]   img_reg_array_14_62_imag;
  reg        [17:0]   img_reg_array_14_63_real;
  reg        [17:0]   img_reg_array_14_63_imag;
  reg        [17:0]   img_reg_array_15_0_real;
  reg        [17:0]   img_reg_array_15_0_imag;
  reg        [17:0]   img_reg_array_15_1_real;
  reg        [17:0]   img_reg_array_15_1_imag;
  reg        [17:0]   img_reg_array_15_2_real;
  reg        [17:0]   img_reg_array_15_2_imag;
  reg        [17:0]   img_reg_array_15_3_real;
  reg        [17:0]   img_reg_array_15_3_imag;
  reg        [17:0]   img_reg_array_15_4_real;
  reg        [17:0]   img_reg_array_15_4_imag;
  reg        [17:0]   img_reg_array_15_5_real;
  reg        [17:0]   img_reg_array_15_5_imag;
  reg        [17:0]   img_reg_array_15_6_real;
  reg        [17:0]   img_reg_array_15_6_imag;
  reg        [17:0]   img_reg_array_15_7_real;
  reg        [17:0]   img_reg_array_15_7_imag;
  reg        [17:0]   img_reg_array_15_8_real;
  reg        [17:0]   img_reg_array_15_8_imag;
  reg        [17:0]   img_reg_array_15_9_real;
  reg        [17:0]   img_reg_array_15_9_imag;
  reg        [17:0]   img_reg_array_15_10_real;
  reg        [17:0]   img_reg_array_15_10_imag;
  reg        [17:0]   img_reg_array_15_11_real;
  reg        [17:0]   img_reg_array_15_11_imag;
  reg        [17:0]   img_reg_array_15_12_real;
  reg        [17:0]   img_reg_array_15_12_imag;
  reg        [17:0]   img_reg_array_15_13_real;
  reg        [17:0]   img_reg_array_15_13_imag;
  reg        [17:0]   img_reg_array_15_14_real;
  reg        [17:0]   img_reg_array_15_14_imag;
  reg        [17:0]   img_reg_array_15_15_real;
  reg        [17:0]   img_reg_array_15_15_imag;
  reg        [17:0]   img_reg_array_15_16_real;
  reg        [17:0]   img_reg_array_15_16_imag;
  reg        [17:0]   img_reg_array_15_17_real;
  reg        [17:0]   img_reg_array_15_17_imag;
  reg        [17:0]   img_reg_array_15_18_real;
  reg        [17:0]   img_reg_array_15_18_imag;
  reg        [17:0]   img_reg_array_15_19_real;
  reg        [17:0]   img_reg_array_15_19_imag;
  reg        [17:0]   img_reg_array_15_20_real;
  reg        [17:0]   img_reg_array_15_20_imag;
  reg        [17:0]   img_reg_array_15_21_real;
  reg        [17:0]   img_reg_array_15_21_imag;
  reg        [17:0]   img_reg_array_15_22_real;
  reg        [17:0]   img_reg_array_15_22_imag;
  reg        [17:0]   img_reg_array_15_23_real;
  reg        [17:0]   img_reg_array_15_23_imag;
  reg        [17:0]   img_reg_array_15_24_real;
  reg        [17:0]   img_reg_array_15_24_imag;
  reg        [17:0]   img_reg_array_15_25_real;
  reg        [17:0]   img_reg_array_15_25_imag;
  reg        [17:0]   img_reg_array_15_26_real;
  reg        [17:0]   img_reg_array_15_26_imag;
  reg        [17:0]   img_reg_array_15_27_real;
  reg        [17:0]   img_reg_array_15_27_imag;
  reg        [17:0]   img_reg_array_15_28_real;
  reg        [17:0]   img_reg_array_15_28_imag;
  reg        [17:0]   img_reg_array_15_29_real;
  reg        [17:0]   img_reg_array_15_29_imag;
  reg        [17:0]   img_reg_array_15_30_real;
  reg        [17:0]   img_reg_array_15_30_imag;
  reg        [17:0]   img_reg_array_15_31_real;
  reg        [17:0]   img_reg_array_15_31_imag;
  reg        [17:0]   img_reg_array_15_32_real;
  reg        [17:0]   img_reg_array_15_32_imag;
  reg        [17:0]   img_reg_array_15_33_real;
  reg        [17:0]   img_reg_array_15_33_imag;
  reg        [17:0]   img_reg_array_15_34_real;
  reg        [17:0]   img_reg_array_15_34_imag;
  reg        [17:0]   img_reg_array_15_35_real;
  reg        [17:0]   img_reg_array_15_35_imag;
  reg        [17:0]   img_reg_array_15_36_real;
  reg        [17:0]   img_reg_array_15_36_imag;
  reg        [17:0]   img_reg_array_15_37_real;
  reg        [17:0]   img_reg_array_15_37_imag;
  reg        [17:0]   img_reg_array_15_38_real;
  reg        [17:0]   img_reg_array_15_38_imag;
  reg        [17:0]   img_reg_array_15_39_real;
  reg        [17:0]   img_reg_array_15_39_imag;
  reg        [17:0]   img_reg_array_15_40_real;
  reg        [17:0]   img_reg_array_15_40_imag;
  reg        [17:0]   img_reg_array_15_41_real;
  reg        [17:0]   img_reg_array_15_41_imag;
  reg        [17:0]   img_reg_array_15_42_real;
  reg        [17:0]   img_reg_array_15_42_imag;
  reg        [17:0]   img_reg_array_15_43_real;
  reg        [17:0]   img_reg_array_15_43_imag;
  reg        [17:0]   img_reg_array_15_44_real;
  reg        [17:0]   img_reg_array_15_44_imag;
  reg        [17:0]   img_reg_array_15_45_real;
  reg        [17:0]   img_reg_array_15_45_imag;
  reg        [17:0]   img_reg_array_15_46_real;
  reg        [17:0]   img_reg_array_15_46_imag;
  reg        [17:0]   img_reg_array_15_47_real;
  reg        [17:0]   img_reg_array_15_47_imag;
  reg        [17:0]   img_reg_array_15_48_real;
  reg        [17:0]   img_reg_array_15_48_imag;
  reg        [17:0]   img_reg_array_15_49_real;
  reg        [17:0]   img_reg_array_15_49_imag;
  reg        [17:0]   img_reg_array_15_50_real;
  reg        [17:0]   img_reg_array_15_50_imag;
  reg        [17:0]   img_reg_array_15_51_real;
  reg        [17:0]   img_reg_array_15_51_imag;
  reg        [17:0]   img_reg_array_15_52_real;
  reg        [17:0]   img_reg_array_15_52_imag;
  reg        [17:0]   img_reg_array_15_53_real;
  reg        [17:0]   img_reg_array_15_53_imag;
  reg        [17:0]   img_reg_array_15_54_real;
  reg        [17:0]   img_reg_array_15_54_imag;
  reg        [17:0]   img_reg_array_15_55_real;
  reg        [17:0]   img_reg_array_15_55_imag;
  reg        [17:0]   img_reg_array_15_56_real;
  reg        [17:0]   img_reg_array_15_56_imag;
  reg        [17:0]   img_reg_array_15_57_real;
  reg        [17:0]   img_reg_array_15_57_imag;
  reg        [17:0]   img_reg_array_15_58_real;
  reg        [17:0]   img_reg_array_15_58_imag;
  reg        [17:0]   img_reg_array_15_59_real;
  reg        [17:0]   img_reg_array_15_59_imag;
  reg        [17:0]   img_reg_array_15_60_real;
  reg        [17:0]   img_reg_array_15_60_imag;
  reg        [17:0]   img_reg_array_15_61_real;
  reg        [17:0]   img_reg_array_15_61_imag;
  reg        [17:0]   img_reg_array_15_62_real;
  reg        [17:0]   img_reg_array_15_62_imag;
  reg        [17:0]   img_reg_array_15_63_real;
  reg        [17:0]   img_reg_array_15_63_imag;
  reg        [17:0]   img_reg_array_16_0_real;
  reg        [17:0]   img_reg_array_16_0_imag;
  reg        [17:0]   img_reg_array_16_1_real;
  reg        [17:0]   img_reg_array_16_1_imag;
  reg        [17:0]   img_reg_array_16_2_real;
  reg        [17:0]   img_reg_array_16_2_imag;
  reg        [17:0]   img_reg_array_16_3_real;
  reg        [17:0]   img_reg_array_16_3_imag;
  reg        [17:0]   img_reg_array_16_4_real;
  reg        [17:0]   img_reg_array_16_4_imag;
  reg        [17:0]   img_reg_array_16_5_real;
  reg        [17:0]   img_reg_array_16_5_imag;
  reg        [17:0]   img_reg_array_16_6_real;
  reg        [17:0]   img_reg_array_16_6_imag;
  reg        [17:0]   img_reg_array_16_7_real;
  reg        [17:0]   img_reg_array_16_7_imag;
  reg        [17:0]   img_reg_array_16_8_real;
  reg        [17:0]   img_reg_array_16_8_imag;
  reg        [17:0]   img_reg_array_16_9_real;
  reg        [17:0]   img_reg_array_16_9_imag;
  reg        [17:0]   img_reg_array_16_10_real;
  reg        [17:0]   img_reg_array_16_10_imag;
  reg        [17:0]   img_reg_array_16_11_real;
  reg        [17:0]   img_reg_array_16_11_imag;
  reg        [17:0]   img_reg_array_16_12_real;
  reg        [17:0]   img_reg_array_16_12_imag;
  reg        [17:0]   img_reg_array_16_13_real;
  reg        [17:0]   img_reg_array_16_13_imag;
  reg        [17:0]   img_reg_array_16_14_real;
  reg        [17:0]   img_reg_array_16_14_imag;
  reg        [17:0]   img_reg_array_16_15_real;
  reg        [17:0]   img_reg_array_16_15_imag;
  reg        [17:0]   img_reg_array_16_16_real;
  reg        [17:0]   img_reg_array_16_16_imag;
  reg        [17:0]   img_reg_array_16_17_real;
  reg        [17:0]   img_reg_array_16_17_imag;
  reg        [17:0]   img_reg_array_16_18_real;
  reg        [17:0]   img_reg_array_16_18_imag;
  reg        [17:0]   img_reg_array_16_19_real;
  reg        [17:0]   img_reg_array_16_19_imag;
  reg        [17:0]   img_reg_array_16_20_real;
  reg        [17:0]   img_reg_array_16_20_imag;
  reg        [17:0]   img_reg_array_16_21_real;
  reg        [17:0]   img_reg_array_16_21_imag;
  reg        [17:0]   img_reg_array_16_22_real;
  reg        [17:0]   img_reg_array_16_22_imag;
  reg        [17:0]   img_reg_array_16_23_real;
  reg        [17:0]   img_reg_array_16_23_imag;
  reg        [17:0]   img_reg_array_16_24_real;
  reg        [17:0]   img_reg_array_16_24_imag;
  reg        [17:0]   img_reg_array_16_25_real;
  reg        [17:0]   img_reg_array_16_25_imag;
  reg        [17:0]   img_reg_array_16_26_real;
  reg        [17:0]   img_reg_array_16_26_imag;
  reg        [17:0]   img_reg_array_16_27_real;
  reg        [17:0]   img_reg_array_16_27_imag;
  reg        [17:0]   img_reg_array_16_28_real;
  reg        [17:0]   img_reg_array_16_28_imag;
  reg        [17:0]   img_reg_array_16_29_real;
  reg        [17:0]   img_reg_array_16_29_imag;
  reg        [17:0]   img_reg_array_16_30_real;
  reg        [17:0]   img_reg_array_16_30_imag;
  reg        [17:0]   img_reg_array_16_31_real;
  reg        [17:0]   img_reg_array_16_31_imag;
  reg        [17:0]   img_reg_array_16_32_real;
  reg        [17:0]   img_reg_array_16_32_imag;
  reg        [17:0]   img_reg_array_16_33_real;
  reg        [17:0]   img_reg_array_16_33_imag;
  reg        [17:0]   img_reg_array_16_34_real;
  reg        [17:0]   img_reg_array_16_34_imag;
  reg        [17:0]   img_reg_array_16_35_real;
  reg        [17:0]   img_reg_array_16_35_imag;
  reg        [17:0]   img_reg_array_16_36_real;
  reg        [17:0]   img_reg_array_16_36_imag;
  reg        [17:0]   img_reg_array_16_37_real;
  reg        [17:0]   img_reg_array_16_37_imag;
  reg        [17:0]   img_reg_array_16_38_real;
  reg        [17:0]   img_reg_array_16_38_imag;
  reg        [17:0]   img_reg_array_16_39_real;
  reg        [17:0]   img_reg_array_16_39_imag;
  reg        [17:0]   img_reg_array_16_40_real;
  reg        [17:0]   img_reg_array_16_40_imag;
  reg        [17:0]   img_reg_array_16_41_real;
  reg        [17:0]   img_reg_array_16_41_imag;
  reg        [17:0]   img_reg_array_16_42_real;
  reg        [17:0]   img_reg_array_16_42_imag;
  reg        [17:0]   img_reg_array_16_43_real;
  reg        [17:0]   img_reg_array_16_43_imag;
  reg        [17:0]   img_reg_array_16_44_real;
  reg        [17:0]   img_reg_array_16_44_imag;
  reg        [17:0]   img_reg_array_16_45_real;
  reg        [17:0]   img_reg_array_16_45_imag;
  reg        [17:0]   img_reg_array_16_46_real;
  reg        [17:0]   img_reg_array_16_46_imag;
  reg        [17:0]   img_reg_array_16_47_real;
  reg        [17:0]   img_reg_array_16_47_imag;
  reg        [17:0]   img_reg_array_16_48_real;
  reg        [17:0]   img_reg_array_16_48_imag;
  reg        [17:0]   img_reg_array_16_49_real;
  reg        [17:0]   img_reg_array_16_49_imag;
  reg        [17:0]   img_reg_array_16_50_real;
  reg        [17:0]   img_reg_array_16_50_imag;
  reg        [17:0]   img_reg_array_16_51_real;
  reg        [17:0]   img_reg_array_16_51_imag;
  reg        [17:0]   img_reg_array_16_52_real;
  reg        [17:0]   img_reg_array_16_52_imag;
  reg        [17:0]   img_reg_array_16_53_real;
  reg        [17:0]   img_reg_array_16_53_imag;
  reg        [17:0]   img_reg_array_16_54_real;
  reg        [17:0]   img_reg_array_16_54_imag;
  reg        [17:0]   img_reg_array_16_55_real;
  reg        [17:0]   img_reg_array_16_55_imag;
  reg        [17:0]   img_reg_array_16_56_real;
  reg        [17:0]   img_reg_array_16_56_imag;
  reg        [17:0]   img_reg_array_16_57_real;
  reg        [17:0]   img_reg_array_16_57_imag;
  reg        [17:0]   img_reg_array_16_58_real;
  reg        [17:0]   img_reg_array_16_58_imag;
  reg        [17:0]   img_reg_array_16_59_real;
  reg        [17:0]   img_reg_array_16_59_imag;
  reg        [17:0]   img_reg_array_16_60_real;
  reg        [17:0]   img_reg_array_16_60_imag;
  reg        [17:0]   img_reg_array_16_61_real;
  reg        [17:0]   img_reg_array_16_61_imag;
  reg        [17:0]   img_reg_array_16_62_real;
  reg        [17:0]   img_reg_array_16_62_imag;
  reg        [17:0]   img_reg_array_16_63_real;
  reg        [17:0]   img_reg_array_16_63_imag;
  reg        [17:0]   img_reg_array_17_0_real;
  reg        [17:0]   img_reg_array_17_0_imag;
  reg        [17:0]   img_reg_array_17_1_real;
  reg        [17:0]   img_reg_array_17_1_imag;
  reg        [17:0]   img_reg_array_17_2_real;
  reg        [17:0]   img_reg_array_17_2_imag;
  reg        [17:0]   img_reg_array_17_3_real;
  reg        [17:0]   img_reg_array_17_3_imag;
  reg        [17:0]   img_reg_array_17_4_real;
  reg        [17:0]   img_reg_array_17_4_imag;
  reg        [17:0]   img_reg_array_17_5_real;
  reg        [17:0]   img_reg_array_17_5_imag;
  reg        [17:0]   img_reg_array_17_6_real;
  reg        [17:0]   img_reg_array_17_6_imag;
  reg        [17:0]   img_reg_array_17_7_real;
  reg        [17:0]   img_reg_array_17_7_imag;
  reg        [17:0]   img_reg_array_17_8_real;
  reg        [17:0]   img_reg_array_17_8_imag;
  reg        [17:0]   img_reg_array_17_9_real;
  reg        [17:0]   img_reg_array_17_9_imag;
  reg        [17:0]   img_reg_array_17_10_real;
  reg        [17:0]   img_reg_array_17_10_imag;
  reg        [17:0]   img_reg_array_17_11_real;
  reg        [17:0]   img_reg_array_17_11_imag;
  reg        [17:0]   img_reg_array_17_12_real;
  reg        [17:0]   img_reg_array_17_12_imag;
  reg        [17:0]   img_reg_array_17_13_real;
  reg        [17:0]   img_reg_array_17_13_imag;
  reg        [17:0]   img_reg_array_17_14_real;
  reg        [17:0]   img_reg_array_17_14_imag;
  reg        [17:0]   img_reg_array_17_15_real;
  reg        [17:0]   img_reg_array_17_15_imag;
  reg        [17:0]   img_reg_array_17_16_real;
  reg        [17:0]   img_reg_array_17_16_imag;
  reg        [17:0]   img_reg_array_17_17_real;
  reg        [17:0]   img_reg_array_17_17_imag;
  reg        [17:0]   img_reg_array_17_18_real;
  reg        [17:0]   img_reg_array_17_18_imag;
  reg        [17:0]   img_reg_array_17_19_real;
  reg        [17:0]   img_reg_array_17_19_imag;
  reg        [17:0]   img_reg_array_17_20_real;
  reg        [17:0]   img_reg_array_17_20_imag;
  reg        [17:0]   img_reg_array_17_21_real;
  reg        [17:0]   img_reg_array_17_21_imag;
  reg        [17:0]   img_reg_array_17_22_real;
  reg        [17:0]   img_reg_array_17_22_imag;
  reg        [17:0]   img_reg_array_17_23_real;
  reg        [17:0]   img_reg_array_17_23_imag;
  reg        [17:0]   img_reg_array_17_24_real;
  reg        [17:0]   img_reg_array_17_24_imag;
  reg        [17:0]   img_reg_array_17_25_real;
  reg        [17:0]   img_reg_array_17_25_imag;
  reg        [17:0]   img_reg_array_17_26_real;
  reg        [17:0]   img_reg_array_17_26_imag;
  reg        [17:0]   img_reg_array_17_27_real;
  reg        [17:0]   img_reg_array_17_27_imag;
  reg        [17:0]   img_reg_array_17_28_real;
  reg        [17:0]   img_reg_array_17_28_imag;
  reg        [17:0]   img_reg_array_17_29_real;
  reg        [17:0]   img_reg_array_17_29_imag;
  reg        [17:0]   img_reg_array_17_30_real;
  reg        [17:0]   img_reg_array_17_30_imag;
  reg        [17:0]   img_reg_array_17_31_real;
  reg        [17:0]   img_reg_array_17_31_imag;
  reg        [17:0]   img_reg_array_17_32_real;
  reg        [17:0]   img_reg_array_17_32_imag;
  reg        [17:0]   img_reg_array_17_33_real;
  reg        [17:0]   img_reg_array_17_33_imag;
  reg        [17:0]   img_reg_array_17_34_real;
  reg        [17:0]   img_reg_array_17_34_imag;
  reg        [17:0]   img_reg_array_17_35_real;
  reg        [17:0]   img_reg_array_17_35_imag;
  reg        [17:0]   img_reg_array_17_36_real;
  reg        [17:0]   img_reg_array_17_36_imag;
  reg        [17:0]   img_reg_array_17_37_real;
  reg        [17:0]   img_reg_array_17_37_imag;
  reg        [17:0]   img_reg_array_17_38_real;
  reg        [17:0]   img_reg_array_17_38_imag;
  reg        [17:0]   img_reg_array_17_39_real;
  reg        [17:0]   img_reg_array_17_39_imag;
  reg        [17:0]   img_reg_array_17_40_real;
  reg        [17:0]   img_reg_array_17_40_imag;
  reg        [17:0]   img_reg_array_17_41_real;
  reg        [17:0]   img_reg_array_17_41_imag;
  reg        [17:0]   img_reg_array_17_42_real;
  reg        [17:0]   img_reg_array_17_42_imag;
  reg        [17:0]   img_reg_array_17_43_real;
  reg        [17:0]   img_reg_array_17_43_imag;
  reg        [17:0]   img_reg_array_17_44_real;
  reg        [17:0]   img_reg_array_17_44_imag;
  reg        [17:0]   img_reg_array_17_45_real;
  reg        [17:0]   img_reg_array_17_45_imag;
  reg        [17:0]   img_reg_array_17_46_real;
  reg        [17:0]   img_reg_array_17_46_imag;
  reg        [17:0]   img_reg_array_17_47_real;
  reg        [17:0]   img_reg_array_17_47_imag;
  reg        [17:0]   img_reg_array_17_48_real;
  reg        [17:0]   img_reg_array_17_48_imag;
  reg        [17:0]   img_reg_array_17_49_real;
  reg        [17:0]   img_reg_array_17_49_imag;
  reg        [17:0]   img_reg_array_17_50_real;
  reg        [17:0]   img_reg_array_17_50_imag;
  reg        [17:0]   img_reg_array_17_51_real;
  reg        [17:0]   img_reg_array_17_51_imag;
  reg        [17:0]   img_reg_array_17_52_real;
  reg        [17:0]   img_reg_array_17_52_imag;
  reg        [17:0]   img_reg_array_17_53_real;
  reg        [17:0]   img_reg_array_17_53_imag;
  reg        [17:0]   img_reg_array_17_54_real;
  reg        [17:0]   img_reg_array_17_54_imag;
  reg        [17:0]   img_reg_array_17_55_real;
  reg        [17:0]   img_reg_array_17_55_imag;
  reg        [17:0]   img_reg_array_17_56_real;
  reg        [17:0]   img_reg_array_17_56_imag;
  reg        [17:0]   img_reg_array_17_57_real;
  reg        [17:0]   img_reg_array_17_57_imag;
  reg        [17:0]   img_reg_array_17_58_real;
  reg        [17:0]   img_reg_array_17_58_imag;
  reg        [17:0]   img_reg_array_17_59_real;
  reg        [17:0]   img_reg_array_17_59_imag;
  reg        [17:0]   img_reg_array_17_60_real;
  reg        [17:0]   img_reg_array_17_60_imag;
  reg        [17:0]   img_reg_array_17_61_real;
  reg        [17:0]   img_reg_array_17_61_imag;
  reg        [17:0]   img_reg_array_17_62_real;
  reg        [17:0]   img_reg_array_17_62_imag;
  reg        [17:0]   img_reg_array_17_63_real;
  reg        [17:0]   img_reg_array_17_63_imag;
  reg        [17:0]   img_reg_array_18_0_real;
  reg        [17:0]   img_reg_array_18_0_imag;
  reg        [17:0]   img_reg_array_18_1_real;
  reg        [17:0]   img_reg_array_18_1_imag;
  reg        [17:0]   img_reg_array_18_2_real;
  reg        [17:0]   img_reg_array_18_2_imag;
  reg        [17:0]   img_reg_array_18_3_real;
  reg        [17:0]   img_reg_array_18_3_imag;
  reg        [17:0]   img_reg_array_18_4_real;
  reg        [17:0]   img_reg_array_18_4_imag;
  reg        [17:0]   img_reg_array_18_5_real;
  reg        [17:0]   img_reg_array_18_5_imag;
  reg        [17:0]   img_reg_array_18_6_real;
  reg        [17:0]   img_reg_array_18_6_imag;
  reg        [17:0]   img_reg_array_18_7_real;
  reg        [17:0]   img_reg_array_18_7_imag;
  reg        [17:0]   img_reg_array_18_8_real;
  reg        [17:0]   img_reg_array_18_8_imag;
  reg        [17:0]   img_reg_array_18_9_real;
  reg        [17:0]   img_reg_array_18_9_imag;
  reg        [17:0]   img_reg_array_18_10_real;
  reg        [17:0]   img_reg_array_18_10_imag;
  reg        [17:0]   img_reg_array_18_11_real;
  reg        [17:0]   img_reg_array_18_11_imag;
  reg        [17:0]   img_reg_array_18_12_real;
  reg        [17:0]   img_reg_array_18_12_imag;
  reg        [17:0]   img_reg_array_18_13_real;
  reg        [17:0]   img_reg_array_18_13_imag;
  reg        [17:0]   img_reg_array_18_14_real;
  reg        [17:0]   img_reg_array_18_14_imag;
  reg        [17:0]   img_reg_array_18_15_real;
  reg        [17:0]   img_reg_array_18_15_imag;
  reg        [17:0]   img_reg_array_18_16_real;
  reg        [17:0]   img_reg_array_18_16_imag;
  reg        [17:0]   img_reg_array_18_17_real;
  reg        [17:0]   img_reg_array_18_17_imag;
  reg        [17:0]   img_reg_array_18_18_real;
  reg        [17:0]   img_reg_array_18_18_imag;
  reg        [17:0]   img_reg_array_18_19_real;
  reg        [17:0]   img_reg_array_18_19_imag;
  reg        [17:0]   img_reg_array_18_20_real;
  reg        [17:0]   img_reg_array_18_20_imag;
  reg        [17:0]   img_reg_array_18_21_real;
  reg        [17:0]   img_reg_array_18_21_imag;
  reg        [17:0]   img_reg_array_18_22_real;
  reg        [17:0]   img_reg_array_18_22_imag;
  reg        [17:0]   img_reg_array_18_23_real;
  reg        [17:0]   img_reg_array_18_23_imag;
  reg        [17:0]   img_reg_array_18_24_real;
  reg        [17:0]   img_reg_array_18_24_imag;
  reg        [17:0]   img_reg_array_18_25_real;
  reg        [17:0]   img_reg_array_18_25_imag;
  reg        [17:0]   img_reg_array_18_26_real;
  reg        [17:0]   img_reg_array_18_26_imag;
  reg        [17:0]   img_reg_array_18_27_real;
  reg        [17:0]   img_reg_array_18_27_imag;
  reg        [17:0]   img_reg_array_18_28_real;
  reg        [17:0]   img_reg_array_18_28_imag;
  reg        [17:0]   img_reg_array_18_29_real;
  reg        [17:0]   img_reg_array_18_29_imag;
  reg        [17:0]   img_reg_array_18_30_real;
  reg        [17:0]   img_reg_array_18_30_imag;
  reg        [17:0]   img_reg_array_18_31_real;
  reg        [17:0]   img_reg_array_18_31_imag;
  reg        [17:0]   img_reg_array_18_32_real;
  reg        [17:0]   img_reg_array_18_32_imag;
  reg        [17:0]   img_reg_array_18_33_real;
  reg        [17:0]   img_reg_array_18_33_imag;
  reg        [17:0]   img_reg_array_18_34_real;
  reg        [17:0]   img_reg_array_18_34_imag;
  reg        [17:0]   img_reg_array_18_35_real;
  reg        [17:0]   img_reg_array_18_35_imag;
  reg        [17:0]   img_reg_array_18_36_real;
  reg        [17:0]   img_reg_array_18_36_imag;
  reg        [17:0]   img_reg_array_18_37_real;
  reg        [17:0]   img_reg_array_18_37_imag;
  reg        [17:0]   img_reg_array_18_38_real;
  reg        [17:0]   img_reg_array_18_38_imag;
  reg        [17:0]   img_reg_array_18_39_real;
  reg        [17:0]   img_reg_array_18_39_imag;
  reg        [17:0]   img_reg_array_18_40_real;
  reg        [17:0]   img_reg_array_18_40_imag;
  reg        [17:0]   img_reg_array_18_41_real;
  reg        [17:0]   img_reg_array_18_41_imag;
  reg        [17:0]   img_reg_array_18_42_real;
  reg        [17:0]   img_reg_array_18_42_imag;
  reg        [17:0]   img_reg_array_18_43_real;
  reg        [17:0]   img_reg_array_18_43_imag;
  reg        [17:0]   img_reg_array_18_44_real;
  reg        [17:0]   img_reg_array_18_44_imag;
  reg        [17:0]   img_reg_array_18_45_real;
  reg        [17:0]   img_reg_array_18_45_imag;
  reg        [17:0]   img_reg_array_18_46_real;
  reg        [17:0]   img_reg_array_18_46_imag;
  reg        [17:0]   img_reg_array_18_47_real;
  reg        [17:0]   img_reg_array_18_47_imag;
  reg        [17:0]   img_reg_array_18_48_real;
  reg        [17:0]   img_reg_array_18_48_imag;
  reg        [17:0]   img_reg_array_18_49_real;
  reg        [17:0]   img_reg_array_18_49_imag;
  reg        [17:0]   img_reg_array_18_50_real;
  reg        [17:0]   img_reg_array_18_50_imag;
  reg        [17:0]   img_reg_array_18_51_real;
  reg        [17:0]   img_reg_array_18_51_imag;
  reg        [17:0]   img_reg_array_18_52_real;
  reg        [17:0]   img_reg_array_18_52_imag;
  reg        [17:0]   img_reg_array_18_53_real;
  reg        [17:0]   img_reg_array_18_53_imag;
  reg        [17:0]   img_reg_array_18_54_real;
  reg        [17:0]   img_reg_array_18_54_imag;
  reg        [17:0]   img_reg_array_18_55_real;
  reg        [17:0]   img_reg_array_18_55_imag;
  reg        [17:0]   img_reg_array_18_56_real;
  reg        [17:0]   img_reg_array_18_56_imag;
  reg        [17:0]   img_reg_array_18_57_real;
  reg        [17:0]   img_reg_array_18_57_imag;
  reg        [17:0]   img_reg_array_18_58_real;
  reg        [17:0]   img_reg_array_18_58_imag;
  reg        [17:0]   img_reg_array_18_59_real;
  reg        [17:0]   img_reg_array_18_59_imag;
  reg        [17:0]   img_reg_array_18_60_real;
  reg        [17:0]   img_reg_array_18_60_imag;
  reg        [17:0]   img_reg_array_18_61_real;
  reg        [17:0]   img_reg_array_18_61_imag;
  reg        [17:0]   img_reg_array_18_62_real;
  reg        [17:0]   img_reg_array_18_62_imag;
  reg        [17:0]   img_reg_array_18_63_real;
  reg        [17:0]   img_reg_array_18_63_imag;
  reg        [17:0]   img_reg_array_19_0_real;
  reg        [17:0]   img_reg_array_19_0_imag;
  reg        [17:0]   img_reg_array_19_1_real;
  reg        [17:0]   img_reg_array_19_1_imag;
  reg        [17:0]   img_reg_array_19_2_real;
  reg        [17:0]   img_reg_array_19_2_imag;
  reg        [17:0]   img_reg_array_19_3_real;
  reg        [17:0]   img_reg_array_19_3_imag;
  reg        [17:0]   img_reg_array_19_4_real;
  reg        [17:0]   img_reg_array_19_4_imag;
  reg        [17:0]   img_reg_array_19_5_real;
  reg        [17:0]   img_reg_array_19_5_imag;
  reg        [17:0]   img_reg_array_19_6_real;
  reg        [17:0]   img_reg_array_19_6_imag;
  reg        [17:0]   img_reg_array_19_7_real;
  reg        [17:0]   img_reg_array_19_7_imag;
  reg        [17:0]   img_reg_array_19_8_real;
  reg        [17:0]   img_reg_array_19_8_imag;
  reg        [17:0]   img_reg_array_19_9_real;
  reg        [17:0]   img_reg_array_19_9_imag;
  reg        [17:0]   img_reg_array_19_10_real;
  reg        [17:0]   img_reg_array_19_10_imag;
  reg        [17:0]   img_reg_array_19_11_real;
  reg        [17:0]   img_reg_array_19_11_imag;
  reg        [17:0]   img_reg_array_19_12_real;
  reg        [17:0]   img_reg_array_19_12_imag;
  reg        [17:0]   img_reg_array_19_13_real;
  reg        [17:0]   img_reg_array_19_13_imag;
  reg        [17:0]   img_reg_array_19_14_real;
  reg        [17:0]   img_reg_array_19_14_imag;
  reg        [17:0]   img_reg_array_19_15_real;
  reg        [17:0]   img_reg_array_19_15_imag;
  reg        [17:0]   img_reg_array_19_16_real;
  reg        [17:0]   img_reg_array_19_16_imag;
  reg        [17:0]   img_reg_array_19_17_real;
  reg        [17:0]   img_reg_array_19_17_imag;
  reg        [17:0]   img_reg_array_19_18_real;
  reg        [17:0]   img_reg_array_19_18_imag;
  reg        [17:0]   img_reg_array_19_19_real;
  reg        [17:0]   img_reg_array_19_19_imag;
  reg        [17:0]   img_reg_array_19_20_real;
  reg        [17:0]   img_reg_array_19_20_imag;
  reg        [17:0]   img_reg_array_19_21_real;
  reg        [17:0]   img_reg_array_19_21_imag;
  reg        [17:0]   img_reg_array_19_22_real;
  reg        [17:0]   img_reg_array_19_22_imag;
  reg        [17:0]   img_reg_array_19_23_real;
  reg        [17:0]   img_reg_array_19_23_imag;
  reg        [17:0]   img_reg_array_19_24_real;
  reg        [17:0]   img_reg_array_19_24_imag;
  reg        [17:0]   img_reg_array_19_25_real;
  reg        [17:0]   img_reg_array_19_25_imag;
  reg        [17:0]   img_reg_array_19_26_real;
  reg        [17:0]   img_reg_array_19_26_imag;
  reg        [17:0]   img_reg_array_19_27_real;
  reg        [17:0]   img_reg_array_19_27_imag;
  reg        [17:0]   img_reg_array_19_28_real;
  reg        [17:0]   img_reg_array_19_28_imag;
  reg        [17:0]   img_reg_array_19_29_real;
  reg        [17:0]   img_reg_array_19_29_imag;
  reg        [17:0]   img_reg_array_19_30_real;
  reg        [17:0]   img_reg_array_19_30_imag;
  reg        [17:0]   img_reg_array_19_31_real;
  reg        [17:0]   img_reg_array_19_31_imag;
  reg        [17:0]   img_reg_array_19_32_real;
  reg        [17:0]   img_reg_array_19_32_imag;
  reg        [17:0]   img_reg_array_19_33_real;
  reg        [17:0]   img_reg_array_19_33_imag;
  reg        [17:0]   img_reg_array_19_34_real;
  reg        [17:0]   img_reg_array_19_34_imag;
  reg        [17:0]   img_reg_array_19_35_real;
  reg        [17:0]   img_reg_array_19_35_imag;
  reg        [17:0]   img_reg_array_19_36_real;
  reg        [17:0]   img_reg_array_19_36_imag;
  reg        [17:0]   img_reg_array_19_37_real;
  reg        [17:0]   img_reg_array_19_37_imag;
  reg        [17:0]   img_reg_array_19_38_real;
  reg        [17:0]   img_reg_array_19_38_imag;
  reg        [17:0]   img_reg_array_19_39_real;
  reg        [17:0]   img_reg_array_19_39_imag;
  reg        [17:0]   img_reg_array_19_40_real;
  reg        [17:0]   img_reg_array_19_40_imag;
  reg        [17:0]   img_reg_array_19_41_real;
  reg        [17:0]   img_reg_array_19_41_imag;
  reg        [17:0]   img_reg_array_19_42_real;
  reg        [17:0]   img_reg_array_19_42_imag;
  reg        [17:0]   img_reg_array_19_43_real;
  reg        [17:0]   img_reg_array_19_43_imag;
  reg        [17:0]   img_reg_array_19_44_real;
  reg        [17:0]   img_reg_array_19_44_imag;
  reg        [17:0]   img_reg_array_19_45_real;
  reg        [17:0]   img_reg_array_19_45_imag;
  reg        [17:0]   img_reg_array_19_46_real;
  reg        [17:0]   img_reg_array_19_46_imag;
  reg        [17:0]   img_reg_array_19_47_real;
  reg        [17:0]   img_reg_array_19_47_imag;
  reg        [17:0]   img_reg_array_19_48_real;
  reg        [17:0]   img_reg_array_19_48_imag;
  reg        [17:0]   img_reg_array_19_49_real;
  reg        [17:0]   img_reg_array_19_49_imag;
  reg        [17:0]   img_reg_array_19_50_real;
  reg        [17:0]   img_reg_array_19_50_imag;
  reg        [17:0]   img_reg_array_19_51_real;
  reg        [17:0]   img_reg_array_19_51_imag;
  reg        [17:0]   img_reg_array_19_52_real;
  reg        [17:0]   img_reg_array_19_52_imag;
  reg        [17:0]   img_reg_array_19_53_real;
  reg        [17:0]   img_reg_array_19_53_imag;
  reg        [17:0]   img_reg_array_19_54_real;
  reg        [17:0]   img_reg_array_19_54_imag;
  reg        [17:0]   img_reg_array_19_55_real;
  reg        [17:0]   img_reg_array_19_55_imag;
  reg        [17:0]   img_reg_array_19_56_real;
  reg        [17:0]   img_reg_array_19_56_imag;
  reg        [17:0]   img_reg_array_19_57_real;
  reg        [17:0]   img_reg_array_19_57_imag;
  reg        [17:0]   img_reg_array_19_58_real;
  reg        [17:0]   img_reg_array_19_58_imag;
  reg        [17:0]   img_reg_array_19_59_real;
  reg        [17:0]   img_reg_array_19_59_imag;
  reg        [17:0]   img_reg_array_19_60_real;
  reg        [17:0]   img_reg_array_19_60_imag;
  reg        [17:0]   img_reg_array_19_61_real;
  reg        [17:0]   img_reg_array_19_61_imag;
  reg        [17:0]   img_reg_array_19_62_real;
  reg        [17:0]   img_reg_array_19_62_imag;
  reg        [17:0]   img_reg_array_19_63_real;
  reg        [17:0]   img_reg_array_19_63_imag;
  reg        [17:0]   img_reg_array_20_0_real;
  reg        [17:0]   img_reg_array_20_0_imag;
  reg        [17:0]   img_reg_array_20_1_real;
  reg        [17:0]   img_reg_array_20_1_imag;
  reg        [17:0]   img_reg_array_20_2_real;
  reg        [17:0]   img_reg_array_20_2_imag;
  reg        [17:0]   img_reg_array_20_3_real;
  reg        [17:0]   img_reg_array_20_3_imag;
  reg        [17:0]   img_reg_array_20_4_real;
  reg        [17:0]   img_reg_array_20_4_imag;
  reg        [17:0]   img_reg_array_20_5_real;
  reg        [17:0]   img_reg_array_20_5_imag;
  reg        [17:0]   img_reg_array_20_6_real;
  reg        [17:0]   img_reg_array_20_6_imag;
  reg        [17:0]   img_reg_array_20_7_real;
  reg        [17:0]   img_reg_array_20_7_imag;
  reg        [17:0]   img_reg_array_20_8_real;
  reg        [17:0]   img_reg_array_20_8_imag;
  reg        [17:0]   img_reg_array_20_9_real;
  reg        [17:0]   img_reg_array_20_9_imag;
  reg        [17:0]   img_reg_array_20_10_real;
  reg        [17:0]   img_reg_array_20_10_imag;
  reg        [17:0]   img_reg_array_20_11_real;
  reg        [17:0]   img_reg_array_20_11_imag;
  reg        [17:0]   img_reg_array_20_12_real;
  reg        [17:0]   img_reg_array_20_12_imag;
  reg        [17:0]   img_reg_array_20_13_real;
  reg        [17:0]   img_reg_array_20_13_imag;
  reg        [17:0]   img_reg_array_20_14_real;
  reg        [17:0]   img_reg_array_20_14_imag;
  reg        [17:0]   img_reg_array_20_15_real;
  reg        [17:0]   img_reg_array_20_15_imag;
  reg        [17:0]   img_reg_array_20_16_real;
  reg        [17:0]   img_reg_array_20_16_imag;
  reg        [17:0]   img_reg_array_20_17_real;
  reg        [17:0]   img_reg_array_20_17_imag;
  reg        [17:0]   img_reg_array_20_18_real;
  reg        [17:0]   img_reg_array_20_18_imag;
  reg        [17:0]   img_reg_array_20_19_real;
  reg        [17:0]   img_reg_array_20_19_imag;
  reg        [17:0]   img_reg_array_20_20_real;
  reg        [17:0]   img_reg_array_20_20_imag;
  reg        [17:0]   img_reg_array_20_21_real;
  reg        [17:0]   img_reg_array_20_21_imag;
  reg        [17:0]   img_reg_array_20_22_real;
  reg        [17:0]   img_reg_array_20_22_imag;
  reg        [17:0]   img_reg_array_20_23_real;
  reg        [17:0]   img_reg_array_20_23_imag;
  reg        [17:0]   img_reg_array_20_24_real;
  reg        [17:0]   img_reg_array_20_24_imag;
  reg        [17:0]   img_reg_array_20_25_real;
  reg        [17:0]   img_reg_array_20_25_imag;
  reg        [17:0]   img_reg_array_20_26_real;
  reg        [17:0]   img_reg_array_20_26_imag;
  reg        [17:0]   img_reg_array_20_27_real;
  reg        [17:0]   img_reg_array_20_27_imag;
  reg        [17:0]   img_reg_array_20_28_real;
  reg        [17:0]   img_reg_array_20_28_imag;
  reg        [17:0]   img_reg_array_20_29_real;
  reg        [17:0]   img_reg_array_20_29_imag;
  reg        [17:0]   img_reg_array_20_30_real;
  reg        [17:0]   img_reg_array_20_30_imag;
  reg        [17:0]   img_reg_array_20_31_real;
  reg        [17:0]   img_reg_array_20_31_imag;
  reg        [17:0]   img_reg_array_20_32_real;
  reg        [17:0]   img_reg_array_20_32_imag;
  reg        [17:0]   img_reg_array_20_33_real;
  reg        [17:0]   img_reg_array_20_33_imag;
  reg        [17:0]   img_reg_array_20_34_real;
  reg        [17:0]   img_reg_array_20_34_imag;
  reg        [17:0]   img_reg_array_20_35_real;
  reg        [17:0]   img_reg_array_20_35_imag;
  reg        [17:0]   img_reg_array_20_36_real;
  reg        [17:0]   img_reg_array_20_36_imag;
  reg        [17:0]   img_reg_array_20_37_real;
  reg        [17:0]   img_reg_array_20_37_imag;
  reg        [17:0]   img_reg_array_20_38_real;
  reg        [17:0]   img_reg_array_20_38_imag;
  reg        [17:0]   img_reg_array_20_39_real;
  reg        [17:0]   img_reg_array_20_39_imag;
  reg        [17:0]   img_reg_array_20_40_real;
  reg        [17:0]   img_reg_array_20_40_imag;
  reg        [17:0]   img_reg_array_20_41_real;
  reg        [17:0]   img_reg_array_20_41_imag;
  reg        [17:0]   img_reg_array_20_42_real;
  reg        [17:0]   img_reg_array_20_42_imag;
  reg        [17:0]   img_reg_array_20_43_real;
  reg        [17:0]   img_reg_array_20_43_imag;
  reg        [17:0]   img_reg_array_20_44_real;
  reg        [17:0]   img_reg_array_20_44_imag;
  reg        [17:0]   img_reg_array_20_45_real;
  reg        [17:0]   img_reg_array_20_45_imag;
  reg        [17:0]   img_reg_array_20_46_real;
  reg        [17:0]   img_reg_array_20_46_imag;
  reg        [17:0]   img_reg_array_20_47_real;
  reg        [17:0]   img_reg_array_20_47_imag;
  reg        [17:0]   img_reg_array_20_48_real;
  reg        [17:0]   img_reg_array_20_48_imag;
  reg        [17:0]   img_reg_array_20_49_real;
  reg        [17:0]   img_reg_array_20_49_imag;
  reg        [17:0]   img_reg_array_20_50_real;
  reg        [17:0]   img_reg_array_20_50_imag;
  reg        [17:0]   img_reg_array_20_51_real;
  reg        [17:0]   img_reg_array_20_51_imag;
  reg        [17:0]   img_reg_array_20_52_real;
  reg        [17:0]   img_reg_array_20_52_imag;
  reg        [17:0]   img_reg_array_20_53_real;
  reg        [17:0]   img_reg_array_20_53_imag;
  reg        [17:0]   img_reg_array_20_54_real;
  reg        [17:0]   img_reg_array_20_54_imag;
  reg        [17:0]   img_reg_array_20_55_real;
  reg        [17:0]   img_reg_array_20_55_imag;
  reg        [17:0]   img_reg_array_20_56_real;
  reg        [17:0]   img_reg_array_20_56_imag;
  reg        [17:0]   img_reg_array_20_57_real;
  reg        [17:0]   img_reg_array_20_57_imag;
  reg        [17:0]   img_reg_array_20_58_real;
  reg        [17:0]   img_reg_array_20_58_imag;
  reg        [17:0]   img_reg_array_20_59_real;
  reg        [17:0]   img_reg_array_20_59_imag;
  reg        [17:0]   img_reg_array_20_60_real;
  reg        [17:0]   img_reg_array_20_60_imag;
  reg        [17:0]   img_reg_array_20_61_real;
  reg        [17:0]   img_reg_array_20_61_imag;
  reg        [17:0]   img_reg_array_20_62_real;
  reg        [17:0]   img_reg_array_20_62_imag;
  reg        [17:0]   img_reg_array_20_63_real;
  reg        [17:0]   img_reg_array_20_63_imag;
  reg        [17:0]   img_reg_array_21_0_real;
  reg        [17:0]   img_reg_array_21_0_imag;
  reg        [17:0]   img_reg_array_21_1_real;
  reg        [17:0]   img_reg_array_21_1_imag;
  reg        [17:0]   img_reg_array_21_2_real;
  reg        [17:0]   img_reg_array_21_2_imag;
  reg        [17:0]   img_reg_array_21_3_real;
  reg        [17:0]   img_reg_array_21_3_imag;
  reg        [17:0]   img_reg_array_21_4_real;
  reg        [17:0]   img_reg_array_21_4_imag;
  reg        [17:0]   img_reg_array_21_5_real;
  reg        [17:0]   img_reg_array_21_5_imag;
  reg        [17:0]   img_reg_array_21_6_real;
  reg        [17:0]   img_reg_array_21_6_imag;
  reg        [17:0]   img_reg_array_21_7_real;
  reg        [17:0]   img_reg_array_21_7_imag;
  reg        [17:0]   img_reg_array_21_8_real;
  reg        [17:0]   img_reg_array_21_8_imag;
  reg        [17:0]   img_reg_array_21_9_real;
  reg        [17:0]   img_reg_array_21_9_imag;
  reg        [17:0]   img_reg_array_21_10_real;
  reg        [17:0]   img_reg_array_21_10_imag;
  reg        [17:0]   img_reg_array_21_11_real;
  reg        [17:0]   img_reg_array_21_11_imag;
  reg        [17:0]   img_reg_array_21_12_real;
  reg        [17:0]   img_reg_array_21_12_imag;
  reg        [17:0]   img_reg_array_21_13_real;
  reg        [17:0]   img_reg_array_21_13_imag;
  reg        [17:0]   img_reg_array_21_14_real;
  reg        [17:0]   img_reg_array_21_14_imag;
  reg        [17:0]   img_reg_array_21_15_real;
  reg        [17:0]   img_reg_array_21_15_imag;
  reg        [17:0]   img_reg_array_21_16_real;
  reg        [17:0]   img_reg_array_21_16_imag;
  reg        [17:0]   img_reg_array_21_17_real;
  reg        [17:0]   img_reg_array_21_17_imag;
  reg        [17:0]   img_reg_array_21_18_real;
  reg        [17:0]   img_reg_array_21_18_imag;
  reg        [17:0]   img_reg_array_21_19_real;
  reg        [17:0]   img_reg_array_21_19_imag;
  reg        [17:0]   img_reg_array_21_20_real;
  reg        [17:0]   img_reg_array_21_20_imag;
  reg        [17:0]   img_reg_array_21_21_real;
  reg        [17:0]   img_reg_array_21_21_imag;
  reg        [17:0]   img_reg_array_21_22_real;
  reg        [17:0]   img_reg_array_21_22_imag;
  reg        [17:0]   img_reg_array_21_23_real;
  reg        [17:0]   img_reg_array_21_23_imag;
  reg        [17:0]   img_reg_array_21_24_real;
  reg        [17:0]   img_reg_array_21_24_imag;
  reg        [17:0]   img_reg_array_21_25_real;
  reg        [17:0]   img_reg_array_21_25_imag;
  reg        [17:0]   img_reg_array_21_26_real;
  reg        [17:0]   img_reg_array_21_26_imag;
  reg        [17:0]   img_reg_array_21_27_real;
  reg        [17:0]   img_reg_array_21_27_imag;
  reg        [17:0]   img_reg_array_21_28_real;
  reg        [17:0]   img_reg_array_21_28_imag;
  reg        [17:0]   img_reg_array_21_29_real;
  reg        [17:0]   img_reg_array_21_29_imag;
  reg        [17:0]   img_reg_array_21_30_real;
  reg        [17:0]   img_reg_array_21_30_imag;
  reg        [17:0]   img_reg_array_21_31_real;
  reg        [17:0]   img_reg_array_21_31_imag;
  reg        [17:0]   img_reg_array_21_32_real;
  reg        [17:0]   img_reg_array_21_32_imag;
  reg        [17:0]   img_reg_array_21_33_real;
  reg        [17:0]   img_reg_array_21_33_imag;
  reg        [17:0]   img_reg_array_21_34_real;
  reg        [17:0]   img_reg_array_21_34_imag;
  reg        [17:0]   img_reg_array_21_35_real;
  reg        [17:0]   img_reg_array_21_35_imag;
  reg        [17:0]   img_reg_array_21_36_real;
  reg        [17:0]   img_reg_array_21_36_imag;
  reg        [17:0]   img_reg_array_21_37_real;
  reg        [17:0]   img_reg_array_21_37_imag;
  reg        [17:0]   img_reg_array_21_38_real;
  reg        [17:0]   img_reg_array_21_38_imag;
  reg        [17:0]   img_reg_array_21_39_real;
  reg        [17:0]   img_reg_array_21_39_imag;
  reg        [17:0]   img_reg_array_21_40_real;
  reg        [17:0]   img_reg_array_21_40_imag;
  reg        [17:0]   img_reg_array_21_41_real;
  reg        [17:0]   img_reg_array_21_41_imag;
  reg        [17:0]   img_reg_array_21_42_real;
  reg        [17:0]   img_reg_array_21_42_imag;
  reg        [17:0]   img_reg_array_21_43_real;
  reg        [17:0]   img_reg_array_21_43_imag;
  reg        [17:0]   img_reg_array_21_44_real;
  reg        [17:0]   img_reg_array_21_44_imag;
  reg        [17:0]   img_reg_array_21_45_real;
  reg        [17:0]   img_reg_array_21_45_imag;
  reg        [17:0]   img_reg_array_21_46_real;
  reg        [17:0]   img_reg_array_21_46_imag;
  reg        [17:0]   img_reg_array_21_47_real;
  reg        [17:0]   img_reg_array_21_47_imag;
  reg        [17:0]   img_reg_array_21_48_real;
  reg        [17:0]   img_reg_array_21_48_imag;
  reg        [17:0]   img_reg_array_21_49_real;
  reg        [17:0]   img_reg_array_21_49_imag;
  reg        [17:0]   img_reg_array_21_50_real;
  reg        [17:0]   img_reg_array_21_50_imag;
  reg        [17:0]   img_reg_array_21_51_real;
  reg        [17:0]   img_reg_array_21_51_imag;
  reg        [17:0]   img_reg_array_21_52_real;
  reg        [17:0]   img_reg_array_21_52_imag;
  reg        [17:0]   img_reg_array_21_53_real;
  reg        [17:0]   img_reg_array_21_53_imag;
  reg        [17:0]   img_reg_array_21_54_real;
  reg        [17:0]   img_reg_array_21_54_imag;
  reg        [17:0]   img_reg_array_21_55_real;
  reg        [17:0]   img_reg_array_21_55_imag;
  reg        [17:0]   img_reg_array_21_56_real;
  reg        [17:0]   img_reg_array_21_56_imag;
  reg        [17:0]   img_reg_array_21_57_real;
  reg        [17:0]   img_reg_array_21_57_imag;
  reg        [17:0]   img_reg_array_21_58_real;
  reg        [17:0]   img_reg_array_21_58_imag;
  reg        [17:0]   img_reg_array_21_59_real;
  reg        [17:0]   img_reg_array_21_59_imag;
  reg        [17:0]   img_reg_array_21_60_real;
  reg        [17:0]   img_reg_array_21_60_imag;
  reg        [17:0]   img_reg_array_21_61_real;
  reg        [17:0]   img_reg_array_21_61_imag;
  reg        [17:0]   img_reg_array_21_62_real;
  reg        [17:0]   img_reg_array_21_62_imag;
  reg        [17:0]   img_reg_array_21_63_real;
  reg        [17:0]   img_reg_array_21_63_imag;
  reg        [17:0]   img_reg_array_22_0_real;
  reg        [17:0]   img_reg_array_22_0_imag;
  reg        [17:0]   img_reg_array_22_1_real;
  reg        [17:0]   img_reg_array_22_1_imag;
  reg        [17:0]   img_reg_array_22_2_real;
  reg        [17:0]   img_reg_array_22_2_imag;
  reg        [17:0]   img_reg_array_22_3_real;
  reg        [17:0]   img_reg_array_22_3_imag;
  reg        [17:0]   img_reg_array_22_4_real;
  reg        [17:0]   img_reg_array_22_4_imag;
  reg        [17:0]   img_reg_array_22_5_real;
  reg        [17:0]   img_reg_array_22_5_imag;
  reg        [17:0]   img_reg_array_22_6_real;
  reg        [17:0]   img_reg_array_22_6_imag;
  reg        [17:0]   img_reg_array_22_7_real;
  reg        [17:0]   img_reg_array_22_7_imag;
  reg        [17:0]   img_reg_array_22_8_real;
  reg        [17:0]   img_reg_array_22_8_imag;
  reg        [17:0]   img_reg_array_22_9_real;
  reg        [17:0]   img_reg_array_22_9_imag;
  reg        [17:0]   img_reg_array_22_10_real;
  reg        [17:0]   img_reg_array_22_10_imag;
  reg        [17:0]   img_reg_array_22_11_real;
  reg        [17:0]   img_reg_array_22_11_imag;
  reg        [17:0]   img_reg_array_22_12_real;
  reg        [17:0]   img_reg_array_22_12_imag;
  reg        [17:0]   img_reg_array_22_13_real;
  reg        [17:0]   img_reg_array_22_13_imag;
  reg        [17:0]   img_reg_array_22_14_real;
  reg        [17:0]   img_reg_array_22_14_imag;
  reg        [17:0]   img_reg_array_22_15_real;
  reg        [17:0]   img_reg_array_22_15_imag;
  reg        [17:0]   img_reg_array_22_16_real;
  reg        [17:0]   img_reg_array_22_16_imag;
  reg        [17:0]   img_reg_array_22_17_real;
  reg        [17:0]   img_reg_array_22_17_imag;
  reg        [17:0]   img_reg_array_22_18_real;
  reg        [17:0]   img_reg_array_22_18_imag;
  reg        [17:0]   img_reg_array_22_19_real;
  reg        [17:0]   img_reg_array_22_19_imag;
  reg        [17:0]   img_reg_array_22_20_real;
  reg        [17:0]   img_reg_array_22_20_imag;
  reg        [17:0]   img_reg_array_22_21_real;
  reg        [17:0]   img_reg_array_22_21_imag;
  reg        [17:0]   img_reg_array_22_22_real;
  reg        [17:0]   img_reg_array_22_22_imag;
  reg        [17:0]   img_reg_array_22_23_real;
  reg        [17:0]   img_reg_array_22_23_imag;
  reg        [17:0]   img_reg_array_22_24_real;
  reg        [17:0]   img_reg_array_22_24_imag;
  reg        [17:0]   img_reg_array_22_25_real;
  reg        [17:0]   img_reg_array_22_25_imag;
  reg        [17:0]   img_reg_array_22_26_real;
  reg        [17:0]   img_reg_array_22_26_imag;
  reg        [17:0]   img_reg_array_22_27_real;
  reg        [17:0]   img_reg_array_22_27_imag;
  reg        [17:0]   img_reg_array_22_28_real;
  reg        [17:0]   img_reg_array_22_28_imag;
  reg        [17:0]   img_reg_array_22_29_real;
  reg        [17:0]   img_reg_array_22_29_imag;
  reg        [17:0]   img_reg_array_22_30_real;
  reg        [17:0]   img_reg_array_22_30_imag;
  reg        [17:0]   img_reg_array_22_31_real;
  reg        [17:0]   img_reg_array_22_31_imag;
  reg        [17:0]   img_reg_array_22_32_real;
  reg        [17:0]   img_reg_array_22_32_imag;
  reg        [17:0]   img_reg_array_22_33_real;
  reg        [17:0]   img_reg_array_22_33_imag;
  reg        [17:0]   img_reg_array_22_34_real;
  reg        [17:0]   img_reg_array_22_34_imag;
  reg        [17:0]   img_reg_array_22_35_real;
  reg        [17:0]   img_reg_array_22_35_imag;
  reg        [17:0]   img_reg_array_22_36_real;
  reg        [17:0]   img_reg_array_22_36_imag;
  reg        [17:0]   img_reg_array_22_37_real;
  reg        [17:0]   img_reg_array_22_37_imag;
  reg        [17:0]   img_reg_array_22_38_real;
  reg        [17:0]   img_reg_array_22_38_imag;
  reg        [17:0]   img_reg_array_22_39_real;
  reg        [17:0]   img_reg_array_22_39_imag;
  reg        [17:0]   img_reg_array_22_40_real;
  reg        [17:0]   img_reg_array_22_40_imag;
  reg        [17:0]   img_reg_array_22_41_real;
  reg        [17:0]   img_reg_array_22_41_imag;
  reg        [17:0]   img_reg_array_22_42_real;
  reg        [17:0]   img_reg_array_22_42_imag;
  reg        [17:0]   img_reg_array_22_43_real;
  reg        [17:0]   img_reg_array_22_43_imag;
  reg        [17:0]   img_reg_array_22_44_real;
  reg        [17:0]   img_reg_array_22_44_imag;
  reg        [17:0]   img_reg_array_22_45_real;
  reg        [17:0]   img_reg_array_22_45_imag;
  reg        [17:0]   img_reg_array_22_46_real;
  reg        [17:0]   img_reg_array_22_46_imag;
  reg        [17:0]   img_reg_array_22_47_real;
  reg        [17:0]   img_reg_array_22_47_imag;
  reg        [17:0]   img_reg_array_22_48_real;
  reg        [17:0]   img_reg_array_22_48_imag;
  reg        [17:0]   img_reg_array_22_49_real;
  reg        [17:0]   img_reg_array_22_49_imag;
  reg        [17:0]   img_reg_array_22_50_real;
  reg        [17:0]   img_reg_array_22_50_imag;
  reg        [17:0]   img_reg_array_22_51_real;
  reg        [17:0]   img_reg_array_22_51_imag;
  reg        [17:0]   img_reg_array_22_52_real;
  reg        [17:0]   img_reg_array_22_52_imag;
  reg        [17:0]   img_reg_array_22_53_real;
  reg        [17:0]   img_reg_array_22_53_imag;
  reg        [17:0]   img_reg_array_22_54_real;
  reg        [17:0]   img_reg_array_22_54_imag;
  reg        [17:0]   img_reg_array_22_55_real;
  reg        [17:0]   img_reg_array_22_55_imag;
  reg        [17:0]   img_reg_array_22_56_real;
  reg        [17:0]   img_reg_array_22_56_imag;
  reg        [17:0]   img_reg_array_22_57_real;
  reg        [17:0]   img_reg_array_22_57_imag;
  reg        [17:0]   img_reg_array_22_58_real;
  reg        [17:0]   img_reg_array_22_58_imag;
  reg        [17:0]   img_reg_array_22_59_real;
  reg        [17:0]   img_reg_array_22_59_imag;
  reg        [17:0]   img_reg_array_22_60_real;
  reg        [17:0]   img_reg_array_22_60_imag;
  reg        [17:0]   img_reg_array_22_61_real;
  reg        [17:0]   img_reg_array_22_61_imag;
  reg        [17:0]   img_reg_array_22_62_real;
  reg        [17:0]   img_reg_array_22_62_imag;
  reg        [17:0]   img_reg_array_22_63_real;
  reg        [17:0]   img_reg_array_22_63_imag;
  reg        [17:0]   img_reg_array_23_0_real;
  reg        [17:0]   img_reg_array_23_0_imag;
  reg        [17:0]   img_reg_array_23_1_real;
  reg        [17:0]   img_reg_array_23_1_imag;
  reg        [17:0]   img_reg_array_23_2_real;
  reg        [17:0]   img_reg_array_23_2_imag;
  reg        [17:0]   img_reg_array_23_3_real;
  reg        [17:0]   img_reg_array_23_3_imag;
  reg        [17:0]   img_reg_array_23_4_real;
  reg        [17:0]   img_reg_array_23_4_imag;
  reg        [17:0]   img_reg_array_23_5_real;
  reg        [17:0]   img_reg_array_23_5_imag;
  reg        [17:0]   img_reg_array_23_6_real;
  reg        [17:0]   img_reg_array_23_6_imag;
  reg        [17:0]   img_reg_array_23_7_real;
  reg        [17:0]   img_reg_array_23_7_imag;
  reg        [17:0]   img_reg_array_23_8_real;
  reg        [17:0]   img_reg_array_23_8_imag;
  reg        [17:0]   img_reg_array_23_9_real;
  reg        [17:0]   img_reg_array_23_9_imag;
  reg        [17:0]   img_reg_array_23_10_real;
  reg        [17:0]   img_reg_array_23_10_imag;
  reg        [17:0]   img_reg_array_23_11_real;
  reg        [17:0]   img_reg_array_23_11_imag;
  reg        [17:0]   img_reg_array_23_12_real;
  reg        [17:0]   img_reg_array_23_12_imag;
  reg        [17:0]   img_reg_array_23_13_real;
  reg        [17:0]   img_reg_array_23_13_imag;
  reg        [17:0]   img_reg_array_23_14_real;
  reg        [17:0]   img_reg_array_23_14_imag;
  reg        [17:0]   img_reg_array_23_15_real;
  reg        [17:0]   img_reg_array_23_15_imag;
  reg        [17:0]   img_reg_array_23_16_real;
  reg        [17:0]   img_reg_array_23_16_imag;
  reg        [17:0]   img_reg_array_23_17_real;
  reg        [17:0]   img_reg_array_23_17_imag;
  reg        [17:0]   img_reg_array_23_18_real;
  reg        [17:0]   img_reg_array_23_18_imag;
  reg        [17:0]   img_reg_array_23_19_real;
  reg        [17:0]   img_reg_array_23_19_imag;
  reg        [17:0]   img_reg_array_23_20_real;
  reg        [17:0]   img_reg_array_23_20_imag;
  reg        [17:0]   img_reg_array_23_21_real;
  reg        [17:0]   img_reg_array_23_21_imag;
  reg        [17:0]   img_reg_array_23_22_real;
  reg        [17:0]   img_reg_array_23_22_imag;
  reg        [17:0]   img_reg_array_23_23_real;
  reg        [17:0]   img_reg_array_23_23_imag;
  reg        [17:0]   img_reg_array_23_24_real;
  reg        [17:0]   img_reg_array_23_24_imag;
  reg        [17:0]   img_reg_array_23_25_real;
  reg        [17:0]   img_reg_array_23_25_imag;
  reg        [17:0]   img_reg_array_23_26_real;
  reg        [17:0]   img_reg_array_23_26_imag;
  reg        [17:0]   img_reg_array_23_27_real;
  reg        [17:0]   img_reg_array_23_27_imag;
  reg        [17:0]   img_reg_array_23_28_real;
  reg        [17:0]   img_reg_array_23_28_imag;
  reg        [17:0]   img_reg_array_23_29_real;
  reg        [17:0]   img_reg_array_23_29_imag;
  reg        [17:0]   img_reg_array_23_30_real;
  reg        [17:0]   img_reg_array_23_30_imag;
  reg        [17:0]   img_reg_array_23_31_real;
  reg        [17:0]   img_reg_array_23_31_imag;
  reg        [17:0]   img_reg_array_23_32_real;
  reg        [17:0]   img_reg_array_23_32_imag;
  reg        [17:0]   img_reg_array_23_33_real;
  reg        [17:0]   img_reg_array_23_33_imag;
  reg        [17:0]   img_reg_array_23_34_real;
  reg        [17:0]   img_reg_array_23_34_imag;
  reg        [17:0]   img_reg_array_23_35_real;
  reg        [17:0]   img_reg_array_23_35_imag;
  reg        [17:0]   img_reg_array_23_36_real;
  reg        [17:0]   img_reg_array_23_36_imag;
  reg        [17:0]   img_reg_array_23_37_real;
  reg        [17:0]   img_reg_array_23_37_imag;
  reg        [17:0]   img_reg_array_23_38_real;
  reg        [17:0]   img_reg_array_23_38_imag;
  reg        [17:0]   img_reg_array_23_39_real;
  reg        [17:0]   img_reg_array_23_39_imag;
  reg        [17:0]   img_reg_array_23_40_real;
  reg        [17:0]   img_reg_array_23_40_imag;
  reg        [17:0]   img_reg_array_23_41_real;
  reg        [17:0]   img_reg_array_23_41_imag;
  reg        [17:0]   img_reg_array_23_42_real;
  reg        [17:0]   img_reg_array_23_42_imag;
  reg        [17:0]   img_reg_array_23_43_real;
  reg        [17:0]   img_reg_array_23_43_imag;
  reg        [17:0]   img_reg_array_23_44_real;
  reg        [17:0]   img_reg_array_23_44_imag;
  reg        [17:0]   img_reg_array_23_45_real;
  reg        [17:0]   img_reg_array_23_45_imag;
  reg        [17:0]   img_reg_array_23_46_real;
  reg        [17:0]   img_reg_array_23_46_imag;
  reg        [17:0]   img_reg_array_23_47_real;
  reg        [17:0]   img_reg_array_23_47_imag;
  reg        [17:0]   img_reg_array_23_48_real;
  reg        [17:0]   img_reg_array_23_48_imag;
  reg        [17:0]   img_reg_array_23_49_real;
  reg        [17:0]   img_reg_array_23_49_imag;
  reg        [17:0]   img_reg_array_23_50_real;
  reg        [17:0]   img_reg_array_23_50_imag;
  reg        [17:0]   img_reg_array_23_51_real;
  reg        [17:0]   img_reg_array_23_51_imag;
  reg        [17:0]   img_reg_array_23_52_real;
  reg        [17:0]   img_reg_array_23_52_imag;
  reg        [17:0]   img_reg_array_23_53_real;
  reg        [17:0]   img_reg_array_23_53_imag;
  reg        [17:0]   img_reg_array_23_54_real;
  reg        [17:0]   img_reg_array_23_54_imag;
  reg        [17:0]   img_reg_array_23_55_real;
  reg        [17:0]   img_reg_array_23_55_imag;
  reg        [17:0]   img_reg_array_23_56_real;
  reg        [17:0]   img_reg_array_23_56_imag;
  reg        [17:0]   img_reg_array_23_57_real;
  reg        [17:0]   img_reg_array_23_57_imag;
  reg        [17:0]   img_reg_array_23_58_real;
  reg        [17:0]   img_reg_array_23_58_imag;
  reg        [17:0]   img_reg_array_23_59_real;
  reg        [17:0]   img_reg_array_23_59_imag;
  reg        [17:0]   img_reg_array_23_60_real;
  reg        [17:0]   img_reg_array_23_60_imag;
  reg        [17:0]   img_reg_array_23_61_real;
  reg        [17:0]   img_reg_array_23_61_imag;
  reg        [17:0]   img_reg_array_23_62_real;
  reg        [17:0]   img_reg_array_23_62_imag;
  reg        [17:0]   img_reg_array_23_63_real;
  reg        [17:0]   img_reg_array_23_63_imag;
  reg        [17:0]   img_reg_array_24_0_real;
  reg        [17:0]   img_reg_array_24_0_imag;
  reg        [17:0]   img_reg_array_24_1_real;
  reg        [17:0]   img_reg_array_24_1_imag;
  reg        [17:0]   img_reg_array_24_2_real;
  reg        [17:0]   img_reg_array_24_2_imag;
  reg        [17:0]   img_reg_array_24_3_real;
  reg        [17:0]   img_reg_array_24_3_imag;
  reg        [17:0]   img_reg_array_24_4_real;
  reg        [17:0]   img_reg_array_24_4_imag;
  reg        [17:0]   img_reg_array_24_5_real;
  reg        [17:0]   img_reg_array_24_5_imag;
  reg        [17:0]   img_reg_array_24_6_real;
  reg        [17:0]   img_reg_array_24_6_imag;
  reg        [17:0]   img_reg_array_24_7_real;
  reg        [17:0]   img_reg_array_24_7_imag;
  reg        [17:0]   img_reg_array_24_8_real;
  reg        [17:0]   img_reg_array_24_8_imag;
  reg        [17:0]   img_reg_array_24_9_real;
  reg        [17:0]   img_reg_array_24_9_imag;
  reg        [17:0]   img_reg_array_24_10_real;
  reg        [17:0]   img_reg_array_24_10_imag;
  reg        [17:0]   img_reg_array_24_11_real;
  reg        [17:0]   img_reg_array_24_11_imag;
  reg        [17:0]   img_reg_array_24_12_real;
  reg        [17:0]   img_reg_array_24_12_imag;
  reg        [17:0]   img_reg_array_24_13_real;
  reg        [17:0]   img_reg_array_24_13_imag;
  reg        [17:0]   img_reg_array_24_14_real;
  reg        [17:0]   img_reg_array_24_14_imag;
  reg        [17:0]   img_reg_array_24_15_real;
  reg        [17:0]   img_reg_array_24_15_imag;
  reg        [17:0]   img_reg_array_24_16_real;
  reg        [17:0]   img_reg_array_24_16_imag;
  reg        [17:0]   img_reg_array_24_17_real;
  reg        [17:0]   img_reg_array_24_17_imag;
  reg        [17:0]   img_reg_array_24_18_real;
  reg        [17:0]   img_reg_array_24_18_imag;
  reg        [17:0]   img_reg_array_24_19_real;
  reg        [17:0]   img_reg_array_24_19_imag;
  reg        [17:0]   img_reg_array_24_20_real;
  reg        [17:0]   img_reg_array_24_20_imag;
  reg        [17:0]   img_reg_array_24_21_real;
  reg        [17:0]   img_reg_array_24_21_imag;
  reg        [17:0]   img_reg_array_24_22_real;
  reg        [17:0]   img_reg_array_24_22_imag;
  reg        [17:0]   img_reg_array_24_23_real;
  reg        [17:0]   img_reg_array_24_23_imag;
  reg        [17:0]   img_reg_array_24_24_real;
  reg        [17:0]   img_reg_array_24_24_imag;
  reg        [17:0]   img_reg_array_24_25_real;
  reg        [17:0]   img_reg_array_24_25_imag;
  reg        [17:0]   img_reg_array_24_26_real;
  reg        [17:0]   img_reg_array_24_26_imag;
  reg        [17:0]   img_reg_array_24_27_real;
  reg        [17:0]   img_reg_array_24_27_imag;
  reg        [17:0]   img_reg_array_24_28_real;
  reg        [17:0]   img_reg_array_24_28_imag;
  reg        [17:0]   img_reg_array_24_29_real;
  reg        [17:0]   img_reg_array_24_29_imag;
  reg        [17:0]   img_reg_array_24_30_real;
  reg        [17:0]   img_reg_array_24_30_imag;
  reg        [17:0]   img_reg_array_24_31_real;
  reg        [17:0]   img_reg_array_24_31_imag;
  reg        [17:0]   img_reg_array_24_32_real;
  reg        [17:0]   img_reg_array_24_32_imag;
  reg        [17:0]   img_reg_array_24_33_real;
  reg        [17:0]   img_reg_array_24_33_imag;
  reg        [17:0]   img_reg_array_24_34_real;
  reg        [17:0]   img_reg_array_24_34_imag;
  reg        [17:0]   img_reg_array_24_35_real;
  reg        [17:0]   img_reg_array_24_35_imag;
  reg        [17:0]   img_reg_array_24_36_real;
  reg        [17:0]   img_reg_array_24_36_imag;
  reg        [17:0]   img_reg_array_24_37_real;
  reg        [17:0]   img_reg_array_24_37_imag;
  reg        [17:0]   img_reg_array_24_38_real;
  reg        [17:0]   img_reg_array_24_38_imag;
  reg        [17:0]   img_reg_array_24_39_real;
  reg        [17:0]   img_reg_array_24_39_imag;
  reg        [17:0]   img_reg_array_24_40_real;
  reg        [17:0]   img_reg_array_24_40_imag;
  reg        [17:0]   img_reg_array_24_41_real;
  reg        [17:0]   img_reg_array_24_41_imag;
  reg        [17:0]   img_reg_array_24_42_real;
  reg        [17:0]   img_reg_array_24_42_imag;
  reg        [17:0]   img_reg_array_24_43_real;
  reg        [17:0]   img_reg_array_24_43_imag;
  reg        [17:0]   img_reg_array_24_44_real;
  reg        [17:0]   img_reg_array_24_44_imag;
  reg        [17:0]   img_reg_array_24_45_real;
  reg        [17:0]   img_reg_array_24_45_imag;
  reg        [17:0]   img_reg_array_24_46_real;
  reg        [17:0]   img_reg_array_24_46_imag;
  reg        [17:0]   img_reg_array_24_47_real;
  reg        [17:0]   img_reg_array_24_47_imag;
  reg        [17:0]   img_reg_array_24_48_real;
  reg        [17:0]   img_reg_array_24_48_imag;
  reg        [17:0]   img_reg_array_24_49_real;
  reg        [17:0]   img_reg_array_24_49_imag;
  reg        [17:0]   img_reg_array_24_50_real;
  reg        [17:0]   img_reg_array_24_50_imag;
  reg        [17:0]   img_reg_array_24_51_real;
  reg        [17:0]   img_reg_array_24_51_imag;
  reg        [17:0]   img_reg_array_24_52_real;
  reg        [17:0]   img_reg_array_24_52_imag;
  reg        [17:0]   img_reg_array_24_53_real;
  reg        [17:0]   img_reg_array_24_53_imag;
  reg        [17:0]   img_reg_array_24_54_real;
  reg        [17:0]   img_reg_array_24_54_imag;
  reg        [17:0]   img_reg_array_24_55_real;
  reg        [17:0]   img_reg_array_24_55_imag;
  reg        [17:0]   img_reg_array_24_56_real;
  reg        [17:0]   img_reg_array_24_56_imag;
  reg        [17:0]   img_reg_array_24_57_real;
  reg        [17:0]   img_reg_array_24_57_imag;
  reg        [17:0]   img_reg_array_24_58_real;
  reg        [17:0]   img_reg_array_24_58_imag;
  reg        [17:0]   img_reg_array_24_59_real;
  reg        [17:0]   img_reg_array_24_59_imag;
  reg        [17:0]   img_reg_array_24_60_real;
  reg        [17:0]   img_reg_array_24_60_imag;
  reg        [17:0]   img_reg_array_24_61_real;
  reg        [17:0]   img_reg_array_24_61_imag;
  reg        [17:0]   img_reg_array_24_62_real;
  reg        [17:0]   img_reg_array_24_62_imag;
  reg        [17:0]   img_reg_array_24_63_real;
  reg        [17:0]   img_reg_array_24_63_imag;
  reg        [17:0]   img_reg_array_25_0_real;
  reg        [17:0]   img_reg_array_25_0_imag;
  reg        [17:0]   img_reg_array_25_1_real;
  reg        [17:0]   img_reg_array_25_1_imag;
  reg        [17:0]   img_reg_array_25_2_real;
  reg        [17:0]   img_reg_array_25_2_imag;
  reg        [17:0]   img_reg_array_25_3_real;
  reg        [17:0]   img_reg_array_25_3_imag;
  reg        [17:0]   img_reg_array_25_4_real;
  reg        [17:0]   img_reg_array_25_4_imag;
  reg        [17:0]   img_reg_array_25_5_real;
  reg        [17:0]   img_reg_array_25_5_imag;
  reg        [17:0]   img_reg_array_25_6_real;
  reg        [17:0]   img_reg_array_25_6_imag;
  reg        [17:0]   img_reg_array_25_7_real;
  reg        [17:0]   img_reg_array_25_7_imag;
  reg        [17:0]   img_reg_array_25_8_real;
  reg        [17:0]   img_reg_array_25_8_imag;
  reg        [17:0]   img_reg_array_25_9_real;
  reg        [17:0]   img_reg_array_25_9_imag;
  reg        [17:0]   img_reg_array_25_10_real;
  reg        [17:0]   img_reg_array_25_10_imag;
  reg        [17:0]   img_reg_array_25_11_real;
  reg        [17:0]   img_reg_array_25_11_imag;
  reg        [17:0]   img_reg_array_25_12_real;
  reg        [17:0]   img_reg_array_25_12_imag;
  reg        [17:0]   img_reg_array_25_13_real;
  reg        [17:0]   img_reg_array_25_13_imag;
  reg        [17:0]   img_reg_array_25_14_real;
  reg        [17:0]   img_reg_array_25_14_imag;
  reg        [17:0]   img_reg_array_25_15_real;
  reg        [17:0]   img_reg_array_25_15_imag;
  reg        [17:0]   img_reg_array_25_16_real;
  reg        [17:0]   img_reg_array_25_16_imag;
  reg        [17:0]   img_reg_array_25_17_real;
  reg        [17:0]   img_reg_array_25_17_imag;
  reg        [17:0]   img_reg_array_25_18_real;
  reg        [17:0]   img_reg_array_25_18_imag;
  reg        [17:0]   img_reg_array_25_19_real;
  reg        [17:0]   img_reg_array_25_19_imag;
  reg        [17:0]   img_reg_array_25_20_real;
  reg        [17:0]   img_reg_array_25_20_imag;
  reg        [17:0]   img_reg_array_25_21_real;
  reg        [17:0]   img_reg_array_25_21_imag;
  reg        [17:0]   img_reg_array_25_22_real;
  reg        [17:0]   img_reg_array_25_22_imag;
  reg        [17:0]   img_reg_array_25_23_real;
  reg        [17:0]   img_reg_array_25_23_imag;
  reg        [17:0]   img_reg_array_25_24_real;
  reg        [17:0]   img_reg_array_25_24_imag;
  reg        [17:0]   img_reg_array_25_25_real;
  reg        [17:0]   img_reg_array_25_25_imag;
  reg        [17:0]   img_reg_array_25_26_real;
  reg        [17:0]   img_reg_array_25_26_imag;
  reg        [17:0]   img_reg_array_25_27_real;
  reg        [17:0]   img_reg_array_25_27_imag;
  reg        [17:0]   img_reg_array_25_28_real;
  reg        [17:0]   img_reg_array_25_28_imag;
  reg        [17:0]   img_reg_array_25_29_real;
  reg        [17:0]   img_reg_array_25_29_imag;
  reg        [17:0]   img_reg_array_25_30_real;
  reg        [17:0]   img_reg_array_25_30_imag;
  reg        [17:0]   img_reg_array_25_31_real;
  reg        [17:0]   img_reg_array_25_31_imag;
  reg        [17:0]   img_reg_array_25_32_real;
  reg        [17:0]   img_reg_array_25_32_imag;
  reg        [17:0]   img_reg_array_25_33_real;
  reg        [17:0]   img_reg_array_25_33_imag;
  reg        [17:0]   img_reg_array_25_34_real;
  reg        [17:0]   img_reg_array_25_34_imag;
  reg        [17:0]   img_reg_array_25_35_real;
  reg        [17:0]   img_reg_array_25_35_imag;
  reg        [17:0]   img_reg_array_25_36_real;
  reg        [17:0]   img_reg_array_25_36_imag;
  reg        [17:0]   img_reg_array_25_37_real;
  reg        [17:0]   img_reg_array_25_37_imag;
  reg        [17:0]   img_reg_array_25_38_real;
  reg        [17:0]   img_reg_array_25_38_imag;
  reg        [17:0]   img_reg_array_25_39_real;
  reg        [17:0]   img_reg_array_25_39_imag;
  reg        [17:0]   img_reg_array_25_40_real;
  reg        [17:0]   img_reg_array_25_40_imag;
  reg        [17:0]   img_reg_array_25_41_real;
  reg        [17:0]   img_reg_array_25_41_imag;
  reg        [17:0]   img_reg_array_25_42_real;
  reg        [17:0]   img_reg_array_25_42_imag;
  reg        [17:0]   img_reg_array_25_43_real;
  reg        [17:0]   img_reg_array_25_43_imag;
  reg        [17:0]   img_reg_array_25_44_real;
  reg        [17:0]   img_reg_array_25_44_imag;
  reg        [17:0]   img_reg_array_25_45_real;
  reg        [17:0]   img_reg_array_25_45_imag;
  reg        [17:0]   img_reg_array_25_46_real;
  reg        [17:0]   img_reg_array_25_46_imag;
  reg        [17:0]   img_reg_array_25_47_real;
  reg        [17:0]   img_reg_array_25_47_imag;
  reg        [17:0]   img_reg_array_25_48_real;
  reg        [17:0]   img_reg_array_25_48_imag;
  reg        [17:0]   img_reg_array_25_49_real;
  reg        [17:0]   img_reg_array_25_49_imag;
  reg        [17:0]   img_reg_array_25_50_real;
  reg        [17:0]   img_reg_array_25_50_imag;
  reg        [17:0]   img_reg_array_25_51_real;
  reg        [17:0]   img_reg_array_25_51_imag;
  reg        [17:0]   img_reg_array_25_52_real;
  reg        [17:0]   img_reg_array_25_52_imag;
  reg        [17:0]   img_reg_array_25_53_real;
  reg        [17:0]   img_reg_array_25_53_imag;
  reg        [17:0]   img_reg_array_25_54_real;
  reg        [17:0]   img_reg_array_25_54_imag;
  reg        [17:0]   img_reg_array_25_55_real;
  reg        [17:0]   img_reg_array_25_55_imag;
  reg        [17:0]   img_reg_array_25_56_real;
  reg        [17:0]   img_reg_array_25_56_imag;
  reg        [17:0]   img_reg_array_25_57_real;
  reg        [17:0]   img_reg_array_25_57_imag;
  reg        [17:0]   img_reg_array_25_58_real;
  reg        [17:0]   img_reg_array_25_58_imag;
  reg        [17:0]   img_reg_array_25_59_real;
  reg        [17:0]   img_reg_array_25_59_imag;
  reg        [17:0]   img_reg_array_25_60_real;
  reg        [17:0]   img_reg_array_25_60_imag;
  reg        [17:0]   img_reg_array_25_61_real;
  reg        [17:0]   img_reg_array_25_61_imag;
  reg        [17:0]   img_reg_array_25_62_real;
  reg        [17:0]   img_reg_array_25_62_imag;
  reg        [17:0]   img_reg_array_25_63_real;
  reg        [17:0]   img_reg_array_25_63_imag;
  reg        [17:0]   img_reg_array_26_0_real;
  reg        [17:0]   img_reg_array_26_0_imag;
  reg        [17:0]   img_reg_array_26_1_real;
  reg        [17:0]   img_reg_array_26_1_imag;
  reg        [17:0]   img_reg_array_26_2_real;
  reg        [17:0]   img_reg_array_26_2_imag;
  reg        [17:0]   img_reg_array_26_3_real;
  reg        [17:0]   img_reg_array_26_3_imag;
  reg        [17:0]   img_reg_array_26_4_real;
  reg        [17:0]   img_reg_array_26_4_imag;
  reg        [17:0]   img_reg_array_26_5_real;
  reg        [17:0]   img_reg_array_26_5_imag;
  reg        [17:0]   img_reg_array_26_6_real;
  reg        [17:0]   img_reg_array_26_6_imag;
  reg        [17:0]   img_reg_array_26_7_real;
  reg        [17:0]   img_reg_array_26_7_imag;
  reg        [17:0]   img_reg_array_26_8_real;
  reg        [17:0]   img_reg_array_26_8_imag;
  reg        [17:0]   img_reg_array_26_9_real;
  reg        [17:0]   img_reg_array_26_9_imag;
  reg        [17:0]   img_reg_array_26_10_real;
  reg        [17:0]   img_reg_array_26_10_imag;
  reg        [17:0]   img_reg_array_26_11_real;
  reg        [17:0]   img_reg_array_26_11_imag;
  reg        [17:0]   img_reg_array_26_12_real;
  reg        [17:0]   img_reg_array_26_12_imag;
  reg        [17:0]   img_reg_array_26_13_real;
  reg        [17:0]   img_reg_array_26_13_imag;
  reg        [17:0]   img_reg_array_26_14_real;
  reg        [17:0]   img_reg_array_26_14_imag;
  reg        [17:0]   img_reg_array_26_15_real;
  reg        [17:0]   img_reg_array_26_15_imag;
  reg        [17:0]   img_reg_array_26_16_real;
  reg        [17:0]   img_reg_array_26_16_imag;
  reg        [17:0]   img_reg_array_26_17_real;
  reg        [17:0]   img_reg_array_26_17_imag;
  reg        [17:0]   img_reg_array_26_18_real;
  reg        [17:0]   img_reg_array_26_18_imag;
  reg        [17:0]   img_reg_array_26_19_real;
  reg        [17:0]   img_reg_array_26_19_imag;
  reg        [17:0]   img_reg_array_26_20_real;
  reg        [17:0]   img_reg_array_26_20_imag;
  reg        [17:0]   img_reg_array_26_21_real;
  reg        [17:0]   img_reg_array_26_21_imag;
  reg        [17:0]   img_reg_array_26_22_real;
  reg        [17:0]   img_reg_array_26_22_imag;
  reg        [17:0]   img_reg_array_26_23_real;
  reg        [17:0]   img_reg_array_26_23_imag;
  reg        [17:0]   img_reg_array_26_24_real;
  reg        [17:0]   img_reg_array_26_24_imag;
  reg        [17:0]   img_reg_array_26_25_real;
  reg        [17:0]   img_reg_array_26_25_imag;
  reg        [17:0]   img_reg_array_26_26_real;
  reg        [17:0]   img_reg_array_26_26_imag;
  reg        [17:0]   img_reg_array_26_27_real;
  reg        [17:0]   img_reg_array_26_27_imag;
  reg        [17:0]   img_reg_array_26_28_real;
  reg        [17:0]   img_reg_array_26_28_imag;
  reg        [17:0]   img_reg_array_26_29_real;
  reg        [17:0]   img_reg_array_26_29_imag;
  reg        [17:0]   img_reg_array_26_30_real;
  reg        [17:0]   img_reg_array_26_30_imag;
  reg        [17:0]   img_reg_array_26_31_real;
  reg        [17:0]   img_reg_array_26_31_imag;
  reg        [17:0]   img_reg_array_26_32_real;
  reg        [17:0]   img_reg_array_26_32_imag;
  reg        [17:0]   img_reg_array_26_33_real;
  reg        [17:0]   img_reg_array_26_33_imag;
  reg        [17:0]   img_reg_array_26_34_real;
  reg        [17:0]   img_reg_array_26_34_imag;
  reg        [17:0]   img_reg_array_26_35_real;
  reg        [17:0]   img_reg_array_26_35_imag;
  reg        [17:0]   img_reg_array_26_36_real;
  reg        [17:0]   img_reg_array_26_36_imag;
  reg        [17:0]   img_reg_array_26_37_real;
  reg        [17:0]   img_reg_array_26_37_imag;
  reg        [17:0]   img_reg_array_26_38_real;
  reg        [17:0]   img_reg_array_26_38_imag;
  reg        [17:0]   img_reg_array_26_39_real;
  reg        [17:0]   img_reg_array_26_39_imag;
  reg        [17:0]   img_reg_array_26_40_real;
  reg        [17:0]   img_reg_array_26_40_imag;
  reg        [17:0]   img_reg_array_26_41_real;
  reg        [17:0]   img_reg_array_26_41_imag;
  reg        [17:0]   img_reg_array_26_42_real;
  reg        [17:0]   img_reg_array_26_42_imag;
  reg        [17:0]   img_reg_array_26_43_real;
  reg        [17:0]   img_reg_array_26_43_imag;
  reg        [17:0]   img_reg_array_26_44_real;
  reg        [17:0]   img_reg_array_26_44_imag;
  reg        [17:0]   img_reg_array_26_45_real;
  reg        [17:0]   img_reg_array_26_45_imag;
  reg        [17:0]   img_reg_array_26_46_real;
  reg        [17:0]   img_reg_array_26_46_imag;
  reg        [17:0]   img_reg_array_26_47_real;
  reg        [17:0]   img_reg_array_26_47_imag;
  reg        [17:0]   img_reg_array_26_48_real;
  reg        [17:0]   img_reg_array_26_48_imag;
  reg        [17:0]   img_reg_array_26_49_real;
  reg        [17:0]   img_reg_array_26_49_imag;
  reg        [17:0]   img_reg_array_26_50_real;
  reg        [17:0]   img_reg_array_26_50_imag;
  reg        [17:0]   img_reg_array_26_51_real;
  reg        [17:0]   img_reg_array_26_51_imag;
  reg        [17:0]   img_reg_array_26_52_real;
  reg        [17:0]   img_reg_array_26_52_imag;
  reg        [17:0]   img_reg_array_26_53_real;
  reg        [17:0]   img_reg_array_26_53_imag;
  reg        [17:0]   img_reg_array_26_54_real;
  reg        [17:0]   img_reg_array_26_54_imag;
  reg        [17:0]   img_reg_array_26_55_real;
  reg        [17:0]   img_reg_array_26_55_imag;
  reg        [17:0]   img_reg_array_26_56_real;
  reg        [17:0]   img_reg_array_26_56_imag;
  reg        [17:0]   img_reg_array_26_57_real;
  reg        [17:0]   img_reg_array_26_57_imag;
  reg        [17:0]   img_reg_array_26_58_real;
  reg        [17:0]   img_reg_array_26_58_imag;
  reg        [17:0]   img_reg_array_26_59_real;
  reg        [17:0]   img_reg_array_26_59_imag;
  reg        [17:0]   img_reg_array_26_60_real;
  reg        [17:0]   img_reg_array_26_60_imag;
  reg        [17:0]   img_reg_array_26_61_real;
  reg        [17:0]   img_reg_array_26_61_imag;
  reg        [17:0]   img_reg_array_26_62_real;
  reg        [17:0]   img_reg_array_26_62_imag;
  reg        [17:0]   img_reg_array_26_63_real;
  reg        [17:0]   img_reg_array_26_63_imag;
  reg        [17:0]   img_reg_array_27_0_real;
  reg        [17:0]   img_reg_array_27_0_imag;
  reg        [17:0]   img_reg_array_27_1_real;
  reg        [17:0]   img_reg_array_27_1_imag;
  reg        [17:0]   img_reg_array_27_2_real;
  reg        [17:0]   img_reg_array_27_2_imag;
  reg        [17:0]   img_reg_array_27_3_real;
  reg        [17:0]   img_reg_array_27_3_imag;
  reg        [17:0]   img_reg_array_27_4_real;
  reg        [17:0]   img_reg_array_27_4_imag;
  reg        [17:0]   img_reg_array_27_5_real;
  reg        [17:0]   img_reg_array_27_5_imag;
  reg        [17:0]   img_reg_array_27_6_real;
  reg        [17:0]   img_reg_array_27_6_imag;
  reg        [17:0]   img_reg_array_27_7_real;
  reg        [17:0]   img_reg_array_27_7_imag;
  reg        [17:0]   img_reg_array_27_8_real;
  reg        [17:0]   img_reg_array_27_8_imag;
  reg        [17:0]   img_reg_array_27_9_real;
  reg        [17:0]   img_reg_array_27_9_imag;
  reg        [17:0]   img_reg_array_27_10_real;
  reg        [17:0]   img_reg_array_27_10_imag;
  reg        [17:0]   img_reg_array_27_11_real;
  reg        [17:0]   img_reg_array_27_11_imag;
  reg        [17:0]   img_reg_array_27_12_real;
  reg        [17:0]   img_reg_array_27_12_imag;
  reg        [17:0]   img_reg_array_27_13_real;
  reg        [17:0]   img_reg_array_27_13_imag;
  reg        [17:0]   img_reg_array_27_14_real;
  reg        [17:0]   img_reg_array_27_14_imag;
  reg        [17:0]   img_reg_array_27_15_real;
  reg        [17:0]   img_reg_array_27_15_imag;
  reg        [17:0]   img_reg_array_27_16_real;
  reg        [17:0]   img_reg_array_27_16_imag;
  reg        [17:0]   img_reg_array_27_17_real;
  reg        [17:0]   img_reg_array_27_17_imag;
  reg        [17:0]   img_reg_array_27_18_real;
  reg        [17:0]   img_reg_array_27_18_imag;
  reg        [17:0]   img_reg_array_27_19_real;
  reg        [17:0]   img_reg_array_27_19_imag;
  reg        [17:0]   img_reg_array_27_20_real;
  reg        [17:0]   img_reg_array_27_20_imag;
  reg        [17:0]   img_reg_array_27_21_real;
  reg        [17:0]   img_reg_array_27_21_imag;
  reg        [17:0]   img_reg_array_27_22_real;
  reg        [17:0]   img_reg_array_27_22_imag;
  reg        [17:0]   img_reg_array_27_23_real;
  reg        [17:0]   img_reg_array_27_23_imag;
  reg        [17:0]   img_reg_array_27_24_real;
  reg        [17:0]   img_reg_array_27_24_imag;
  reg        [17:0]   img_reg_array_27_25_real;
  reg        [17:0]   img_reg_array_27_25_imag;
  reg        [17:0]   img_reg_array_27_26_real;
  reg        [17:0]   img_reg_array_27_26_imag;
  reg        [17:0]   img_reg_array_27_27_real;
  reg        [17:0]   img_reg_array_27_27_imag;
  reg        [17:0]   img_reg_array_27_28_real;
  reg        [17:0]   img_reg_array_27_28_imag;
  reg        [17:0]   img_reg_array_27_29_real;
  reg        [17:0]   img_reg_array_27_29_imag;
  reg        [17:0]   img_reg_array_27_30_real;
  reg        [17:0]   img_reg_array_27_30_imag;
  reg        [17:0]   img_reg_array_27_31_real;
  reg        [17:0]   img_reg_array_27_31_imag;
  reg        [17:0]   img_reg_array_27_32_real;
  reg        [17:0]   img_reg_array_27_32_imag;
  reg        [17:0]   img_reg_array_27_33_real;
  reg        [17:0]   img_reg_array_27_33_imag;
  reg        [17:0]   img_reg_array_27_34_real;
  reg        [17:0]   img_reg_array_27_34_imag;
  reg        [17:0]   img_reg_array_27_35_real;
  reg        [17:0]   img_reg_array_27_35_imag;
  reg        [17:0]   img_reg_array_27_36_real;
  reg        [17:0]   img_reg_array_27_36_imag;
  reg        [17:0]   img_reg_array_27_37_real;
  reg        [17:0]   img_reg_array_27_37_imag;
  reg        [17:0]   img_reg_array_27_38_real;
  reg        [17:0]   img_reg_array_27_38_imag;
  reg        [17:0]   img_reg_array_27_39_real;
  reg        [17:0]   img_reg_array_27_39_imag;
  reg        [17:0]   img_reg_array_27_40_real;
  reg        [17:0]   img_reg_array_27_40_imag;
  reg        [17:0]   img_reg_array_27_41_real;
  reg        [17:0]   img_reg_array_27_41_imag;
  reg        [17:0]   img_reg_array_27_42_real;
  reg        [17:0]   img_reg_array_27_42_imag;
  reg        [17:0]   img_reg_array_27_43_real;
  reg        [17:0]   img_reg_array_27_43_imag;
  reg        [17:0]   img_reg_array_27_44_real;
  reg        [17:0]   img_reg_array_27_44_imag;
  reg        [17:0]   img_reg_array_27_45_real;
  reg        [17:0]   img_reg_array_27_45_imag;
  reg        [17:0]   img_reg_array_27_46_real;
  reg        [17:0]   img_reg_array_27_46_imag;
  reg        [17:0]   img_reg_array_27_47_real;
  reg        [17:0]   img_reg_array_27_47_imag;
  reg        [17:0]   img_reg_array_27_48_real;
  reg        [17:0]   img_reg_array_27_48_imag;
  reg        [17:0]   img_reg_array_27_49_real;
  reg        [17:0]   img_reg_array_27_49_imag;
  reg        [17:0]   img_reg_array_27_50_real;
  reg        [17:0]   img_reg_array_27_50_imag;
  reg        [17:0]   img_reg_array_27_51_real;
  reg        [17:0]   img_reg_array_27_51_imag;
  reg        [17:0]   img_reg_array_27_52_real;
  reg        [17:0]   img_reg_array_27_52_imag;
  reg        [17:0]   img_reg_array_27_53_real;
  reg        [17:0]   img_reg_array_27_53_imag;
  reg        [17:0]   img_reg_array_27_54_real;
  reg        [17:0]   img_reg_array_27_54_imag;
  reg        [17:0]   img_reg_array_27_55_real;
  reg        [17:0]   img_reg_array_27_55_imag;
  reg        [17:0]   img_reg_array_27_56_real;
  reg        [17:0]   img_reg_array_27_56_imag;
  reg        [17:0]   img_reg_array_27_57_real;
  reg        [17:0]   img_reg_array_27_57_imag;
  reg        [17:0]   img_reg_array_27_58_real;
  reg        [17:0]   img_reg_array_27_58_imag;
  reg        [17:0]   img_reg_array_27_59_real;
  reg        [17:0]   img_reg_array_27_59_imag;
  reg        [17:0]   img_reg_array_27_60_real;
  reg        [17:0]   img_reg_array_27_60_imag;
  reg        [17:0]   img_reg_array_27_61_real;
  reg        [17:0]   img_reg_array_27_61_imag;
  reg        [17:0]   img_reg_array_27_62_real;
  reg        [17:0]   img_reg_array_27_62_imag;
  reg        [17:0]   img_reg_array_27_63_real;
  reg        [17:0]   img_reg_array_27_63_imag;
  reg        [17:0]   img_reg_array_28_0_real;
  reg        [17:0]   img_reg_array_28_0_imag;
  reg        [17:0]   img_reg_array_28_1_real;
  reg        [17:0]   img_reg_array_28_1_imag;
  reg        [17:0]   img_reg_array_28_2_real;
  reg        [17:0]   img_reg_array_28_2_imag;
  reg        [17:0]   img_reg_array_28_3_real;
  reg        [17:0]   img_reg_array_28_3_imag;
  reg        [17:0]   img_reg_array_28_4_real;
  reg        [17:0]   img_reg_array_28_4_imag;
  reg        [17:0]   img_reg_array_28_5_real;
  reg        [17:0]   img_reg_array_28_5_imag;
  reg        [17:0]   img_reg_array_28_6_real;
  reg        [17:0]   img_reg_array_28_6_imag;
  reg        [17:0]   img_reg_array_28_7_real;
  reg        [17:0]   img_reg_array_28_7_imag;
  reg        [17:0]   img_reg_array_28_8_real;
  reg        [17:0]   img_reg_array_28_8_imag;
  reg        [17:0]   img_reg_array_28_9_real;
  reg        [17:0]   img_reg_array_28_9_imag;
  reg        [17:0]   img_reg_array_28_10_real;
  reg        [17:0]   img_reg_array_28_10_imag;
  reg        [17:0]   img_reg_array_28_11_real;
  reg        [17:0]   img_reg_array_28_11_imag;
  reg        [17:0]   img_reg_array_28_12_real;
  reg        [17:0]   img_reg_array_28_12_imag;
  reg        [17:0]   img_reg_array_28_13_real;
  reg        [17:0]   img_reg_array_28_13_imag;
  reg        [17:0]   img_reg_array_28_14_real;
  reg        [17:0]   img_reg_array_28_14_imag;
  reg        [17:0]   img_reg_array_28_15_real;
  reg        [17:0]   img_reg_array_28_15_imag;
  reg        [17:0]   img_reg_array_28_16_real;
  reg        [17:0]   img_reg_array_28_16_imag;
  reg        [17:0]   img_reg_array_28_17_real;
  reg        [17:0]   img_reg_array_28_17_imag;
  reg        [17:0]   img_reg_array_28_18_real;
  reg        [17:0]   img_reg_array_28_18_imag;
  reg        [17:0]   img_reg_array_28_19_real;
  reg        [17:0]   img_reg_array_28_19_imag;
  reg        [17:0]   img_reg_array_28_20_real;
  reg        [17:0]   img_reg_array_28_20_imag;
  reg        [17:0]   img_reg_array_28_21_real;
  reg        [17:0]   img_reg_array_28_21_imag;
  reg        [17:0]   img_reg_array_28_22_real;
  reg        [17:0]   img_reg_array_28_22_imag;
  reg        [17:0]   img_reg_array_28_23_real;
  reg        [17:0]   img_reg_array_28_23_imag;
  reg        [17:0]   img_reg_array_28_24_real;
  reg        [17:0]   img_reg_array_28_24_imag;
  reg        [17:0]   img_reg_array_28_25_real;
  reg        [17:0]   img_reg_array_28_25_imag;
  reg        [17:0]   img_reg_array_28_26_real;
  reg        [17:0]   img_reg_array_28_26_imag;
  reg        [17:0]   img_reg_array_28_27_real;
  reg        [17:0]   img_reg_array_28_27_imag;
  reg        [17:0]   img_reg_array_28_28_real;
  reg        [17:0]   img_reg_array_28_28_imag;
  reg        [17:0]   img_reg_array_28_29_real;
  reg        [17:0]   img_reg_array_28_29_imag;
  reg        [17:0]   img_reg_array_28_30_real;
  reg        [17:0]   img_reg_array_28_30_imag;
  reg        [17:0]   img_reg_array_28_31_real;
  reg        [17:0]   img_reg_array_28_31_imag;
  reg        [17:0]   img_reg_array_28_32_real;
  reg        [17:0]   img_reg_array_28_32_imag;
  reg        [17:0]   img_reg_array_28_33_real;
  reg        [17:0]   img_reg_array_28_33_imag;
  reg        [17:0]   img_reg_array_28_34_real;
  reg        [17:0]   img_reg_array_28_34_imag;
  reg        [17:0]   img_reg_array_28_35_real;
  reg        [17:0]   img_reg_array_28_35_imag;
  reg        [17:0]   img_reg_array_28_36_real;
  reg        [17:0]   img_reg_array_28_36_imag;
  reg        [17:0]   img_reg_array_28_37_real;
  reg        [17:0]   img_reg_array_28_37_imag;
  reg        [17:0]   img_reg_array_28_38_real;
  reg        [17:0]   img_reg_array_28_38_imag;
  reg        [17:0]   img_reg_array_28_39_real;
  reg        [17:0]   img_reg_array_28_39_imag;
  reg        [17:0]   img_reg_array_28_40_real;
  reg        [17:0]   img_reg_array_28_40_imag;
  reg        [17:0]   img_reg_array_28_41_real;
  reg        [17:0]   img_reg_array_28_41_imag;
  reg        [17:0]   img_reg_array_28_42_real;
  reg        [17:0]   img_reg_array_28_42_imag;
  reg        [17:0]   img_reg_array_28_43_real;
  reg        [17:0]   img_reg_array_28_43_imag;
  reg        [17:0]   img_reg_array_28_44_real;
  reg        [17:0]   img_reg_array_28_44_imag;
  reg        [17:0]   img_reg_array_28_45_real;
  reg        [17:0]   img_reg_array_28_45_imag;
  reg        [17:0]   img_reg_array_28_46_real;
  reg        [17:0]   img_reg_array_28_46_imag;
  reg        [17:0]   img_reg_array_28_47_real;
  reg        [17:0]   img_reg_array_28_47_imag;
  reg        [17:0]   img_reg_array_28_48_real;
  reg        [17:0]   img_reg_array_28_48_imag;
  reg        [17:0]   img_reg_array_28_49_real;
  reg        [17:0]   img_reg_array_28_49_imag;
  reg        [17:0]   img_reg_array_28_50_real;
  reg        [17:0]   img_reg_array_28_50_imag;
  reg        [17:0]   img_reg_array_28_51_real;
  reg        [17:0]   img_reg_array_28_51_imag;
  reg        [17:0]   img_reg_array_28_52_real;
  reg        [17:0]   img_reg_array_28_52_imag;
  reg        [17:0]   img_reg_array_28_53_real;
  reg        [17:0]   img_reg_array_28_53_imag;
  reg        [17:0]   img_reg_array_28_54_real;
  reg        [17:0]   img_reg_array_28_54_imag;
  reg        [17:0]   img_reg_array_28_55_real;
  reg        [17:0]   img_reg_array_28_55_imag;
  reg        [17:0]   img_reg_array_28_56_real;
  reg        [17:0]   img_reg_array_28_56_imag;
  reg        [17:0]   img_reg_array_28_57_real;
  reg        [17:0]   img_reg_array_28_57_imag;
  reg        [17:0]   img_reg_array_28_58_real;
  reg        [17:0]   img_reg_array_28_58_imag;
  reg        [17:0]   img_reg_array_28_59_real;
  reg        [17:0]   img_reg_array_28_59_imag;
  reg        [17:0]   img_reg_array_28_60_real;
  reg        [17:0]   img_reg_array_28_60_imag;
  reg        [17:0]   img_reg_array_28_61_real;
  reg        [17:0]   img_reg_array_28_61_imag;
  reg        [17:0]   img_reg_array_28_62_real;
  reg        [17:0]   img_reg_array_28_62_imag;
  reg        [17:0]   img_reg_array_28_63_real;
  reg        [17:0]   img_reg_array_28_63_imag;
  reg        [17:0]   img_reg_array_29_0_real;
  reg        [17:0]   img_reg_array_29_0_imag;
  reg        [17:0]   img_reg_array_29_1_real;
  reg        [17:0]   img_reg_array_29_1_imag;
  reg        [17:0]   img_reg_array_29_2_real;
  reg        [17:0]   img_reg_array_29_2_imag;
  reg        [17:0]   img_reg_array_29_3_real;
  reg        [17:0]   img_reg_array_29_3_imag;
  reg        [17:0]   img_reg_array_29_4_real;
  reg        [17:0]   img_reg_array_29_4_imag;
  reg        [17:0]   img_reg_array_29_5_real;
  reg        [17:0]   img_reg_array_29_5_imag;
  reg        [17:0]   img_reg_array_29_6_real;
  reg        [17:0]   img_reg_array_29_6_imag;
  reg        [17:0]   img_reg_array_29_7_real;
  reg        [17:0]   img_reg_array_29_7_imag;
  reg        [17:0]   img_reg_array_29_8_real;
  reg        [17:0]   img_reg_array_29_8_imag;
  reg        [17:0]   img_reg_array_29_9_real;
  reg        [17:0]   img_reg_array_29_9_imag;
  reg        [17:0]   img_reg_array_29_10_real;
  reg        [17:0]   img_reg_array_29_10_imag;
  reg        [17:0]   img_reg_array_29_11_real;
  reg        [17:0]   img_reg_array_29_11_imag;
  reg        [17:0]   img_reg_array_29_12_real;
  reg        [17:0]   img_reg_array_29_12_imag;
  reg        [17:0]   img_reg_array_29_13_real;
  reg        [17:0]   img_reg_array_29_13_imag;
  reg        [17:0]   img_reg_array_29_14_real;
  reg        [17:0]   img_reg_array_29_14_imag;
  reg        [17:0]   img_reg_array_29_15_real;
  reg        [17:0]   img_reg_array_29_15_imag;
  reg        [17:0]   img_reg_array_29_16_real;
  reg        [17:0]   img_reg_array_29_16_imag;
  reg        [17:0]   img_reg_array_29_17_real;
  reg        [17:0]   img_reg_array_29_17_imag;
  reg        [17:0]   img_reg_array_29_18_real;
  reg        [17:0]   img_reg_array_29_18_imag;
  reg        [17:0]   img_reg_array_29_19_real;
  reg        [17:0]   img_reg_array_29_19_imag;
  reg        [17:0]   img_reg_array_29_20_real;
  reg        [17:0]   img_reg_array_29_20_imag;
  reg        [17:0]   img_reg_array_29_21_real;
  reg        [17:0]   img_reg_array_29_21_imag;
  reg        [17:0]   img_reg_array_29_22_real;
  reg        [17:0]   img_reg_array_29_22_imag;
  reg        [17:0]   img_reg_array_29_23_real;
  reg        [17:0]   img_reg_array_29_23_imag;
  reg        [17:0]   img_reg_array_29_24_real;
  reg        [17:0]   img_reg_array_29_24_imag;
  reg        [17:0]   img_reg_array_29_25_real;
  reg        [17:0]   img_reg_array_29_25_imag;
  reg        [17:0]   img_reg_array_29_26_real;
  reg        [17:0]   img_reg_array_29_26_imag;
  reg        [17:0]   img_reg_array_29_27_real;
  reg        [17:0]   img_reg_array_29_27_imag;
  reg        [17:0]   img_reg_array_29_28_real;
  reg        [17:0]   img_reg_array_29_28_imag;
  reg        [17:0]   img_reg_array_29_29_real;
  reg        [17:0]   img_reg_array_29_29_imag;
  reg        [17:0]   img_reg_array_29_30_real;
  reg        [17:0]   img_reg_array_29_30_imag;
  reg        [17:0]   img_reg_array_29_31_real;
  reg        [17:0]   img_reg_array_29_31_imag;
  reg        [17:0]   img_reg_array_29_32_real;
  reg        [17:0]   img_reg_array_29_32_imag;
  reg        [17:0]   img_reg_array_29_33_real;
  reg        [17:0]   img_reg_array_29_33_imag;
  reg        [17:0]   img_reg_array_29_34_real;
  reg        [17:0]   img_reg_array_29_34_imag;
  reg        [17:0]   img_reg_array_29_35_real;
  reg        [17:0]   img_reg_array_29_35_imag;
  reg        [17:0]   img_reg_array_29_36_real;
  reg        [17:0]   img_reg_array_29_36_imag;
  reg        [17:0]   img_reg_array_29_37_real;
  reg        [17:0]   img_reg_array_29_37_imag;
  reg        [17:0]   img_reg_array_29_38_real;
  reg        [17:0]   img_reg_array_29_38_imag;
  reg        [17:0]   img_reg_array_29_39_real;
  reg        [17:0]   img_reg_array_29_39_imag;
  reg        [17:0]   img_reg_array_29_40_real;
  reg        [17:0]   img_reg_array_29_40_imag;
  reg        [17:0]   img_reg_array_29_41_real;
  reg        [17:0]   img_reg_array_29_41_imag;
  reg        [17:0]   img_reg_array_29_42_real;
  reg        [17:0]   img_reg_array_29_42_imag;
  reg        [17:0]   img_reg_array_29_43_real;
  reg        [17:0]   img_reg_array_29_43_imag;
  reg        [17:0]   img_reg_array_29_44_real;
  reg        [17:0]   img_reg_array_29_44_imag;
  reg        [17:0]   img_reg_array_29_45_real;
  reg        [17:0]   img_reg_array_29_45_imag;
  reg        [17:0]   img_reg_array_29_46_real;
  reg        [17:0]   img_reg_array_29_46_imag;
  reg        [17:0]   img_reg_array_29_47_real;
  reg        [17:0]   img_reg_array_29_47_imag;
  reg        [17:0]   img_reg_array_29_48_real;
  reg        [17:0]   img_reg_array_29_48_imag;
  reg        [17:0]   img_reg_array_29_49_real;
  reg        [17:0]   img_reg_array_29_49_imag;
  reg        [17:0]   img_reg_array_29_50_real;
  reg        [17:0]   img_reg_array_29_50_imag;
  reg        [17:0]   img_reg_array_29_51_real;
  reg        [17:0]   img_reg_array_29_51_imag;
  reg        [17:0]   img_reg_array_29_52_real;
  reg        [17:0]   img_reg_array_29_52_imag;
  reg        [17:0]   img_reg_array_29_53_real;
  reg        [17:0]   img_reg_array_29_53_imag;
  reg        [17:0]   img_reg_array_29_54_real;
  reg        [17:0]   img_reg_array_29_54_imag;
  reg        [17:0]   img_reg_array_29_55_real;
  reg        [17:0]   img_reg_array_29_55_imag;
  reg        [17:0]   img_reg_array_29_56_real;
  reg        [17:0]   img_reg_array_29_56_imag;
  reg        [17:0]   img_reg_array_29_57_real;
  reg        [17:0]   img_reg_array_29_57_imag;
  reg        [17:0]   img_reg_array_29_58_real;
  reg        [17:0]   img_reg_array_29_58_imag;
  reg        [17:0]   img_reg_array_29_59_real;
  reg        [17:0]   img_reg_array_29_59_imag;
  reg        [17:0]   img_reg_array_29_60_real;
  reg        [17:0]   img_reg_array_29_60_imag;
  reg        [17:0]   img_reg_array_29_61_real;
  reg        [17:0]   img_reg_array_29_61_imag;
  reg        [17:0]   img_reg_array_29_62_real;
  reg        [17:0]   img_reg_array_29_62_imag;
  reg        [17:0]   img_reg_array_29_63_real;
  reg        [17:0]   img_reg_array_29_63_imag;
  reg        [17:0]   img_reg_array_30_0_real;
  reg        [17:0]   img_reg_array_30_0_imag;
  reg        [17:0]   img_reg_array_30_1_real;
  reg        [17:0]   img_reg_array_30_1_imag;
  reg        [17:0]   img_reg_array_30_2_real;
  reg        [17:0]   img_reg_array_30_2_imag;
  reg        [17:0]   img_reg_array_30_3_real;
  reg        [17:0]   img_reg_array_30_3_imag;
  reg        [17:0]   img_reg_array_30_4_real;
  reg        [17:0]   img_reg_array_30_4_imag;
  reg        [17:0]   img_reg_array_30_5_real;
  reg        [17:0]   img_reg_array_30_5_imag;
  reg        [17:0]   img_reg_array_30_6_real;
  reg        [17:0]   img_reg_array_30_6_imag;
  reg        [17:0]   img_reg_array_30_7_real;
  reg        [17:0]   img_reg_array_30_7_imag;
  reg        [17:0]   img_reg_array_30_8_real;
  reg        [17:0]   img_reg_array_30_8_imag;
  reg        [17:0]   img_reg_array_30_9_real;
  reg        [17:0]   img_reg_array_30_9_imag;
  reg        [17:0]   img_reg_array_30_10_real;
  reg        [17:0]   img_reg_array_30_10_imag;
  reg        [17:0]   img_reg_array_30_11_real;
  reg        [17:0]   img_reg_array_30_11_imag;
  reg        [17:0]   img_reg_array_30_12_real;
  reg        [17:0]   img_reg_array_30_12_imag;
  reg        [17:0]   img_reg_array_30_13_real;
  reg        [17:0]   img_reg_array_30_13_imag;
  reg        [17:0]   img_reg_array_30_14_real;
  reg        [17:0]   img_reg_array_30_14_imag;
  reg        [17:0]   img_reg_array_30_15_real;
  reg        [17:0]   img_reg_array_30_15_imag;
  reg        [17:0]   img_reg_array_30_16_real;
  reg        [17:0]   img_reg_array_30_16_imag;
  reg        [17:0]   img_reg_array_30_17_real;
  reg        [17:0]   img_reg_array_30_17_imag;
  reg        [17:0]   img_reg_array_30_18_real;
  reg        [17:0]   img_reg_array_30_18_imag;
  reg        [17:0]   img_reg_array_30_19_real;
  reg        [17:0]   img_reg_array_30_19_imag;
  reg        [17:0]   img_reg_array_30_20_real;
  reg        [17:0]   img_reg_array_30_20_imag;
  reg        [17:0]   img_reg_array_30_21_real;
  reg        [17:0]   img_reg_array_30_21_imag;
  reg        [17:0]   img_reg_array_30_22_real;
  reg        [17:0]   img_reg_array_30_22_imag;
  reg        [17:0]   img_reg_array_30_23_real;
  reg        [17:0]   img_reg_array_30_23_imag;
  reg        [17:0]   img_reg_array_30_24_real;
  reg        [17:0]   img_reg_array_30_24_imag;
  reg        [17:0]   img_reg_array_30_25_real;
  reg        [17:0]   img_reg_array_30_25_imag;
  reg        [17:0]   img_reg_array_30_26_real;
  reg        [17:0]   img_reg_array_30_26_imag;
  reg        [17:0]   img_reg_array_30_27_real;
  reg        [17:0]   img_reg_array_30_27_imag;
  reg        [17:0]   img_reg_array_30_28_real;
  reg        [17:0]   img_reg_array_30_28_imag;
  reg        [17:0]   img_reg_array_30_29_real;
  reg        [17:0]   img_reg_array_30_29_imag;
  reg        [17:0]   img_reg_array_30_30_real;
  reg        [17:0]   img_reg_array_30_30_imag;
  reg        [17:0]   img_reg_array_30_31_real;
  reg        [17:0]   img_reg_array_30_31_imag;
  reg        [17:0]   img_reg_array_30_32_real;
  reg        [17:0]   img_reg_array_30_32_imag;
  reg        [17:0]   img_reg_array_30_33_real;
  reg        [17:0]   img_reg_array_30_33_imag;
  reg        [17:0]   img_reg_array_30_34_real;
  reg        [17:0]   img_reg_array_30_34_imag;
  reg        [17:0]   img_reg_array_30_35_real;
  reg        [17:0]   img_reg_array_30_35_imag;
  reg        [17:0]   img_reg_array_30_36_real;
  reg        [17:0]   img_reg_array_30_36_imag;
  reg        [17:0]   img_reg_array_30_37_real;
  reg        [17:0]   img_reg_array_30_37_imag;
  reg        [17:0]   img_reg_array_30_38_real;
  reg        [17:0]   img_reg_array_30_38_imag;
  reg        [17:0]   img_reg_array_30_39_real;
  reg        [17:0]   img_reg_array_30_39_imag;
  reg        [17:0]   img_reg_array_30_40_real;
  reg        [17:0]   img_reg_array_30_40_imag;
  reg        [17:0]   img_reg_array_30_41_real;
  reg        [17:0]   img_reg_array_30_41_imag;
  reg        [17:0]   img_reg_array_30_42_real;
  reg        [17:0]   img_reg_array_30_42_imag;
  reg        [17:0]   img_reg_array_30_43_real;
  reg        [17:0]   img_reg_array_30_43_imag;
  reg        [17:0]   img_reg_array_30_44_real;
  reg        [17:0]   img_reg_array_30_44_imag;
  reg        [17:0]   img_reg_array_30_45_real;
  reg        [17:0]   img_reg_array_30_45_imag;
  reg        [17:0]   img_reg_array_30_46_real;
  reg        [17:0]   img_reg_array_30_46_imag;
  reg        [17:0]   img_reg_array_30_47_real;
  reg        [17:0]   img_reg_array_30_47_imag;
  reg        [17:0]   img_reg_array_30_48_real;
  reg        [17:0]   img_reg_array_30_48_imag;
  reg        [17:0]   img_reg_array_30_49_real;
  reg        [17:0]   img_reg_array_30_49_imag;
  reg        [17:0]   img_reg_array_30_50_real;
  reg        [17:0]   img_reg_array_30_50_imag;
  reg        [17:0]   img_reg_array_30_51_real;
  reg        [17:0]   img_reg_array_30_51_imag;
  reg        [17:0]   img_reg_array_30_52_real;
  reg        [17:0]   img_reg_array_30_52_imag;
  reg        [17:0]   img_reg_array_30_53_real;
  reg        [17:0]   img_reg_array_30_53_imag;
  reg        [17:0]   img_reg_array_30_54_real;
  reg        [17:0]   img_reg_array_30_54_imag;
  reg        [17:0]   img_reg_array_30_55_real;
  reg        [17:0]   img_reg_array_30_55_imag;
  reg        [17:0]   img_reg_array_30_56_real;
  reg        [17:0]   img_reg_array_30_56_imag;
  reg        [17:0]   img_reg_array_30_57_real;
  reg        [17:0]   img_reg_array_30_57_imag;
  reg        [17:0]   img_reg_array_30_58_real;
  reg        [17:0]   img_reg_array_30_58_imag;
  reg        [17:0]   img_reg_array_30_59_real;
  reg        [17:0]   img_reg_array_30_59_imag;
  reg        [17:0]   img_reg_array_30_60_real;
  reg        [17:0]   img_reg_array_30_60_imag;
  reg        [17:0]   img_reg_array_30_61_real;
  reg        [17:0]   img_reg_array_30_61_imag;
  reg        [17:0]   img_reg_array_30_62_real;
  reg        [17:0]   img_reg_array_30_62_imag;
  reg        [17:0]   img_reg_array_30_63_real;
  reg        [17:0]   img_reg_array_30_63_imag;
  reg        [17:0]   img_reg_array_31_0_real;
  reg        [17:0]   img_reg_array_31_0_imag;
  reg        [17:0]   img_reg_array_31_1_real;
  reg        [17:0]   img_reg_array_31_1_imag;
  reg        [17:0]   img_reg_array_31_2_real;
  reg        [17:0]   img_reg_array_31_2_imag;
  reg        [17:0]   img_reg_array_31_3_real;
  reg        [17:0]   img_reg_array_31_3_imag;
  reg        [17:0]   img_reg_array_31_4_real;
  reg        [17:0]   img_reg_array_31_4_imag;
  reg        [17:0]   img_reg_array_31_5_real;
  reg        [17:0]   img_reg_array_31_5_imag;
  reg        [17:0]   img_reg_array_31_6_real;
  reg        [17:0]   img_reg_array_31_6_imag;
  reg        [17:0]   img_reg_array_31_7_real;
  reg        [17:0]   img_reg_array_31_7_imag;
  reg        [17:0]   img_reg_array_31_8_real;
  reg        [17:0]   img_reg_array_31_8_imag;
  reg        [17:0]   img_reg_array_31_9_real;
  reg        [17:0]   img_reg_array_31_9_imag;
  reg        [17:0]   img_reg_array_31_10_real;
  reg        [17:0]   img_reg_array_31_10_imag;
  reg        [17:0]   img_reg_array_31_11_real;
  reg        [17:0]   img_reg_array_31_11_imag;
  reg        [17:0]   img_reg_array_31_12_real;
  reg        [17:0]   img_reg_array_31_12_imag;
  reg        [17:0]   img_reg_array_31_13_real;
  reg        [17:0]   img_reg_array_31_13_imag;
  reg        [17:0]   img_reg_array_31_14_real;
  reg        [17:0]   img_reg_array_31_14_imag;
  reg        [17:0]   img_reg_array_31_15_real;
  reg        [17:0]   img_reg_array_31_15_imag;
  reg        [17:0]   img_reg_array_31_16_real;
  reg        [17:0]   img_reg_array_31_16_imag;
  reg        [17:0]   img_reg_array_31_17_real;
  reg        [17:0]   img_reg_array_31_17_imag;
  reg        [17:0]   img_reg_array_31_18_real;
  reg        [17:0]   img_reg_array_31_18_imag;
  reg        [17:0]   img_reg_array_31_19_real;
  reg        [17:0]   img_reg_array_31_19_imag;
  reg        [17:0]   img_reg_array_31_20_real;
  reg        [17:0]   img_reg_array_31_20_imag;
  reg        [17:0]   img_reg_array_31_21_real;
  reg        [17:0]   img_reg_array_31_21_imag;
  reg        [17:0]   img_reg_array_31_22_real;
  reg        [17:0]   img_reg_array_31_22_imag;
  reg        [17:0]   img_reg_array_31_23_real;
  reg        [17:0]   img_reg_array_31_23_imag;
  reg        [17:0]   img_reg_array_31_24_real;
  reg        [17:0]   img_reg_array_31_24_imag;
  reg        [17:0]   img_reg_array_31_25_real;
  reg        [17:0]   img_reg_array_31_25_imag;
  reg        [17:0]   img_reg_array_31_26_real;
  reg        [17:0]   img_reg_array_31_26_imag;
  reg        [17:0]   img_reg_array_31_27_real;
  reg        [17:0]   img_reg_array_31_27_imag;
  reg        [17:0]   img_reg_array_31_28_real;
  reg        [17:0]   img_reg_array_31_28_imag;
  reg        [17:0]   img_reg_array_31_29_real;
  reg        [17:0]   img_reg_array_31_29_imag;
  reg        [17:0]   img_reg_array_31_30_real;
  reg        [17:0]   img_reg_array_31_30_imag;
  reg        [17:0]   img_reg_array_31_31_real;
  reg        [17:0]   img_reg_array_31_31_imag;
  reg        [17:0]   img_reg_array_31_32_real;
  reg        [17:0]   img_reg_array_31_32_imag;
  reg        [17:0]   img_reg_array_31_33_real;
  reg        [17:0]   img_reg_array_31_33_imag;
  reg        [17:0]   img_reg_array_31_34_real;
  reg        [17:0]   img_reg_array_31_34_imag;
  reg        [17:0]   img_reg_array_31_35_real;
  reg        [17:0]   img_reg_array_31_35_imag;
  reg        [17:0]   img_reg_array_31_36_real;
  reg        [17:0]   img_reg_array_31_36_imag;
  reg        [17:0]   img_reg_array_31_37_real;
  reg        [17:0]   img_reg_array_31_37_imag;
  reg        [17:0]   img_reg_array_31_38_real;
  reg        [17:0]   img_reg_array_31_38_imag;
  reg        [17:0]   img_reg_array_31_39_real;
  reg        [17:0]   img_reg_array_31_39_imag;
  reg        [17:0]   img_reg_array_31_40_real;
  reg        [17:0]   img_reg_array_31_40_imag;
  reg        [17:0]   img_reg_array_31_41_real;
  reg        [17:0]   img_reg_array_31_41_imag;
  reg        [17:0]   img_reg_array_31_42_real;
  reg        [17:0]   img_reg_array_31_42_imag;
  reg        [17:0]   img_reg_array_31_43_real;
  reg        [17:0]   img_reg_array_31_43_imag;
  reg        [17:0]   img_reg_array_31_44_real;
  reg        [17:0]   img_reg_array_31_44_imag;
  reg        [17:0]   img_reg_array_31_45_real;
  reg        [17:0]   img_reg_array_31_45_imag;
  reg        [17:0]   img_reg_array_31_46_real;
  reg        [17:0]   img_reg_array_31_46_imag;
  reg        [17:0]   img_reg_array_31_47_real;
  reg        [17:0]   img_reg_array_31_47_imag;
  reg        [17:0]   img_reg_array_31_48_real;
  reg        [17:0]   img_reg_array_31_48_imag;
  reg        [17:0]   img_reg_array_31_49_real;
  reg        [17:0]   img_reg_array_31_49_imag;
  reg        [17:0]   img_reg_array_31_50_real;
  reg        [17:0]   img_reg_array_31_50_imag;
  reg        [17:0]   img_reg_array_31_51_real;
  reg        [17:0]   img_reg_array_31_51_imag;
  reg        [17:0]   img_reg_array_31_52_real;
  reg        [17:0]   img_reg_array_31_52_imag;
  reg        [17:0]   img_reg_array_31_53_real;
  reg        [17:0]   img_reg_array_31_53_imag;
  reg        [17:0]   img_reg_array_31_54_real;
  reg        [17:0]   img_reg_array_31_54_imag;
  reg        [17:0]   img_reg_array_31_55_real;
  reg        [17:0]   img_reg_array_31_55_imag;
  reg        [17:0]   img_reg_array_31_56_real;
  reg        [17:0]   img_reg_array_31_56_imag;
  reg        [17:0]   img_reg_array_31_57_real;
  reg        [17:0]   img_reg_array_31_57_imag;
  reg        [17:0]   img_reg_array_31_58_real;
  reg        [17:0]   img_reg_array_31_58_imag;
  reg        [17:0]   img_reg_array_31_59_real;
  reg        [17:0]   img_reg_array_31_59_imag;
  reg        [17:0]   img_reg_array_31_60_real;
  reg        [17:0]   img_reg_array_31_60_imag;
  reg        [17:0]   img_reg_array_31_61_real;
  reg        [17:0]   img_reg_array_31_61_imag;
  reg        [17:0]   img_reg_array_31_62_real;
  reg        [17:0]   img_reg_array_31_62_imag;
  reg        [17:0]   img_reg_array_31_63_real;
  reg        [17:0]   img_reg_array_31_63_imag;
  reg        [17:0]   img_reg_array_32_0_real;
  reg        [17:0]   img_reg_array_32_0_imag;
  reg        [17:0]   img_reg_array_32_1_real;
  reg        [17:0]   img_reg_array_32_1_imag;
  reg        [17:0]   img_reg_array_32_2_real;
  reg        [17:0]   img_reg_array_32_2_imag;
  reg        [17:0]   img_reg_array_32_3_real;
  reg        [17:0]   img_reg_array_32_3_imag;
  reg        [17:0]   img_reg_array_32_4_real;
  reg        [17:0]   img_reg_array_32_4_imag;
  reg        [17:0]   img_reg_array_32_5_real;
  reg        [17:0]   img_reg_array_32_5_imag;
  reg        [17:0]   img_reg_array_32_6_real;
  reg        [17:0]   img_reg_array_32_6_imag;
  reg        [17:0]   img_reg_array_32_7_real;
  reg        [17:0]   img_reg_array_32_7_imag;
  reg        [17:0]   img_reg_array_32_8_real;
  reg        [17:0]   img_reg_array_32_8_imag;
  reg        [17:0]   img_reg_array_32_9_real;
  reg        [17:0]   img_reg_array_32_9_imag;
  reg        [17:0]   img_reg_array_32_10_real;
  reg        [17:0]   img_reg_array_32_10_imag;
  reg        [17:0]   img_reg_array_32_11_real;
  reg        [17:0]   img_reg_array_32_11_imag;
  reg        [17:0]   img_reg_array_32_12_real;
  reg        [17:0]   img_reg_array_32_12_imag;
  reg        [17:0]   img_reg_array_32_13_real;
  reg        [17:0]   img_reg_array_32_13_imag;
  reg        [17:0]   img_reg_array_32_14_real;
  reg        [17:0]   img_reg_array_32_14_imag;
  reg        [17:0]   img_reg_array_32_15_real;
  reg        [17:0]   img_reg_array_32_15_imag;
  reg        [17:0]   img_reg_array_32_16_real;
  reg        [17:0]   img_reg_array_32_16_imag;
  reg        [17:0]   img_reg_array_32_17_real;
  reg        [17:0]   img_reg_array_32_17_imag;
  reg        [17:0]   img_reg_array_32_18_real;
  reg        [17:0]   img_reg_array_32_18_imag;
  reg        [17:0]   img_reg_array_32_19_real;
  reg        [17:0]   img_reg_array_32_19_imag;
  reg        [17:0]   img_reg_array_32_20_real;
  reg        [17:0]   img_reg_array_32_20_imag;
  reg        [17:0]   img_reg_array_32_21_real;
  reg        [17:0]   img_reg_array_32_21_imag;
  reg        [17:0]   img_reg_array_32_22_real;
  reg        [17:0]   img_reg_array_32_22_imag;
  reg        [17:0]   img_reg_array_32_23_real;
  reg        [17:0]   img_reg_array_32_23_imag;
  reg        [17:0]   img_reg_array_32_24_real;
  reg        [17:0]   img_reg_array_32_24_imag;
  reg        [17:0]   img_reg_array_32_25_real;
  reg        [17:0]   img_reg_array_32_25_imag;
  reg        [17:0]   img_reg_array_32_26_real;
  reg        [17:0]   img_reg_array_32_26_imag;
  reg        [17:0]   img_reg_array_32_27_real;
  reg        [17:0]   img_reg_array_32_27_imag;
  reg        [17:0]   img_reg_array_32_28_real;
  reg        [17:0]   img_reg_array_32_28_imag;
  reg        [17:0]   img_reg_array_32_29_real;
  reg        [17:0]   img_reg_array_32_29_imag;
  reg        [17:0]   img_reg_array_32_30_real;
  reg        [17:0]   img_reg_array_32_30_imag;
  reg        [17:0]   img_reg_array_32_31_real;
  reg        [17:0]   img_reg_array_32_31_imag;
  reg        [17:0]   img_reg_array_32_32_real;
  reg        [17:0]   img_reg_array_32_32_imag;
  reg        [17:0]   img_reg_array_32_33_real;
  reg        [17:0]   img_reg_array_32_33_imag;
  reg        [17:0]   img_reg_array_32_34_real;
  reg        [17:0]   img_reg_array_32_34_imag;
  reg        [17:0]   img_reg_array_32_35_real;
  reg        [17:0]   img_reg_array_32_35_imag;
  reg        [17:0]   img_reg_array_32_36_real;
  reg        [17:0]   img_reg_array_32_36_imag;
  reg        [17:0]   img_reg_array_32_37_real;
  reg        [17:0]   img_reg_array_32_37_imag;
  reg        [17:0]   img_reg_array_32_38_real;
  reg        [17:0]   img_reg_array_32_38_imag;
  reg        [17:0]   img_reg_array_32_39_real;
  reg        [17:0]   img_reg_array_32_39_imag;
  reg        [17:0]   img_reg_array_32_40_real;
  reg        [17:0]   img_reg_array_32_40_imag;
  reg        [17:0]   img_reg_array_32_41_real;
  reg        [17:0]   img_reg_array_32_41_imag;
  reg        [17:0]   img_reg_array_32_42_real;
  reg        [17:0]   img_reg_array_32_42_imag;
  reg        [17:0]   img_reg_array_32_43_real;
  reg        [17:0]   img_reg_array_32_43_imag;
  reg        [17:0]   img_reg_array_32_44_real;
  reg        [17:0]   img_reg_array_32_44_imag;
  reg        [17:0]   img_reg_array_32_45_real;
  reg        [17:0]   img_reg_array_32_45_imag;
  reg        [17:0]   img_reg_array_32_46_real;
  reg        [17:0]   img_reg_array_32_46_imag;
  reg        [17:0]   img_reg_array_32_47_real;
  reg        [17:0]   img_reg_array_32_47_imag;
  reg        [17:0]   img_reg_array_32_48_real;
  reg        [17:0]   img_reg_array_32_48_imag;
  reg        [17:0]   img_reg_array_32_49_real;
  reg        [17:0]   img_reg_array_32_49_imag;
  reg        [17:0]   img_reg_array_32_50_real;
  reg        [17:0]   img_reg_array_32_50_imag;
  reg        [17:0]   img_reg_array_32_51_real;
  reg        [17:0]   img_reg_array_32_51_imag;
  reg        [17:0]   img_reg_array_32_52_real;
  reg        [17:0]   img_reg_array_32_52_imag;
  reg        [17:0]   img_reg_array_32_53_real;
  reg        [17:0]   img_reg_array_32_53_imag;
  reg        [17:0]   img_reg_array_32_54_real;
  reg        [17:0]   img_reg_array_32_54_imag;
  reg        [17:0]   img_reg_array_32_55_real;
  reg        [17:0]   img_reg_array_32_55_imag;
  reg        [17:0]   img_reg_array_32_56_real;
  reg        [17:0]   img_reg_array_32_56_imag;
  reg        [17:0]   img_reg_array_32_57_real;
  reg        [17:0]   img_reg_array_32_57_imag;
  reg        [17:0]   img_reg_array_32_58_real;
  reg        [17:0]   img_reg_array_32_58_imag;
  reg        [17:0]   img_reg_array_32_59_real;
  reg        [17:0]   img_reg_array_32_59_imag;
  reg        [17:0]   img_reg_array_32_60_real;
  reg        [17:0]   img_reg_array_32_60_imag;
  reg        [17:0]   img_reg_array_32_61_real;
  reg        [17:0]   img_reg_array_32_61_imag;
  reg        [17:0]   img_reg_array_32_62_real;
  reg        [17:0]   img_reg_array_32_62_imag;
  reg        [17:0]   img_reg_array_32_63_real;
  reg        [17:0]   img_reg_array_32_63_imag;
  reg        [17:0]   img_reg_array_33_0_real;
  reg        [17:0]   img_reg_array_33_0_imag;
  reg        [17:0]   img_reg_array_33_1_real;
  reg        [17:0]   img_reg_array_33_1_imag;
  reg        [17:0]   img_reg_array_33_2_real;
  reg        [17:0]   img_reg_array_33_2_imag;
  reg        [17:0]   img_reg_array_33_3_real;
  reg        [17:0]   img_reg_array_33_3_imag;
  reg        [17:0]   img_reg_array_33_4_real;
  reg        [17:0]   img_reg_array_33_4_imag;
  reg        [17:0]   img_reg_array_33_5_real;
  reg        [17:0]   img_reg_array_33_5_imag;
  reg        [17:0]   img_reg_array_33_6_real;
  reg        [17:0]   img_reg_array_33_6_imag;
  reg        [17:0]   img_reg_array_33_7_real;
  reg        [17:0]   img_reg_array_33_7_imag;
  reg        [17:0]   img_reg_array_33_8_real;
  reg        [17:0]   img_reg_array_33_8_imag;
  reg        [17:0]   img_reg_array_33_9_real;
  reg        [17:0]   img_reg_array_33_9_imag;
  reg        [17:0]   img_reg_array_33_10_real;
  reg        [17:0]   img_reg_array_33_10_imag;
  reg        [17:0]   img_reg_array_33_11_real;
  reg        [17:0]   img_reg_array_33_11_imag;
  reg        [17:0]   img_reg_array_33_12_real;
  reg        [17:0]   img_reg_array_33_12_imag;
  reg        [17:0]   img_reg_array_33_13_real;
  reg        [17:0]   img_reg_array_33_13_imag;
  reg        [17:0]   img_reg_array_33_14_real;
  reg        [17:0]   img_reg_array_33_14_imag;
  reg        [17:0]   img_reg_array_33_15_real;
  reg        [17:0]   img_reg_array_33_15_imag;
  reg        [17:0]   img_reg_array_33_16_real;
  reg        [17:0]   img_reg_array_33_16_imag;
  reg        [17:0]   img_reg_array_33_17_real;
  reg        [17:0]   img_reg_array_33_17_imag;
  reg        [17:0]   img_reg_array_33_18_real;
  reg        [17:0]   img_reg_array_33_18_imag;
  reg        [17:0]   img_reg_array_33_19_real;
  reg        [17:0]   img_reg_array_33_19_imag;
  reg        [17:0]   img_reg_array_33_20_real;
  reg        [17:0]   img_reg_array_33_20_imag;
  reg        [17:0]   img_reg_array_33_21_real;
  reg        [17:0]   img_reg_array_33_21_imag;
  reg        [17:0]   img_reg_array_33_22_real;
  reg        [17:0]   img_reg_array_33_22_imag;
  reg        [17:0]   img_reg_array_33_23_real;
  reg        [17:0]   img_reg_array_33_23_imag;
  reg        [17:0]   img_reg_array_33_24_real;
  reg        [17:0]   img_reg_array_33_24_imag;
  reg        [17:0]   img_reg_array_33_25_real;
  reg        [17:0]   img_reg_array_33_25_imag;
  reg        [17:0]   img_reg_array_33_26_real;
  reg        [17:0]   img_reg_array_33_26_imag;
  reg        [17:0]   img_reg_array_33_27_real;
  reg        [17:0]   img_reg_array_33_27_imag;
  reg        [17:0]   img_reg_array_33_28_real;
  reg        [17:0]   img_reg_array_33_28_imag;
  reg        [17:0]   img_reg_array_33_29_real;
  reg        [17:0]   img_reg_array_33_29_imag;
  reg        [17:0]   img_reg_array_33_30_real;
  reg        [17:0]   img_reg_array_33_30_imag;
  reg        [17:0]   img_reg_array_33_31_real;
  reg        [17:0]   img_reg_array_33_31_imag;
  reg        [17:0]   img_reg_array_33_32_real;
  reg        [17:0]   img_reg_array_33_32_imag;
  reg        [17:0]   img_reg_array_33_33_real;
  reg        [17:0]   img_reg_array_33_33_imag;
  reg        [17:0]   img_reg_array_33_34_real;
  reg        [17:0]   img_reg_array_33_34_imag;
  reg        [17:0]   img_reg_array_33_35_real;
  reg        [17:0]   img_reg_array_33_35_imag;
  reg        [17:0]   img_reg_array_33_36_real;
  reg        [17:0]   img_reg_array_33_36_imag;
  reg        [17:0]   img_reg_array_33_37_real;
  reg        [17:0]   img_reg_array_33_37_imag;
  reg        [17:0]   img_reg_array_33_38_real;
  reg        [17:0]   img_reg_array_33_38_imag;
  reg        [17:0]   img_reg_array_33_39_real;
  reg        [17:0]   img_reg_array_33_39_imag;
  reg        [17:0]   img_reg_array_33_40_real;
  reg        [17:0]   img_reg_array_33_40_imag;
  reg        [17:0]   img_reg_array_33_41_real;
  reg        [17:0]   img_reg_array_33_41_imag;
  reg        [17:0]   img_reg_array_33_42_real;
  reg        [17:0]   img_reg_array_33_42_imag;
  reg        [17:0]   img_reg_array_33_43_real;
  reg        [17:0]   img_reg_array_33_43_imag;
  reg        [17:0]   img_reg_array_33_44_real;
  reg        [17:0]   img_reg_array_33_44_imag;
  reg        [17:0]   img_reg_array_33_45_real;
  reg        [17:0]   img_reg_array_33_45_imag;
  reg        [17:0]   img_reg_array_33_46_real;
  reg        [17:0]   img_reg_array_33_46_imag;
  reg        [17:0]   img_reg_array_33_47_real;
  reg        [17:0]   img_reg_array_33_47_imag;
  reg        [17:0]   img_reg_array_33_48_real;
  reg        [17:0]   img_reg_array_33_48_imag;
  reg        [17:0]   img_reg_array_33_49_real;
  reg        [17:0]   img_reg_array_33_49_imag;
  reg        [17:0]   img_reg_array_33_50_real;
  reg        [17:0]   img_reg_array_33_50_imag;
  reg        [17:0]   img_reg_array_33_51_real;
  reg        [17:0]   img_reg_array_33_51_imag;
  reg        [17:0]   img_reg_array_33_52_real;
  reg        [17:0]   img_reg_array_33_52_imag;
  reg        [17:0]   img_reg_array_33_53_real;
  reg        [17:0]   img_reg_array_33_53_imag;
  reg        [17:0]   img_reg_array_33_54_real;
  reg        [17:0]   img_reg_array_33_54_imag;
  reg        [17:0]   img_reg_array_33_55_real;
  reg        [17:0]   img_reg_array_33_55_imag;
  reg        [17:0]   img_reg_array_33_56_real;
  reg        [17:0]   img_reg_array_33_56_imag;
  reg        [17:0]   img_reg_array_33_57_real;
  reg        [17:0]   img_reg_array_33_57_imag;
  reg        [17:0]   img_reg_array_33_58_real;
  reg        [17:0]   img_reg_array_33_58_imag;
  reg        [17:0]   img_reg_array_33_59_real;
  reg        [17:0]   img_reg_array_33_59_imag;
  reg        [17:0]   img_reg_array_33_60_real;
  reg        [17:0]   img_reg_array_33_60_imag;
  reg        [17:0]   img_reg_array_33_61_real;
  reg        [17:0]   img_reg_array_33_61_imag;
  reg        [17:0]   img_reg_array_33_62_real;
  reg        [17:0]   img_reg_array_33_62_imag;
  reg        [17:0]   img_reg_array_33_63_real;
  reg        [17:0]   img_reg_array_33_63_imag;
  reg        [17:0]   img_reg_array_34_0_real;
  reg        [17:0]   img_reg_array_34_0_imag;
  reg        [17:0]   img_reg_array_34_1_real;
  reg        [17:0]   img_reg_array_34_1_imag;
  reg        [17:0]   img_reg_array_34_2_real;
  reg        [17:0]   img_reg_array_34_2_imag;
  reg        [17:0]   img_reg_array_34_3_real;
  reg        [17:0]   img_reg_array_34_3_imag;
  reg        [17:0]   img_reg_array_34_4_real;
  reg        [17:0]   img_reg_array_34_4_imag;
  reg        [17:0]   img_reg_array_34_5_real;
  reg        [17:0]   img_reg_array_34_5_imag;
  reg        [17:0]   img_reg_array_34_6_real;
  reg        [17:0]   img_reg_array_34_6_imag;
  reg        [17:0]   img_reg_array_34_7_real;
  reg        [17:0]   img_reg_array_34_7_imag;
  reg        [17:0]   img_reg_array_34_8_real;
  reg        [17:0]   img_reg_array_34_8_imag;
  reg        [17:0]   img_reg_array_34_9_real;
  reg        [17:0]   img_reg_array_34_9_imag;
  reg        [17:0]   img_reg_array_34_10_real;
  reg        [17:0]   img_reg_array_34_10_imag;
  reg        [17:0]   img_reg_array_34_11_real;
  reg        [17:0]   img_reg_array_34_11_imag;
  reg        [17:0]   img_reg_array_34_12_real;
  reg        [17:0]   img_reg_array_34_12_imag;
  reg        [17:0]   img_reg_array_34_13_real;
  reg        [17:0]   img_reg_array_34_13_imag;
  reg        [17:0]   img_reg_array_34_14_real;
  reg        [17:0]   img_reg_array_34_14_imag;
  reg        [17:0]   img_reg_array_34_15_real;
  reg        [17:0]   img_reg_array_34_15_imag;
  reg        [17:0]   img_reg_array_34_16_real;
  reg        [17:0]   img_reg_array_34_16_imag;
  reg        [17:0]   img_reg_array_34_17_real;
  reg        [17:0]   img_reg_array_34_17_imag;
  reg        [17:0]   img_reg_array_34_18_real;
  reg        [17:0]   img_reg_array_34_18_imag;
  reg        [17:0]   img_reg_array_34_19_real;
  reg        [17:0]   img_reg_array_34_19_imag;
  reg        [17:0]   img_reg_array_34_20_real;
  reg        [17:0]   img_reg_array_34_20_imag;
  reg        [17:0]   img_reg_array_34_21_real;
  reg        [17:0]   img_reg_array_34_21_imag;
  reg        [17:0]   img_reg_array_34_22_real;
  reg        [17:0]   img_reg_array_34_22_imag;
  reg        [17:0]   img_reg_array_34_23_real;
  reg        [17:0]   img_reg_array_34_23_imag;
  reg        [17:0]   img_reg_array_34_24_real;
  reg        [17:0]   img_reg_array_34_24_imag;
  reg        [17:0]   img_reg_array_34_25_real;
  reg        [17:0]   img_reg_array_34_25_imag;
  reg        [17:0]   img_reg_array_34_26_real;
  reg        [17:0]   img_reg_array_34_26_imag;
  reg        [17:0]   img_reg_array_34_27_real;
  reg        [17:0]   img_reg_array_34_27_imag;
  reg        [17:0]   img_reg_array_34_28_real;
  reg        [17:0]   img_reg_array_34_28_imag;
  reg        [17:0]   img_reg_array_34_29_real;
  reg        [17:0]   img_reg_array_34_29_imag;
  reg        [17:0]   img_reg_array_34_30_real;
  reg        [17:0]   img_reg_array_34_30_imag;
  reg        [17:0]   img_reg_array_34_31_real;
  reg        [17:0]   img_reg_array_34_31_imag;
  reg        [17:0]   img_reg_array_34_32_real;
  reg        [17:0]   img_reg_array_34_32_imag;
  reg        [17:0]   img_reg_array_34_33_real;
  reg        [17:0]   img_reg_array_34_33_imag;
  reg        [17:0]   img_reg_array_34_34_real;
  reg        [17:0]   img_reg_array_34_34_imag;
  reg        [17:0]   img_reg_array_34_35_real;
  reg        [17:0]   img_reg_array_34_35_imag;
  reg        [17:0]   img_reg_array_34_36_real;
  reg        [17:0]   img_reg_array_34_36_imag;
  reg        [17:0]   img_reg_array_34_37_real;
  reg        [17:0]   img_reg_array_34_37_imag;
  reg        [17:0]   img_reg_array_34_38_real;
  reg        [17:0]   img_reg_array_34_38_imag;
  reg        [17:0]   img_reg_array_34_39_real;
  reg        [17:0]   img_reg_array_34_39_imag;
  reg        [17:0]   img_reg_array_34_40_real;
  reg        [17:0]   img_reg_array_34_40_imag;
  reg        [17:0]   img_reg_array_34_41_real;
  reg        [17:0]   img_reg_array_34_41_imag;
  reg        [17:0]   img_reg_array_34_42_real;
  reg        [17:0]   img_reg_array_34_42_imag;
  reg        [17:0]   img_reg_array_34_43_real;
  reg        [17:0]   img_reg_array_34_43_imag;
  reg        [17:0]   img_reg_array_34_44_real;
  reg        [17:0]   img_reg_array_34_44_imag;
  reg        [17:0]   img_reg_array_34_45_real;
  reg        [17:0]   img_reg_array_34_45_imag;
  reg        [17:0]   img_reg_array_34_46_real;
  reg        [17:0]   img_reg_array_34_46_imag;
  reg        [17:0]   img_reg_array_34_47_real;
  reg        [17:0]   img_reg_array_34_47_imag;
  reg        [17:0]   img_reg_array_34_48_real;
  reg        [17:0]   img_reg_array_34_48_imag;
  reg        [17:0]   img_reg_array_34_49_real;
  reg        [17:0]   img_reg_array_34_49_imag;
  reg        [17:0]   img_reg_array_34_50_real;
  reg        [17:0]   img_reg_array_34_50_imag;
  reg        [17:0]   img_reg_array_34_51_real;
  reg        [17:0]   img_reg_array_34_51_imag;
  reg        [17:0]   img_reg_array_34_52_real;
  reg        [17:0]   img_reg_array_34_52_imag;
  reg        [17:0]   img_reg_array_34_53_real;
  reg        [17:0]   img_reg_array_34_53_imag;
  reg        [17:0]   img_reg_array_34_54_real;
  reg        [17:0]   img_reg_array_34_54_imag;
  reg        [17:0]   img_reg_array_34_55_real;
  reg        [17:0]   img_reg_array_34_55_imag;
  reg        [17:0]   img_reg_array_34_56_real;
  reg        [17:0]   img_reg_array_34_56_imag;
  reg        [17:0]   img_reg_array_34_57_real;
  reg        [17:0]   img_reg_array_34_57_imag;
  reg        [17:0]   img_reg_array_34_58_real;
  reg        [17:0]   img_reg_array_34_58_imag;
  reg        [17:0]   img_reg_array_34_59_real;
  reg        [17:0]   img_reg_array_34_59_imag;
  reg        [17:0]   img_reg_array_34_60_real;
  reg        [17:0]   img_reg_array_34_60_imag;
  reg        [17:0]   img_reg_array_34_61_real;
  reg        [17:0]   img_reg_array_34_61_imag;
  reg        [17:0]   img_reg_array_34_62_real;
  reg        [17:0]   img_reg_array_34_62_imag;
  reg        [17:0]   img_reg_array_34_63_real;
  reg        [17:0]   img_reg_array_34_63_imag;
  reg        [17:0]   img_reg_array_35_0_real;
  reg        [17:0]   img_reg_array_35_0_imag;
  reg        [17:0]   img_reg_array_35_1_real;
  reg        [17:0]   img_reg_array_35_1_imag;
  reg        [17:0]   img_reg_array_35_2_real;
  reg        [17:0]   img_reg_array_35_2_imag;
  reg        [17:0]   img_reg_array_35_3_real;
  reg        [17:0]   img_reg_array_35_3_imag;
  reg        [17:0]   img_reg_array_35_4_real;
  reg        [17:0]   img_reg_array_35_4_imag;
  reg        [17:0]   img_reg_array_35_5_real;
  reg        [17:0]   img_reg_array_35_5_imag;
  reg        [17:0]   img_reg_array_35_6_real;
  reg        [17:0]   img_reg_array_35_6_imag;
  reg        [17:0]   img_reg_array_35_7_real;
  reg        [17:0]   img_reg_array_35_7_imag;
  reg        [17:0]   img_reg_array_35_8_real;
  reg        [17:0]   img_reg_array_35_8_imag;
  reg        [17:0]   img_reg_array_35_9_real;
  reg        [17:0]   img_reg_array_35_9_imag;
  reg        [17:0]   img_reg_array_35_10_real;
  reg        [17:0]   img_reg_array_35_10_imag;
  reg        [17:0]   img_reg_array_35_11_real;
  reg        [17:0]   img_reg_array_35_11_imag;
  reg        [17:0]   img_reg_array_35_12_real;
  reg        [17:0]   img_reg_array_35_12_imag;
  reg        [17:0]   img_reg_array_35_13_real;
  reg        [17:0]   img_reg_array_35_13_imag;
  reg        [17:0]   img_reg_array_35_14_real;
  reg        [17:0]   img_reg_array_35_14_imag;
  reg        [17:0]   img_reg_array_35_15_real;
  reg        [17:0]   img_reg_array_35_15_imag;
  reg        [17:0]   img_reg_array_35_16_real;
  reg        [17:0]   img_reg_array_35_16_imag;
  reg        [17:0]   img_reg_array_35_17_real;
  reg        [17:0]   img_reg_array_35_17_imag;
  reg        [17:0]   img_reg_array_35_18_real;
  reg        [17:0]   img_reg_array_35_18_imag;
  reg        [17:0]   img_reg_array_35_19_real;
  reg        [17:0]   img_reg_array_35_19_imag;
  reg        [17:0]   img_reg_array_35_20_real;
  reg        [17:0]   img_reg_array_35_20_imag;
  reg        [17:0]   img_reg_array_35_21_real;
  reg        [17:0]   img_reg_array_35_21_imag;
  reg        [17:0]   img_reg_array_35_22_real;
  reg        [17:0]   img_reg_array_35_22_imag;
  reg        [17:0]   img_reg_array_35_23_real;
  reg        [17:0]   img_reg_array_35_23_imag;
  reg        [17:0]   img_reg_array_35_24_real;
  reg        [17:0]   img_reg_array_35_24_imag;
  reg        [17:0]   img_reg_array_35_25_real;
  reg        [17:0]   img_reg_array_35_25_imag;
  reg        [17:0]   img_reg_array_35_26_real;
  reg        [17:0]   img_reg_array_35_26_imag;
  reg        [17:0]   img_reg_array_35_27_real;
  reg        [17:0]   img_reg_array_35_27_imag;
  reg        [17:0]   img_reg_array_35_28_real;
  reg        [17:0]   img_reg_array_35_28_imag;
  reg        [17:0]   img_reg_array_35_29_real;
  reg        [17:0]   img_reg_array_35_29_imag;
  reg        [17:0]   img_reg_array_35_30_real;
  reg        [17:0]   img_reg_array_35_30_imag;
  reg        [17:0]   img_reg_array_35_31_real;
  reg        [17:0]   img_reg_array_35_31_imag;
  reg        [17:0]   img_reg_array_35_32_real;
  reg        [17:0]   img_reg_array_35_32_imag;
  reg        [17:0]   img_reg_array_35_33_real;
  reg        [17:0]   img_reg_array_35_33_imag;
  reg        [17:0]   img_reg_array_35_34_real;
  reg        [17:0]   img_reg_array_35_34_imag;
  reg        [17:0]   img_reg_array_35_35_real;
  reg        [17:0]   img_reg_array_35_35_imag;
  reg        [17:0]   img_reg_array_35_36_real;
  reg        [17:0]   img_reg_array_35_36_imag;
  reg        [17:0]   img_reg_array_35_37_real;
  reg        [17:0]   img_reg_array_35_37_imag;
  reg        [17:0]   img_reg_array_35_38_real;
  reg        [17:0]   img_reg_array_35_38_imag;
  reg        [17:0]   img_reg_array_35_39_real;
  reg        [17:0]   img_reg_array_35_39_imag;
  reg        [17:0]   img_reg_array_35_40_real;
  reg        [17:0]   img_reg_array_35_40_imag;
  reg        [17:0]   img_reg_array_35_41_real;
  reg        [17:0]   img_reg_array_35_41_imag;
  reg        [17:0]   img_reg_array_35_42_real;
  reg        [17:0]   img_reg_array_35_42_imag;
  reg        [17:0]   img_reg_array_35_43_real;
  reg        [17:0]   img_reg_array_35_43_imag;
  reg        [17:0]   img_reg_array_35_44_real;
  reg        [17:0]   img_reg_array_35_44_imag;
  reg        [17:0]   img_reg_array_35_45_real;
  reg        [17:0]   img_reg_array_35_45_imag;
  reg        [17:0]   img_reg_array_35_46_real;
  reg        [17:0]   img_reg_array_35_46_imag;
  reg        [17:0]   img_reg_array_35_47_real;
  reg        [17:0]   img_reg_array_35_47_imag;
  reg        [17:0]   img_reg_array_35_48_real;
  reg        [17:0]   img_reg_array_35_48_imag;
  reg        [17:0]   img_reg_array_35_49_real;
  reg        [17:0]   img_reg_array_35_49_imag;
  reg        [17:0]   img_reg_array_35_50_real;
  reg        [17:0]   img_reg_array_35_50_imag;
  reg        [17:0]   img_reg_array_35_51_real;
  reg        [17:0]   img_reg_array_35_51_imag;
  reg        [17:0]   img_reg_array_35_52_real;
  reg        [17:0]   img_reg_array_35_52_imag;
  reg        [17:0]   img_reg_array_35_53_real;
  reg        [17:0]   img_reg_array_35_53_imag;
  reg        [17:0]   img_reg_array_35_54_real;
  reg        [17:0]   img_reg_array_35_54_imag;
  reg        [17:0]   img_reg_array_35_55_real;
  reg        [17:0]   img_reg_array_35_55_imag;
  reg        [17:0]   img_reg_array_35_56_real;
  reg        [17:0]   img_reg_array_35_56_imag;
  reg        [17:0]   img_reg_array_35_57_real;
  reg        [17:0]   img_reg_array_35_57_imag;
  reg        [17:0]   img_reg_array_35_58_real;
  reg        [17:0]   img_reg_array_35_58_imag;
  reg        [17:0]   img_reg_array_35_59_real;
  reg        [17:0]   img_reg_array_35_59_imag;
  reg        [17:0]   img_reg_array_35_60_real;
  reg        [17:0]   img_reg_array_35_60_imag;
  reg        [17:0]   img_reg_array_35_61_real;
  reg        [17:0]   img_reg_array_35_61_imag;
  reg        [17:0]   img_reg_array_35_62_real;
  reg        [17:0]   img_reg_array_35_62_imag;
  reg        [17:0]   img_reg_array_35_63_real;
  reg        [17:0]   img_reg_array_35_63_imag;
  reg        [17:0]   img_reg_array_36_0_real;
  reg        [17:0]   img_reg_array_36_0_imag;
  reg        [17:0]   img_reg_array_36_1_real;
  reg        [17:0]   img_reg_array_36_1_imag;
  reg        [17:0]   img_reg_array_36_2_real;
  reg        [17:0]   img_reg_array_36_2_imag;
  reg        [17:0]   img_reg_array_36_3_real;
  reg        [17:0]   img_reg_array_36_3_imag;
  reg        [17:0]   img_reg_array_36_4_real;
  reg        [17:0]   img_reg_array_36_4_imag;
  reg        [17:0]   img_reg_array_36_5_real;
  reg        [17:0]   img_reg_array_36_5_imag;
  reg        [17:0]   img_reg_array_36_6_real;
  reg        [17:0]   img_reg_array_36_6_imag;
  reg        [17:0]   img_reg_array_36_7_real;
  reg        [17:0]   img_reg_array_36_7_imag;
  reg        [17:0]   img_reg_array_36_8_real;
  reg        [17:0]   img_reg_array_36_8_imag;
  reg        [17:0]   img_reg_array_36_9_real;
  reg        [17:0]   img_reg_array_36_9_imag;
  reg        [17:0]   img_reg_array_36_10_real;
  reg        [17:0]   img_reg_array_36_10_imag;
  reg        [17:0]   img_reg_array_36_11_real;
  reg        [17:0]   img_reg_array_36_11_imag;
  reg        [17:0]   img_reg_array_36_12_real;
  reg        [17:0]   img_reg_array_36_12_imag;
  reg        [17:0]   img_reg_array_36_13_real;
  reg        [17:0]   img_reg_array_36_13_imag;
  reg        [17:0]   img_reg_array_36_14_real;
  reg        [17:0]   img_reg_array_36_14_imag;
  reg        [17:0]   img_reg_array_36_15_real;
  reg        [17:0]   img_reg_array_36_15_imag;
  reg        [17:0]   img_reg_array_36_16_real;
  reg        [17:0]   img_reg_array_36_16_imag;
  reg        [17:0]   img_reg_array_36_17_real;
  reg        [17:0]   img_reg_array_36_17_imag;
  reg        [17:0]   img_reg_array_36_18_real;
  reg        [17:0]   img_reg_array_36_18_imag;
  reg        [17:0]   img_reg_array_36_19_real;
  reg        [17:0]   img_reg_array_36_19_imag;
  reg        [17:0]   img_reg_array_36_20_real;
  reg        [17:0]   img_reg_array_36_20_imag;
  reg        [17:0]   img_reg_array_36_21_real;
  reg        [17:0]   img_reg_array_36_21_imag;
  reg        [17:0]   img_reg_array_36_22_real;
  reg        [17:0]   img_reg_array_36_22_imag;
  reg        [17:0]   img_reg_array_36_23_real;
  reg        [17:0]   img_reg_array_36_23_imag;
  reg        [17:0]   img_reg_array_36_24_real;
  reg        [17:0]   img_reg_array_36_24_imag;
  reg        [17:0]   img_reg_array_36_25_real;
  reg        [17:0]   img_reg_array_36_25_imag;
  reg        [17:0]   img_reg_array_36_26_real;
  reg        [17:0]   img_reg_array_36_26_imag;
  reg        [17:0]   img_reg_array_36_27_real;
  reg        [17:0]   img_reg_array_36_27_imag;
  reg        [17:0]   img_reg_array_36_28_real;
  reg        [17:0]   img_reg_array_36_28_imag;
  reg        [17:0]   img_reg_array_36_29_real;
  reg        [17:0]   img_reg_array_36_29_imag;
  reg        [17:0]   img_reg_array_36_30_real;
  reg        [17:0]   img_reg_array_36_30_imag;
  reg        [17:0]   img_reg_array_36_31_real;
  reg        [17:0]   img_reg_array_36_31_imag;
  reg        [17:0]   img_reg_array_36_32_real;
  reg        [17:0]   img_reg_array_36_32_imag;
  reg        [17:0]   img_reg_array_36_33_real;
  reg        [17:0]   img_reg_array_36_33_imag;
  reg        [17:0]   img_reg_array_36_34_real;
  reg        [17:0]   img_reg_array_36_34_imag;
  reg        [17:0]   img_reg_array_36_35_real;
  reg        [17:0]   img_reg_array_36_35_imag;
  reg        [17:0]   img_reg_array_36_36_real;
  reg        [17:0]   img_reg_array_36_36_imag;
  reg        [17:0]   img_reg_array_36_37_real;
  reg        [17:0]   img_reg_array_36_37_imag;
  reg        [17:0]   img_reg_array_36_38_real;
  reg        [17:0]   img_reg_array_36_38_imag;
  reg        [17:0]   img_reg_array_36_39_real;
  reg        [17:0]   img_reg_array_36_39_imag;
  reg        [17:0]   img_reg_array_36_40_real;
  reg        [17:0]   img_reg_array_36_40_imag;
  reg        [17:0]   img_reg_array_36_41_real;
  reg        [17:0]   img_reg_array_36_41_imag;
  reg        [17:0]   img_reg_array_36_42_real;
  reg        [17:0]   img_reg_array_36_42_imag;
  reg        [17:0]   img_reg_array_36_43_real;
  reg        [17:0]   img_reg_array_36_43_imag;
  reg        [17:0]   img_reg_array_36_44_real;
  reg        [17:0]   img_reg_array_36_44_imag;
  reg        [17:0]   img_reg_array_36_45_real;
  reg        [17:0]   img_reg_array_36_45_imag;
  reg        [17:0]   img_reg_array_36_46_real;
  reg        [17:0]   img_reg_array_36_46_imag;
  reg        [17:0]   img_reg_array_36_47_real;
  reg        [17:0]   img_reg_array_36_47_imag;
  reg        [17:0]   img_reg_array_36_48_real;
  reg        [17:0]   img_reg_array_36_48_imag;
  reg        [17:0]   img_reg_array_36_49_real;
  reg        [17:0]   img_reg_array_36_49_imag;
  reg        [17:0]   img_reg_array_36_50_real;
  reg        [17:0]   img_reg_array_36_50_imag;
  reg        [17:0]   img_reg_array_36_51_real;
  reg        [17:0]   img_reg_array_36_51_imag;
  reg        [17:0]   img_reg_array_36_52_real;
  reg        [17:0]   img_reg_array_36_52_imag;
  reg        [17:0]   img_reg_array_36_53_real;
  reg        [17:0]   img_reg_array_36_53_imag;
  reg        [17:0]   img_reg_array_36_54_real;
  reg        [17:0]   img_reg_array_36_54_imag;
  reg        [17:0]   img_reg_array_36_55_real;
  reg        [17:0]   img_reg_array_36_55_imag;
  reg        [17:0]   img_reg_array_36_56_real;
  reg        [17:0]   img_reg_array_36_56_imag;
  reg        [17:0]   img_reg_array_36_57_real;
  reg        [17:0]   img_reg_array_36_57_imag;
  reg        [17:0]   img_reg_array_36_58_real;
  reg        [17:0]   img_reg_array_36_58_imag;
  reg        [17:0]   img_reg_array_36_59_real;
  reg        [17:0]   img_reg_array_36_59_imag;
  reg        [17:0]   img_reg_array_36_60_real;
  reg        [17:0]   img_reg_array_36_60_imag;
  reg        [17:0]   img_reg_array_36_61_real;
  reg        [17:0]   img_reg_array_36_61_imag;
  reg        [17:0]   img_reg_array_36_62_real;
  reg        [17:0]   img_reg_array_36_62_imag;
  reg        [17:0]   img_reg_array_36_63_real;
  reg        [17:0]   img_reg_array_36_63_imag;
  reg        [17:0]   img_reg_array_37_0_real;
  reg        [17:0]   img_reg_array_37_0_imag;
  reg        [17:0]   img_reg_array_37_1_real;
  reg        [17:0]   img_reg_array_37_1_imag;
  reg        [17:0]   img_reg_array_37_2_real;
  reg        [17:0]   img_reg_array_37_2_imag;
  reg        [17:0]   img_reg_array_37_3_real;
  reg        [17:0]   img_reg_array_37_3_imag;
  reg        [17:0]   img_reg_array_37_4_real;
  reg        [17:0]   img_reg_array_37_4_imag;
  reg        [17:0]   img_reg_array_37_5_real;
  reg        [17:0]   img_reg_array_37_5_imag;
  reg        [17:0]   img_reg_array_37_6_real;
  reg        [17:0]   img_reg_array_37_6_imag;
  reg        [17:0]   img_reg_array_37_7_real;
  reg        [17:0]   img_reg_array_37_7_imag;
  reg        [17:0]   img_reg_array_37_8_real;
  reg        [17:0]   img_reg_array_37_8_imag;
  reg        [17:0]   img_reg_array_37_9_real;
  reg        [17:0]   img_reg_array_37_9_imag;
  reg        [17:0]   img_reg_array_37_10_real;
  reg        [17:0]   img_reg_array_37_10_imag;
  reg        [17:0]   img_reg_array_37_11_real;
  reg        [17:0]   img_reg_array_37_11_imag;
  reg        [17:0]   img_reg_array_37_12_real;
  reg        [17:0]   img_reg_array_37_12_imag;
  reg        [17:0]   img_reg_array_37_13_real;
  reg        [17:0]   img_reg_array_37_13_imag;
  reg        [17:0]   img_reg_array_37_14_real;
  reg        [17:0]   img_reg_array_37_14_imag;
  reg        [17:0]   img_reg_array_37_15_real;
  reg        [17:0]   img_reg_array_37_15_imag;
  reg        [17:0]   img_reg_array_37_16_real;
  reg        [17:0]   img_reg_array_37_16_imag;
  reg        [17:0]   img_reg_array_37_17_real;
  reg        [17:0]   img_reg_array_37_17_imag;
  reg        [17:0]   img_reg_array_37_18_real;
  reg        [17:0]   img_reg_array_37_18_imag;
  reg        [17:0]   img_reg_array_37_19_real;
  reg        [17:0]   img_reg_array_37_19_imag;
  reg        [17:0]   img_reg_array_37_20_real;
  reg        [17:0]   img_reg_array_37_20_imag;
  reg        [17:0]   img_reg_array_37_21_real;
  reg        [17:0]   img_reg_array_37_21_imag;
  reg        [17:0]   img_reg_array_37_22_real;
  reg        [17:0]   img_reg_array_37_22_imag;
  reg        [17:0]   img_reg_array_37_23_real;
  reg        [17:0]   img_reg_array_37_23_imag;
  reg        [17:0]   img_reg_array_37_24_real;
  reg        [17:0]   img_reg_array_37_24_imag;
  reg        [17:0]   img_reg_array_37_25_real;
  reg        [17:0]   img_reg_array_37_25_imag;
  reg        [17:0]   img_reg_array_37_26_real;
  reg        [17:0]   img_reg_array_37_26_imag;
  reg        [17:0]   img_reg_array_37_27_real;
  reg        [17:0]   img_reg_array_37_27_imag;
  reg        [17:0]   img_reg_array_37_28_real;
  reg        [17:0]   img_reg_array_37_28_imag;
  reg        [17:0]   img_reg_array_37_29_real;
  reg        [17:0]   img_reg_array_37_29_imag;
  reg        [17:0]   img_reg_array_37_30_real;
  reg        [17:0]   img_reg_array_37_30_imag;
  reg        [17:0]   img_reg_array_37_31_real;
  reg        [17:0]   img_reg_array_37_31_imag;
  reg        [17:0]   img_reg_array_37_32_real;
  reg        [17:0]   img_reg_array_37_32_imag;
  reg        [17:0]   img_reg_array_37_33_real;
  reg        [17:0]   img_reg_array_37_33_imag;
  reg        [17:0]   img_reg_array_37_34_real;
  reg        [17:0]   img_reg_array_37_34_imag;
  reg        [17:0]   img_reg_array_37_35_real;
  reg        [17:0]   img_reg_array_37_35_imag;
  reg        [17:0]   img_reg_array_37_36_real;
  reg        [17:0]   img_reg_array_37_36_imag;
  reg        [17:0]   img_reg_array_37_37_real;
  reg        [17:0]   img_reg_array_37_37_imag;
  reg        [17:0]   img_reg_array_37_38_real;
  reg        [17:0]   img_reg_array_37_38_imag;
  reg        [17:0]   img_reg_array_37_39_real;
  reg        [17:0]   img_reg_array_37_39_imag;
  reg        [17:0]   img_reg_array_37_40_real;
  reg        [17:0]   img_reg_array_37_40_imag;
  reg        [17:0]   img_reg_array_37_41_real;
  reg        [17:0]   img_reg_array_37_41_imag;
  reg        [17:0]   img_reg_array_37_42_real;
  reg        [17:0]   img_reg_array_37_42_imag;
  reg        [17:0]   img_reg_array_37_43_real;
  reg        [17:0]   img_reg_array_37_43_imag;
  reg        [17:0]   img_reg_array_37_44_real;
  reg        [17:0]   img_reg_array_37_44_imag;
  reg        [17:0]   img_reg_array_37_45_real;
  reg        [17:0]   img_reg_array_37_45_imag;
  reg        [17:0]   img_reg_array_37_46_real;
  reg        [17:0]   img_reg_array_37_46_imag;
  reg        [17:0]   img_reg_array_37_47_real;
  reg        [17:0]   img_reg_array_37_47_imag;
  reg        [17:0]   img_reg_array_37_48_real;
  reg        [17:0]   img_reg_array_37_48_imag;
  reg        [17:0]   img_reg_array_37_49_real;
  reg        [17:0]   img_reg_array_37_49_imag;
  reg        [17:0]   img_reg_array_37_50_real;
  reg        [17:0]   img_reg_array_37_50_imag;
  reg        [17:0]   img_reg_array_37_51_real;
  reg        [17:0]   img_reg_array_37_51_imag;
  reg        [17:0]   img_reg_array_37_52_real;
  reg        [17:0]   img_reg_array_37_52_imag;
  reg        [17:0]   img_reg_array_37_53_real;
  reg        [17:0]   img_reg_array_37_53_imag;
  reg        [17:0]   img_reg_array_37_54_real;
  reg        [17:0]   img_reg_array_37_54_imag;
  reg        [17:0]   img_reg_array_37_55_real;
  reg        [17:0]   img_reg_array_37_55_imag;
  reg        [17:0]   img_reg_array_37_56_real;
  reg        [17:0]   img_reg_array_37_56_imag;
  reg        [17:0]   img_reg_array_37_57_real;
  reg        [17:0]   img_reg_array_37_57_imag;
  reg        [17:0]   img_reg_array_37_58_real;
  reg        [17:0]   img_reg_array_37_58_imag;
  reg        [17:0]   img_reg_array_37_59_real;
  reg        [17:0]   img_reg_array_37_59_imag;
  reg        [17:0]   img_reg_array_37_60_real;
  reg        [17:0]   img_reg_array_37_60_imag;
  reg        [17:0]   img_reg_array_37_61_real;
  reg        [17:0]   img_reg_array_37_61_imag;
  reg        [17:0]   img_reg_array_37_62_real;
  reg        [17:0]   img_reg_array_37_62_imag;
  reg        [17:0]   img_reg_array_37_63_real;
  reg        [17:0]   img_reg_array_37_63_imag;
  reg        [17:0]   img_reg_array_38_0_real;
  reg        [17:0]   img_reg_array_38_0_imag;
  reg        [17:0]   img_reg_array_38_1_real;
  reg        [17:0]   img_reg_array_38_1_imag;
  reg        [17:0]   img_reg_array_38_2_real;
  reg        [17:0]   img_reg_array_38_2_imag;
  reg        [17:0]   img_reg_array_38_3_real;
  reg        [17:0]   img_reg_array_38_3_imag;
  reg        [17:0]   img_reg_array_38_4_real;
  reg        [17:0]   img_reg_array_38_4_imag;
  reg        [17:0]   img_reg_array_38_5_real;
  reg        [17:0]   img_reg_array_38_5_imag;
  reg        [17:0]   img_reg_array_38_6_real;
  reg        [17:0]   img_reg_array_38_6_imag;
  reg        [17:0]   img_reg_array_38_7_real;
  reg        [17:0]   img_reg_array_38_7_imag;
  reg        [17:0]   img_reg_array_38_8_real;
  reg        [17:0]   img_reg_array_38_8_imag;
  reg        [17:0]   img_reg_array_38_9_real;
  reg        [17:0]   img_reg_array_38_9_imag;
  reg        [17:0]   img_reg_array_38_10_real;
  reg        [17:0]   img_reg_array_38_10_imag;
  reg        [17:0]   img_reg_array_38_11_real;
  reg        [17:0]   img_reg_array_38_11_imag;
  reg        [17:0]   img_reg_array_38_12_real;
  reg        [17:0]   img_reg_array_38_12_imag;
  reg        [17:0]   img_reg_array_38_13_real;
  reg        [17:0]   img_reg_array_38_13_imag;
  reg        [17:0]   img_reg_array_38_14_real;
  reg        [17:0]   img_reg_array_38_14_imag;
  reg        [17:0]   img_reg_array_38_15_real;
  reg        [17:0]   img_reg_array_38_15_imag;
  reg        [17:0]   img_reg_array_38_16_real;
  reg        [17:0]   img_reg_array_38_16_imag;
  reg        [17:0]   img_reg_array_38_17_real;
  reg        [17:0]   img_reg_array_38_17_imag;
  reg        [17:0]   img_reg_array_38_18_real;
  reg        [17:0]   img_reg_array_38_18_imag;
  reg        [17:0]   img_reg_array_38_19_real;
  reg        [17:0]   img_reg_array_38_19_imag;
  reg        [17:0]   img_reg_array_38_20_real;
  reg        [17:0]   img_reg_array_38_20_imag;
  reg        [17:0]   img_reg_array_38_21_real;
  reg        [17:0]   img_reg_array_38_21_imag;
  reg        [17:0]   img_reg_array_38_22_real;
  reg        [17:0]   img_reg_array_38_22_imag;
  reg        [17:0]   img_reg_array_38_23_real;
  reg        [17:0]   img_reg_array_38_23_imag;
  reg        [17:0]   img_reg_array_38_24_real;
  reg        [17:0]   img_reg_array_38_24_imag;
  reg        [17:0]   img_reg_array_38_25_real;
  reg        [17:0]   img_reg_array_38_25_imag;
  reg        [17:0]   img_reg_array_38_26_real;
  reg        [17:0]   img_reg_array_38_26_imag;
  reg        [17:0]   img_reg_array_38_27_real;
  reg        [17:0]   img_reg_array_38_27_imag;
  reg        [17:0]   img_reg_array_38_28_real;
  reg        [17:0]   img_reg_array_38_28_imag;
  reg        [17:0]   img_reg_array_38_29_real;
  reg        [17:0]   img_reg_array_38_29_imag;
  reg        [17:0]   img_reg_array_38_30_real;
  reg        [17:0]   img_reg_array_38_30_imag;
  reg        [17:0]   img_reg_array_38_31_real;
  reg        [17:0]   img_reg_array_38_31_imag;
  reg        [17:0]   img_reg_array_38_32_real;
  reg        [17:0]   img_reg_array_38_32_imag;
  reg        [17:0]   img_reg_array_38_33_real;
  reg        [17:0]   img_reg_array_38_33_imag;
  reg        [17:0]   img_reg_array_38_34_real;
  reg        [17:0]   img_reg_array_38_34_imag;
  reg        [17:0]   img_reg_array_38_35_real;
  reg        [17:0]   img_reg_array_38_35_imag;
  reg        [17:0]   img_reg_array_38_36_real;
  reg        [17:0]   img_reg_array_38_36_imag;
  reg        [17:0]   img_reg_array_38_37_real;
  reg        [17:0]   img_reg_array_38_37_imag;
  reg        [17:0]   img_reg_array_38_38_real;
  reg        [17:0]   img_reg_array_38_38_imag;
  reg        [17:0]   img_reg_array_38_39_real;
  reg        [17:0]   img_reg_array_38_39_imag;
  reg        [17:0]   img_reg_array_38_40_real;
  reg        [17:0]   img_reg_array_38_40_imag;
  reg        [17:0]   img_reg_array_38_41_real;
  reg        [17:0]   img_reg_array_38_41_imag;
  reg        [17:0]   img_reg_array_38_42_real;
  reg        [17:0]   img_reg_array_38_42_imag;
  reg        [17:0]   img_reg_array_38_43_real;
  reg        [17:0]   img_reg_array_38_43_imag;
  reg        [17:0]   img_reg_array_38_44_real;
  reg        [17:0]   img_reg_array_38_44_imag;
  reg        [17:0]   img_reg_array_38_45_real;
  reg        [17:0]   img_reg_array_38_45_imag;
  reg        [17:0]   img_reg_array_38_46_real;
  reg        [17:0]   img_reg_array_38_46_imag;
  reg        [17:0]   img_reg_array_38_47_real;
  reg        [17:0]   img_reg_array_38_47_imag;
  reg        [17:0]   img_reg_array_38_48_real;
  reg        [17:0]   img_reg_array_38_48_imag;
  reg        [17:0]   img_reg_array_38_49_real;
  reg        [17:0]   img_reg_array_38_49_imag;
  reg        [17:0]   img_reg_array_38_50_real;
  reg        [17:0]   img_reg_array_38_50_imag;
  reg        [17:0]   img_reg_array_38_51_real;
  reg        [17:0]   img_reg_array_38_51_imag;
  reg        [17:0]   img_reg_array_38_52_real;
  reg        [17:0]   img_reg_array_38_52_imag;
  reg        [17:0]   img_reg_array_38_53_real;
  reg        [17:0]   img_reg_array_38_53_imag;
  reg        [17:0]   img_reg_array_38_54_real;
  reg        [17:0]   img_reg_array_38_54_imag;
  reg        [17:0]   img_reg_array_38_55_real;
  reg        [17:0]   img_reg_array_38_55_imag;
  reg        [17:0]   img_reg_array_38_56_real;
  reg        [17:0]   img_reg_array_38_56_imag;
  reg        [17:0]   img_reg_array_38_57_real;
  reg        [17:0]   img_reg_array_38_57_imag;
  reg        [17:0]   img_reg_array_38_58_real;
  reg        [17:0]   img_reg_array_38_58_imag;
  reg        [17:0]   img_reg_array_38_59_real;
  reg        [17:0]   img_reg_array_38_59_imag;
  reg        [17:0]   img_reg_array_38_60_real;
  reg        [17:0]   img_reg_array_38_60_imag;
  reg        [17:0]   img_reg_array_38_61_real;
  reg        [17:0]   img_reg_array_38_61_imag;
  reg        [17:0]   img_reg_array_38_62_real;
  reg        [17:0]   img_reg_array_38_62_imag;
  reg        [17:0]   img_reg_array_38_63_real;
  reg        [17:0]   img_reg_array_38_63_imag;
  reg        [17:0]   img_reg_array_39_0_real;
  reg        [17:0]   img_reg_array_39_0_imag;
  reg        [17:0]   img_reg_array_39_1_real;
  reg        [17:0]   img_reg_array_39_1_imag;
  reg        [17:0]   img_reg_array_39_2_real;
  reg        [17:0]   img_reg_array_39_2_imag;
  reg        [17:0]   img_reg_array_39_3_real;
  reg        [17:0]   img_reg_array_39_3_imag;
  reg        [17:0]   img_reg_array_39_4_real;
  reg        [17:0]   img_reg_array_39_4_imag;
  reg        [17:0]   img_reg_array_39_5_real;
  reg        [17:0]   img_reg_array_39_5_imag;
  reg        [17:0]   img_reg_array_39_6_real;
  reg        [17:0]   img_reg_array_39_6_imag;
  reg        [17:0]   img_reg_array_39_7_real;
  reg        [17:0]   img_reg_array_39_7_imag;
  reg        [17:0]   img_reg_array_39_8_real;
  reg        [17:0]   img_reg_array_39_8_imag;
  reg        [17:0]   img_reg_array_39_9_real;
  reg        [17:0]   img_reg_array_39_9_imag;
  reg        [17:0]   img_reg_array_39_10_real;
  reg        [17:0]   img_reg_array_39_10_imag;
  reg        [17:0]   img_reg_array_39_11_real;
  reg        [17:0]   img_reg_array_39_11_imag;
  reg        [17:0]   img_reg_array_39_12_real;
  reg        [17:0]   img_reg_array_39_12_imag;
  reg        [17:0]   img_reg_array_39_13_real;
  reg        [17:0]   img_reg_array_39_13_imag;
  reg        [17:0]   img_reg_array_39_14_real;
  reg        [17:0]   img_reg_array_39_14_imag;
  reg        [17:0]   img_reg_array_39_15_real;
  reg        [17:0]   img_reg_array_39_15_imag;
  reg        [17:0]   img_reg_array_39_16_real;
  reg        [17:0]   img_reg_array_39_16_imag;
  reg        [17:0]   img_reg_array_39_17_real;
  reg        [17:0]   img_reg_array_39_17_imag;
  reg        [17:0]   img_reg_array_39_18_real;
  reg        [17:0]   img_reg_array_39_18_imag;
  reg        [17:0]   img_reg_array_39_19_real;
  reg        [17:0]   img_reg_array_39_19_imag;
  reg        [17:0]   img_reg_array_39_20_real;
  reg        [17:0]   img_reg_array_39_20_imag;
  reg        [17:0]   img_reg_array_39_21_real;
  reg        [17:0]   img_reg_array_39_21_imag;
  reg        [17:0]   img_reg_array_39_22_real;
  reg        [17:0]   img_reg_array_39_22_imag;
  reg        [17:0]   img_reg_array_39_23_real;
  reg        [17:0]   img_reg_array_39_23_imag;
  reg        [17:0]   img_reg_array_39_24_real;
  reg        [17:0]   img_reg_array_39_24_imag;
  reg        [17:0]   img_reg_array_39_25_real;
  reg        [17:0]   img_reg_array_39_25_imag;
  reg        [17:0]   img_reg_array_39_26_real;
  reg        [17:0]   img_reg_array_39_26_imag;
  reg        [17:0]   img_reg_array_39_27_real;
  reg        [17:0]   img_reg_array_39_27_imag;
  reg        [17:0]   img_reg_array_39_28_real;
  reg        [17:0]   img_reg_array_39_28_imag;
  reg        [17:0]   img_reg_array_39_29_real;
  reg        [17:0]   img_reg_array_39_29_imag;
  reg        [17:0]   img_reg_array_39_30_real;
  reg        [17:0]   img_reg_array_39_30_imag;
  reg        [17:0]   img_reg_array_39_31_real;
  reg        [17:0]   img_reg_array_39_31_imag;
  reg        [17:0]   img_reg_array_39_32_real;
  reg        [17:0]   img_reg_array_39_32_imag;
  reg        [17:0]   img_reg_array_39_33_real;
  reg        [17:0]   img_reg_array_39_33_imag;
  reg        [17:0]   img_reg_array_39_34_real;
  reg        [17:0]   img_reg_array_39_34_imag;
  reg        [17:0]   img_reg_array_39_35_real;
  reg        [17:0]   img_reg_array_39_35_imag;
  reg        [17:0]   img_reg_array_39_36_real;
  reg        [17:0]   img_reg_array_39_36_imag;
  reg        [17:0]   img_reg_array_39_37_real;
  reg        [17:0]   img_reg_array_39_37_imag;
  reg        [17:0]   img_reg_array_39_38_real;
  reg        [17:0]   img_reg_array_39_38_imag;
  reg        [17:0]   img_reg_array_39_39_real;
  reg        [17:0]   img_reg_array_39_39_imag;
  reg        [17:0]   img_reg_array_39_40_real;
  reg        [17:0]   img_reg_array_39_40_imag;
  reg        [17:0]   img_reg_array_39_41_real;
  reg        [17:0]   img_reg_array_39_41_imag;
  reg        [17:0]   img_reg_array_39_42_real;
  reg        [17:0]   img_reg_array_39_42_imag;
  reg        [17:0]   img_reg_array_39_43_real;
  reg        [17:0]   img_reg_array_39_43_imag;
  reg        [17:0]   img_reg_array_39_44_real;
  reg        [17:0]   img_reg_array_39_44_imag;
  reg        [17:0]   img_reg_array_39_45_real;
  reg        [17:0]   img_reg_array_39_45_imag;
  reg        [17:0]   img_reg_array_39_46_real;
  reg        [17:0]   img_reg_array_39_46_imag;
  reg        [17:0]   img_reg_array_39_47_real;
  reg        [17:0]   img_reg_array_39_47_imag;
  reg        [17:0]   img_reg_array_39_48_real;
  reg        [17:0]   img_reg_array_39_48_imag;
  reg        [17:0]   img_reg_array_39_49_real;
  reg        [17:0]   img_reg_array_39_49_imag;
  reg        [17:0]   img_reg_array_39_50_real;
  reg        [17:0]   img_reg_array_39_50_imag;
  reg        [17:0]   img_reg_array_39_51_real;
  reg        [17:0]   img_reg_array_39_51_imag;
  reg        [17:0]   img_reg_array_39_52_real;
  reg        [17:0]   img_reg_array_39_52_imag;
  reg        [17:0]   img_reg_array_39_53_real;
  reg        [17:0]   img_reg_array_39_53_imag;
  reg        [17:0]   img_reg_array_39_54_real;
  reg        [17:0]   img_reg_array_39_54_imag;
  reg        [17:0]   img_reg_array_39_55_real;
  reg        [17:0]   img_reg_array_39_55_imag;
  reg        [17:0]   img_reg_array_39_56_real;
  reg        [17:0]   img_reg_array_39_56_imag;
  reg        [17:0]   img_reg_array_39_57_real;
  reg        [17:0]   img_reg_array_39_57_imag;
  reg        [17:0]   img_reg_array_39_58_real;
  reg        [17:0]   img_reg_array_39_58_imag;
  reg        [17:0]   img_reg_array_39_59_real;
  reg        [17:0]   img_reg_array_39_59_imag;
  reg        [17:0]   img_reg_array_39_60_real;
  reg        [17:0]   img_reg_array_39_60_imag;
  reg        [17:0]   img_reg_array_39_61_real;
  reg        [17:0]   img_reg_array_39_61_imag;
  reg        [17:0]   img_reg_array_39_62_real;
  reg        [17:0]   img_reg_array_39_62_imag;
  reg        [17:0]   img_reg_array_39_63_real;
  reg        [17:0]   img_reg_array_39_63_imag;
  reg        [17:0]   img_reg_array_40_0_real;
  reg        [17:0]   img_reg_array_40_0_imag;
  reg        [17:0]   img_reg_array_40_1_real;
  reg        [17:0]   img_reg_array_40_1_imag;
  reg        [17:0]   img_reg_array_40_2_real;
  reg        [17:0]   img_reg_array_40_2_imag;
  reg        [17:0]   img_reg_array_40_3_real;
  reg        [17:0]   img_reg_array_40_3_imag;
  reg        [17:0]   img_reg_array_40_4_real;
  reg        [17:0]   img_reg_array_40_4_imag;
  reg        [17:0]   img_reg_array_40_5_real;
  reg        [17:0]   img_reg_array_40_5_imag;
  reg        [17:0]   img_reg_array_40_6_real;
  reg        [17:0]   img_reg_array_40_6_imag;
  reg        [17:0]   img_reg_array_40_7_real;
  reg        [17:0]   img_reg_array_40_7_imag;
  reg        [17:0]   img_reg_array_40_8_real;
  reg        [17:0]   img_reg_array_40_8_imag;
  reg        [17:0]   img_reg_array_40_9_real;
  reg        [17:0]   img_reg_array_40_9_imag;
  reg        [17:0]   img_reg_array_40_10_real;
  reg        [17:0]   img_reg_array_40_10_imag;
  reg        [17:0]   img_reg_array_40_11_real;
  reg        [17:0]   img_reg_array_40_11_imag;
  reg        [17:0]   img_reg_array_40_12_real;
  reg        [17:0]   img_reg_array_40_12_imag;
  reg        [17:0]   img_reg_array_40_13_real;
  reg        [17:0]   img_reg_array_40_13_imag;
  reg        [17:0]   img_reg_array_40_14_real;
  reg        [17:0]   img_reg_array_40_14_imag;
  reg        [17:0]   img_reg_array_40_15_real;
  reg        [17:0]   img_reg_array_40_15_imag;
  reg        [17:0]   img_reg_array_40_16_real;
  reg        [17:0]   img_reg_array_40_16_imag;
  reg        [17:0]   img_reg_array_40_17_real;
  reg        [17:0]   img_reg_array_40_17_imag;
  reg        [17:0]   img_reg_array_40_18_real;
  reg        [17:0]   img_reg_array_40_18_imag;
  reg        [17:0]   img_reg_array_40_19_real;
  reg        [17:0]   img_reg_array_40_19_imag;
  reg        [17:0]   img_reg_array_40_20_real;
  reg        [17:0]   img_reg_array_40_20_imag;
  reg        [17:0]   img_reg_array_40_21_real;
  reg        [17:0]   img_reg_array_40_21_imag;
  reg        [17:0]   img_reg_array_40_22_real;
  reg        [17:0]   img_reg_array_40_22_imag;
  reg        [17:0]   img_reg_array_40_23_real;
  reg        [17:0]   img_reg_array_40_23_imag;
  reg        [17:0]   img_reg_array_40_24_real;
  reg        [17:0]   img_reg_array_40_24_imag;
  reg        [17:0]   img_reg_array_40_25_real;
  reg        [17:0]   img_reg_array_40_25_imag;
  reg        [17:0]   img_reg_array_40_26_real;
  reg        [17:0]   img_reg_array_40_26_imag;
  reg        [17:0]   img_reg_array_40_27_real;
  reg        [17:0]   img_reg_array_40_27_imag;
  reg        [17:0]   img_reg_array_40_28_real;
  reg        [17:0]   img_reg_array_40_28_imag;
  reg        [17:0]   img_reg_array_40_29_real;
  reg        [17:0]   img_reg_array_40_29_imag;
  reg        [17:0]   img_reg_array_40_30_real;
  reg        [17:0]   img_reg_array_40_30_imag;
  reg        [17:0]   img_reg_array_40_31_real;
  reg        [17:0]   img_reg_array_40_31_imag;
  reg        [17:0]   img_reg_array_40_32_real;
  reg        [17:0]   img_reg_array_40_32_imag;
  reg        [17:0]   img_reg_array_40_33_real;
  reg        [17:0]   img_reg_array_40_33_imag;
  reg        [17:0]   img_reg_array_40_34_real;
  reg        [17:0]   img_reg_array_40_34_imag;
  reg        [17:0]   img_reg_array_40_35_real;
  reg        [17:0]   img_reg_array_40_35_imag;
  reg        [17:0]   img_reg_array_40_36_real;
  reg        [17:0]   img_reg_array_40_36_imag;
  reg        [17:0]   img_reg_array_40_37_real;
  reg        [17:0]   img_reg_array_40_37_imag;
  reg        [17:0]   img_reg_array_40_38_real;
  reg        [17:0]   img_reg_array_40_38_imag;
  reg        [17:0]   img_reg_array_40_39_real;
  reg        [17:0]   img_reg_array_40_39_imag;
  reg        [17:0]   img_reg_array_40_40_real;
  reg        [17:0]   img_reg_array_40_40_imag;
  reg        [17:0]   img_reg_array_40_41_real;
  reg        [17:0]   img_reg_array_40_41_imag;
  reg        [17:0]   img_reg_array_40_42_real;
  reg        [17:0]   img_reg_array_40_42_imag;
  reg        [17:0]   img_reg_array_40_43_real;
  reg        [17:0]   img_reg_array_40_43_imag;
  reg        [17:0]   img_reg_array_40_44_real;
  reg        [17:0]   img_reg_array_40_44_imag;
  reg        [17:0]   img_reg_array_40_45_real;
  reg        [17:0]   img_reg_array_40_45_imag;
  reg        [17:0]   img_reg_array_40_46_real;
  reg        [17:0]   img_reg_array_40_46_imag;
  reg        [17:0]   img_reg_array_40_47_real;
  reg        [17:0]   img_reg_array_40_47_imag;
  reg        [17:0]   img_reg_array_40_48_real;
  reg        [17:0]   img_reg_array_40_48_imag;
  reg        [17:0]   img_reg_array_40_49_real;
  reg        [17:0]   img_reg_array_40_49_imag;
  reg        [17:0]   img_reg_array_40_50_real;
  reg        [17:0]   img_reg_array_40_50_imag;
  reg        [17:0]   img_reg_array_40_51_real;
  reg        [17:0]   img_reg_array_40_51_imag;
  reg        [17:0]   img_reg_array_40_52_real;
  reg        [17:0]   img_reg_array_40_52_imag;
  reg        [17:0]   img_reg_array_40_53_real;
  reg        [17:0]   img_reg_array_40_53_imag;
  reg        [17:0]   img_reg_array_40_54_real;
  reg        [17:0]   img_reg_array_40_54_imag;
  reg        [17:0]   img_reg_array_40_55_real;
  reg        [17:0]   img_reg_array_40_55_imag;
  reg        [17:0]   img_reg_array_40_56_real;
  reg        [17:0]   img_reg_array_40_56_imag;
  reg        [17:0]   img_reg_array_40_57_real;
  reg        [17:0]   img_reg_array_40_57_imag;
  reg        [17:0]   img_reg_array_40_58_real;
  reg        [17:0]   img_reg_array_40_58_imag;
  reg        [17:0]   img_reg_array_40_59_real;
  reg        [17:0]   img_reg_array_40_59_imag;
  reg        [17:0]   img_reg_array_40_60_real;
  reg        [17:0]   img_reg_array_40_60_imag;
  reg        [17:0]   img_reg_array_40_61_real;
  reg        [17:0]   img_reg_array_40_61_imag;
  reg        [17:0]   img_reg_array_40_62_real;
  reg        [17:0]   img_reg_array_40_62_imag;
  reg        [17:0]   img_reg_array_40_63_real;
  reg        [17:0]   img_reg_array_40_63_imag;
  reg        [17:0]   img_reg_array_41_0_real;
  reg        [17:0]   img_reg_array_41_0_imag;
  reg        [17:0]   img_reg_array_41_1_real;
  reg        [17:0]   img_reg_array_41_1_imag;
  reg        [17:0]   img_reg_array_41_2_real;
  reg        [17:0]   img_reg_array_41_2_imag;
  reg        [17:0]   img_reg_array_41_3_real;
  reg        [17:0]   img_reg_array_41_3_imag;
  reg        [17:0]   img_reg_array_41_4_real;
  reg        [17:0]   img_reg_array_41_4_imag;
  reg        [17:0]   img_reg_array_41_5_real;
  reg        [17:0]   img_reg_array_41_5_imag;
  reg        [17:0]   img_reg_array_41_6_real;
  reg        [17:0]   img_reg_array_41_6_imag;
  reg        [17:0]   img_reg_array_41_7_real;
  reg        [17:0]   img_reg_array_41_7_imag;
  reg        [17:0]   img_reg_array_41_8_real;
  reg        [17:0]   img_reg_array_41_8_imag;
  reg        [17:0]   img_reg_array_41_9_real;
  reg        [17:0]   img_reg_array_41_9_imag;
  reg        [17:0]   img_reg_array_41_10_real;
  reg        [17:0]   img_reg_array_41_10_imag;
  reg        [17:0]   img_reg_array_41_11_real;
  reg        [17:0]   img_reg_array_41_11_imag;
  reg        [17:0]   img_reg_array_41_12_real;
  reg        [17:0]   img_reg_array_41_12_imag;
  reg        [17:0]   img_reg_array_41_13_real;
  reg        [17:0]   img_reg_array_41_13_imag;
  reg        [17:0]   img_reg_array_41_14_real;
  reg        [17:0]   img_reg_array_41_14_imag;
  reg        [17:0]   img_reg_array_41_15_real;
  reg        [17:0]   img_reg_array_41_15_imag;
  reg        [17:0]   img_reg_array_41_16_real;
  reg        [17:0]   img_reg_array_41_16_imag;
  reg        [17:0]   img_reg_array_41_17_real;
  reg        [17:0]   img_reg_array_41_17_imag;
  reg        [17:0]   img_reg_array_41_18_real;
  reg        [17:0]   img_reg_array_41_18_imag;
  reg        [17:0]   img_reg_array_41_19_real;
  reg        [17:0]   img_reg_array_41_19_imag;
  reg        [17:0]   img_reg_array_41_20_real;
  reg        [17:0]   img_reg_array_41_20_imag;
  reg        [17:0]   img_reg_array_41_21_real;
  reg        [17:0]   img_reg_array_41_21_imag;
  reg        [17:0]   img_reg_array_41_22_real;
  reg        [17:0]   img_reg_array_41_22_imag;
  reg        [17:0]   img_reg_array_41_23_real;
  reg        [17:0]   img_reg_array_41_23_imag;
  reg        [17:0]   img_reg_array_41_24_real;
  reg        [17:0]   img_reg_array_41_24_imag;
  reg        [17:0]   img_reg_array_41_25_real;
  reg        [17:0]   img_reg_array_41_25_imag;
  reg        [17:0]   img_reg_array_41_26_real;
  reg        [17:0]   img_reg_array_41_26_imag;
  reg        [17:0]   img_reg_array_41_27_real;
  reg        [17:0]   img_reg_array_41_27_imag;
  reg        [17:0]   img_reg_array_41_28_real;
  reg        [17:0]   img_reg_array_41_28_imag;
  reg        [17:0]   img_reg_array_41_29_real;
  reg        [17:0]   img_reg_array_41_29_imag;
  reg        [17:0]   img_reg_array_41_30_real;
  reg        [17:0]   img_reg_array_41_30_imag;
  reg        [17:0]   img_reg_array_41_31_real;
  reg        [17:0]   img_reg_array_41_31_imag;
  reg        [17:0]   img_reg_array_41_32_real;
  reg        [17:0]   img_reg_array_41_32_imag;
  reg        [17:0]   img_reg_array_41_33_real;
  reg        [17:0]   img_reg_array_41_33_imag;
  reg        [17:0]   img_reg_array_41_34_real;
  reg        [17:0]   img_reg_array_41_34_imag;
  reg        [17:0]   img_reg_array_41_35_real;
  reg        [17:0]   img_reg_array_41_35_imag;
  reg        [17:0]   img_reg_array_41_36_real;
  reg        [17:0]   img_reg_array_41_36_imag;
  reg        [17:0]   img_reg_array_41_37_real;
  reg        [17:0]   img_reg_array_41_37_imag;
  reg        [17:0]   img_reg_array_41_38_real;
  reg        [17:0]   img_reg_array_41_38_imag;
  reg        [17:0]   img_reg_array_41_39_real;
  reg        [17:0]   img_reg_array_41_39_imag;
  reg        [17:0]   img_reg_array_41_40_real;
  reg        [17:0]   img_reg_array_41_40_imag;
  reg        [17:0]   img_reg_array_41_41_real;
  reg        [17:0]   img_reg_array_41_41_imag;
  reg        [17:0]   img_reg_array_41_42_real;
  reg        [17:0]   img_reg_array_41_42_imag;
  reg        [17:0]   img_reg_array_41_43_real;
  reg        [17:0]   img_reg_array_41_43_imag;
  reg        [17:0]   img_reg_array_41_44_real;
  reg        [17:0]   img_reg_array_41_44_imag;
  reg        [17:0]   img_reg_array_41_45_real;
  reg        [17:0]   img_reg_array_41_45_imag;
  reg        [17:0]   img_reg_array_41_46_real;
  reg        [17:0]   img_reg_array_41_46_imag;
  reg        [17:0]   img_reg_array_41_47_real;
  reg        [17:0]   img_reg_array_41_47_imag;
  reg        [17:0]   img_reg_array_41_48_real;
  reg        [17:0]   img_reg_array_41_48_imag;
  reg        [17:0]   img_reg_array_41_49_real;
  reg        [17:0]   img_reg_array_41_49_imag;
  reg        [17:0]   img_reg_array_41_50_real;
  reg        [17:0]   img_reg_array_41_50_imag;
  reg        [17:0]   img_reg_array_41_51_real;
  reg        [17:0]   img_reg_array_41_51_imag;
  reg        [17:0]   img_reg_array_41_52_real;
  reg        [17:0]   img_reg_array_41_52_imag;
  reg        [17:0]   img_reg_array_41_53_real;
  reg        [17:0]   img_reg_array_41_53_imag;
  reg        [17:0]   img_reg_array_41_54_real;
  reg        [17:0]   img_reg_array_41_54_imag;
  reg        [17:0]   img_reg_array_41_55_real;
  reg        [17:0]   img_reg_array_41_55_imag;
  reg        [17:0]   img_reg_array_41_56_real;
  reg        [17:0]   img_reg_array_41_56_imag;
  reg        [17:0]   img_reg_array_41_57_real;
  reg        [17:0]   img_reg_array_41_57_imag;
  reg        [17:0]   img_reg_array_41_58_real;
  reg        [17:0]   img_reg_array_41_58_imag;
  reg        [17:0]   img_reg_array_41_59_real;
  reg        [17:0]   img_reg_array_41_59_imag;
  reg        [17:0]   img_reg_array_41_60_real;
  reg        [17:0]   img_reg_array_41_60_imag;
  reg        [17:0]   img_reg_array_41_61_real;
  reg        [17:0]   img_reg_array_41_61_imag;
  reg        [17:0]   img_reg_array_41_62_real;
  reg        [17:0]   img_reg_array_41_62_imag;
  reg        [17:0]   img_reg_array_41_63_real;
  reg        [17:0]   img_reg_array_41_63_imag;
  reg        [17:0]   img_reg_array_42_0_real;
  reg        [17:0]   img_reg_array_42_0_imag;
  reg        [17:0]   img_reg_array_42_1_real;
  reg        [17:0]   img_reg_array_42_1_imag;
  reg        [17:0]   img_reg_array_42_2_real;
  reg        [17:0]   img_reg_array_42_2_imag;
  reg        [17:0]   img_reg_array_42_3_real;
  reg        [17:0]   img_reg_array_42_3_imag;
  reg        [17:0]   img_reg_array_42_4_real;
  reg        [17:0]   img_reg_array_42_4_imag;
  reg        [17:0]   img_reg_array_42_5_real;
  reg        [17:0]   img_reg_array_42_5_imag;
  reg        [17:0]   img_reg_array_42_6_real;
  reg        [17:0]   img_reg_array_42_6_imag;
  reg        [17:0]   img_reg_array_42_7_real;
  reg        [17:0]   img_reg_array_42_7_imag;
  reg        [17:0]   img_reg_array_42_8_real;
  reg        [17:0]   img_reg_array_42_8_imag;
  reg        [17:0]   img_reg_array_42_9_real;
  reg        [17:0]   img_reg_array_42_9_imag;
  reg        [17:0]   img_reg_array_42_10_real;
  reg        [17:0]   img_reg_array_42_10_imag;
  reg        [17:0]   img_reg_array_42_11_real;
  reg        [17:0]   img_reg_array_42_11_imag;
  reg        [17:0]   img_reg_array_42_12_real;
  reg        [17:0]   img_reg_array_42_12_imag;
  reg        [17:0]   img_reg_array_42_13_real;
  reg        [17:0]   img_reg_array_42_13_imag;
  reg        [17:0]   img_reg_array_42_14_real;
  reg        [17:0]   img_reg_array_42_14_imag;
  reg        [17:0]   img_reg_array_42_15_real;
  reg        [17:0]   img_reg_array_42_15_imag;
  reg        [17:0]   img_reg_array_42_16_real;
  reg        [17:0]   img_reg_array_42_16_imag;
  reg        [17:0]   img_reg_array_42_17_real;
  reg        [17:0]   img_reg_array_42_17_imag;
  reg        [17:0]   img_reg_array_42_18_real;
  reg        [17:0]   img_reg_array_42_18_imag;
  reg        [17:0]   img_reg_array_42_19_real;
  reg        [17:0]   img_reg_array_42_19_imag;
  reg        [17:0]   img_reg_array_42_20_real;
  reg        [17:0]   img_reg_array_42_20_imag;
  reg        [17:0]   img_reg_array_42_21_real;
  reg        [17:0]   img_reg_array_42_21_imag;
  reg        [17:0]   img_reg_array_42_22_real;
  reg        [17:0]   img_reg_array_42_22_imag;
  reg        [17:0]   img_reg_array_42_23_real;
  reg        [17:0]   img_reg_array_42_23_imag;
  reg        [17:0]   img_reg_array_42_24_real;
  reg        [17:0]   img_reg_array_42_24_imag;
  reg        [17:0]   img_reg_array_42_25_real;
  reg        [17:0]   img_reg_array_42_25_imag;
  reg        [17:0]   img_reg_array_42_26_real;
  reg        [17:0]   img_reg_array_42_26_imag;
  reg        [17:0]   img_reg_array_42_27_real;
  reg        [17:0]   img_reg_array_42_27_imag;
  reg        [17:0]   img_reg_array_42_28_real;
  reg        [17:0]   img_reg_array_42_28_imag;
  reg        [17:0]   img_reg_array_42_29_real;
  reg        [17:0]   img_reg_array_42_29_imag;
  reg        [17:0]   img_reg_array_42_30_real;
  reg        [17:0]   img_reg_array_42_30_imag;
  reg        [17:0]   img_reg_array_42_31_real;
  reg        [17:0]   img_reg_array_42_31_imag;
  reg        [17:0]   img_reg_array_42_32_real;
  reg        [17:0]   img_reg_array_42_32_imag;
  reg        [17:0]   img_reg_array_42_33_real;
  reg        [17:0]   img_reg_array_42_33_imag;
  reg        [17:0]   img_reg_array_42_34_real;
  reg        [17:0]   img_reg_array_42_34_imag;
  reg        [17:0]   img_reg_array_42_35_real;
  reg        [17:0]   img_reg_array_42_35_imag;
  reg        [17:0]   img_reg_array_42_36_real;
  reg        [17:0]   img_reg_array_42_36_imag;
  reg        [17:0]   img_reg_array_42_37_real;
  reg        [17:0]   img_reg_array_42_37_imag;
  reg        [17:0]   img_reg_array_42_38_real;
  reg        [17:0]   img_reg_array_42_38_imag;
  reg        [17:0]   img_reg_array_42_39_real;
  reg        [17:0]   img_reg_array_42_39_imag;
  reg        [17:0]   img_reg_array_42_40_real;
  reg        [17:0]   img_reg_array_42_40_imag;
  reg        [17:0]   img_reg_array_42_41_real;
  reg        [17:0]   img_reg_array_42_41_imag;
  reg        [17:0]   img_reg_array_42_42_real;
  reg        [17:0]   img_reg_array_42_42_imag;
  reg        [17:0]   img_reg_array_42_43_real;
  reg        [17:0]   img_reg_array_42_43_imag;
  reg        [17:0]   img_reg_array_42_44_real;
  reg        [17:0]   img_reg_array_42_44_imag;
  reg        [17:0]   img_reg_array_42_45_real;
  reg        [17:0]   img_reg_array_42_45_imag;
  reg        [17:0]   img_reg_array_42_46_real;
  reg        [17:0]   img_reg_array_42_46_imag;
  reg        [17:0]   img_reg_array_42_47_real;
  reg        [17:0]   img_reg_array_42_47_imag;
  reg        [17:0]   img_reg_array_42_48_real;
  reg        [17:0]   img_reg_array_42_48_imag;
  reg        [17:0]   img_reg_array_42_49_real;
  reg        [17:0]   img_reg_array_42_49_imag;
  reg        [17:0]   img_reg_array_42_50_real;
  reg        [17:0]   img_reg_array_42_50_imag;
  reg        [17:0]   img_reg_array_42_51_real;
  reg        [17:0]   img_reg_array_42_51_imag;
  reg        [17:0]   img_reg_array_42_52_real;
  reg        [17:0]   img_reg_array_42_52_imag;
  reg        [17:0]   img_reg_array_42_53_real;
  reg        [17:0]   img_reg_array_42_53_imag;
  reg        [17:0]   img_reg_array_42_54_real;
  reg        [17:0]   img_reg_array_42_54_imag;
  reg        [17:0]   img_reg_array_42_55_real;
  reg        [17:0]   img_reg_array_42_55_imag;
  reg        [17:0]   img_reg_array_42_56_real;
  reg        [17:0]   img_reg_array_42_56_imag;
  reg        [17:0]   img_reg_array_42_57_real;
  reg        [17:0]   img_reg_array_42_57_imag;
  reg        [17:0]   img_reg_array_42_58_real;
  reg        [17:0]   img_reg_array_42_58_imag;
  reg        [17:0]   img_reg_array_42_59_real;
  reg        [17:0]   img_reg_array_42_59_imag;
  reg        [17:0]   img_reg_array_42_60_real;
  reg        [17:0]   img_reg_array_42_60_imag;
  reg        [17:0]   img_reg_array_42_61_real;
  reg        [17:0]   img_reg_array_42_61_imag;
  reg        [17:0]   img_reg_array_42_62_real;
  reg        [17:0]   img_reg_array_42_62_imag;
  reg        [17:0]   img_reg_array_42_63_real;
  reg        [17:0]   img_reg_array_42_63_imag;
  reg        [17:0]   img_reg_array_43_0_real;
  reg        [17:0]   img_reg_array_43_0_imag;
  reg        [17:0]   img_reg_array_43_1_real;
  reg        [17:0]   img_reg_array_43_1_imag;
  reg        [17:0]   img_reg_array_43_2_real;
  reg        [17:0]   img_reg_array_43_2_imag;
  reg        [17:0]   img_reg_array_43_3_real;
  reg        [17:0]   img_reg_array_43_3_imag;
  reg        [17:0]   img_reg_array_43_4_real;
  reg        [17:0]   img_reg_array_43_4_imag;
  reg        [17:0]   img_reg_array_43_5_real;
  reg        [17:0]   img_reg_array_43_5_imag;
  reg        [17:0]   img_reg_array_43_6_real;
  reg        [17:0]   img_reg_array_43_6_imag;
  reg        [17:0]   img_reg_array_43_7_real;
  reg        [17:0]   img_reg_array_43_7_imag;
  reg        [17:0]   img_reg_array_43_8_real;
  reg        [17:0]   img_reg_array_43_8_imag;
  reg        [17:0]   img_reg_array_43_9_real;
  reg        [17:0]   img_reg_array_43_9_imag;
  reg        [17:0]   img_reg_array_43_10_real;
  reg        [17:0]   img_reg_array_43_10_imag;
  reg        [17:0]   img_reg_array_43_11_real;
  reg        [17:0]   img_reg_array_43_11_imag;
  reg        [17:0]   img_reg_array_43_12_real;
  reg        [17:0]   img_reg_array_43_12_imag;
  reg        [17:0]   img_reg_array_43_13_real;
  reg        [17:0]   img_reg_array_43_13_imag;
  reg        [17:0]   img_reg_array_43_14_real;
  reg        [17:0]   img_reg_array_43_14_imag;
  reg        [17:0]   img_reg_array_43_15_real;
  reg        [17:0]   img_reg_array_43_15_imag;
  reg        [17:0]   img_reg_array_43_16_real;
  reg        [17:0]   img_reg_array_43_16_imag;
  reg        [17:0]   img_reg_array_43_17_real;
  reg        [17:0]   img_reg_array_43_17_imag;
  reg        [17:0]   img_reg_array_43_18_real;
  reg        [17:0]   img_reg_array_43_18_imag;
  reg        [17:0]   img_reg_array_43_19_real;
  reg        [17:0]   img_reg_array_43_19_imag;
  reg        [17:0]   img_reg_array_43_20_real;
  reg        [17:0]   img_reg_array_43_20_imag;
  reg        [17:0]   img_reg_array_43_21_real;
  reg        [17:0]   img_reg_array_43_21_imag;
  reg        [17:0]   img_reg_array_43_22_real;
  reg        [17:0]   img_reg_array_43_22_imag;
  reg        [17:0]   img_reg_array_43_23_real;
  reg        [17:0]   img_reg_array_43_23_imag;
  reg        [17:0]   img_reg_array_43_24_real;
  reg        [17:0]   img_reg_array_43_24_imag;
  reg        [17:0]   img_reg_array_43_25_real;
  reg        [17:0]   img_reg_array_43_25_imag;
  reg        [17:0]   img_reg_array_43_26_real;
  reg        [17:0]   img_reg_array_43_26_imag;
  reg        [17:0]   img_reg_array_43_27_real;
  reg        [17:0]   img_reg_array_43_27_imag;
  reg        [17:0]   img_reg_array_43_28_real;
  reg        [17:0]   img_reg_array_43_28_imag;
  reg        [17:0]   img_reg_array_43_29_real;
  reg        [17:0]   img_reg_array_43_29_imag;
  reg        [17:0]   img_reg_array_43_30_real;
  reg        [17:0]   img_reg_array_43_30_imag;
  reg        [17:0]   img_reg_array_43_31_real;
  reg        [17:0]   img_reg_array_43_31_imag;
  reg        [17:0]   img_reg_array_43_32_real;
  reg        [17:0]   img_reg_array_43_32_imag;
  reg        [17:0]   img_reg_array_43_33_real;
  reg        [17:0]   img_reg_array_43_33_imag;
  reg        [17:0]   img_reg_array_43_34_real;
  reg        [17:0]   img_reg_array_43_34_imag;
  reg        [17:0]   img_reg_array_43_35_real;
  reg        [17:0]   img_reg_array_43_35_imag;
  reg        [17:0]   img_reg_array_43_36_real;
  reg        [17:0]   img_reg_array_43_36_imag;
  reg        [17:0]   img_reg_array_43_37_real;
  reg        [17:0]   img_reg_array_43_37_imag;
  reg        [17:0]   img_reg_array_43_38_real;
  reg        [17:0]   img_reg_array_43_38_imag;
  reg        [17:0]   img_reg_array_43_39_real;
  reg        [17:0]   img_reg_array_43_39_imag;
  reg        [17:0]   img_reg_array_43_40_real;
  reg        [17:0]   img_reg_array_43_40_imag;
  reg        [17:0]   img_reg_array_43_41_real;
  reg        [17:0]   img_reg_array_43_41_imag;
  reg        [17:0]   img_reg_array_43_42_real;
  reg        [17:0]   img_reg_array_43_42_imag;
  reg        [17:0]   img_reg_array_43_43_real;
  reg        [17:0]   img_reg_array_43_43_imag;
  reg        [17:0]   img_reg_array_43_44_real;
  reg        [17:0]   img_reg_array_43_44_imag;
  reg        [17:0]   img_reg_array_43_45_real;
  reg        [17:0]   img_reg_array_43_45_imag;
  reg        [17:0]   img_reg_array_43_46_real;
  reg        [17:0]   img_reg_array_43_46_imag;
  reg        [17:0]   img_reg_array_43_47_real;
  reg        [17:0]   img_reg_array_43_47_imag;
  reg        [17:0]   img_reg_array_43_48_real;
  reg        [17:0]   img_reg_array_43_48_imag;
  reg        [17:0]   img_reg_array_43_49_real;
  reg        [17:0]   img_reg_array_43_49_imag;
  reg        [17:0]   img_reg_array_43_50_real;
  reg        [17:0]   img_reg_array_43_50_imag;
  reg        [17:0]   img_reg_array_43_51_real;
  reg        [17:0]   img_reg_array_43_51_imag;
  reg        [17:0]   img_reg_array_43_52_real;
  reg        [17:0]   img_reg_array_43_52_imag;
  reg        [17:0]   img_reg_array_43_53_real;
  reg        [17:0]   img_reg_array_43_53_imag;
  reg        [17:0]   img_reg_array_43_54_real;
  reg        [17:0]   img_reg_array_43_54_imag;
  reg        [17:0]   img_reg_array_43_55_real;
  reg        [17:0]   img_reg_array_43_55_imag;
  reg        [17:0]   img_reg_array_43_56_real;
  reg        [17:0]   img_reg_array_43_56_imag;
  reg        [17:0]   img_reg_array_43_57_real;
  reg        [17:0]   img_reg_array_43_57_imag;
  reg        [17:0]   img_reg_array_43_58_real;
  reg        [17:0]   img_reg_array_43_58_imag;
  reg        [17:0]   img_reg_array_43_59_real;
  reg        [17:0]   img_reg_array_43_59_imag;
  reg        [17:0]   img_reg_array_43_60_real;
  reg        [17:0]   img_reg_array_43_60_imag;
  reg        [17:0]   img_reg_array_43_61_real;
  reg        [17:0]   img_reg_array_43_61_imag;
  reg        [17:0]   img_reg_array_43_62_real;
  reg        [17:0]   img_reg_array_43_62_imag;
  reg        [17:0]   img_reg_array_43_63_real;
  reg        [17:0]   img_reg_array_43_63_imag;
  reg        [17:0]   img_reg_array_44_0_real;
  reg        [17:0]   img_reg_array_44_0_imag;
  reg        [17:0]   img_reg_array_44_1_real;
  reg        [17:0]   img_reg_array_44_1_imag;
  reg        [17:0]   img_reg_array_44_2_real;
  reg        [17:0]   img_reg_array_44_2_imag;
  reg        [17:0]   img_reg_array_44_3_real;
  reg        [17:0]   img_reg_array_44_3_imag;
  reg        [17:0]   img_reg_array_44_4_real;
  reg        [17:0]   img_reg_array_44_4_imag;
  reg        [17:0]   img_reg_array_44_5_real;
  reg        [17:0]   img_reg_array_44_5_imag;
  reg        [17:0]   img_reg_array_44_6_real;
  reg        [17:0]   img_reg_array_44_6_imag;
  reg        [17:0]   img_reg_array_44_7_real;
  reg        [17:0]   img_reg_array_44_7_imag;
  reg        [17:0]   img_reg_array_44_8_real;
  reg        [17:0]   img_reg_array_44_8_imag;
  reg        [17:0]   img_reg_array_44_9_real;
  reg        [17:0]   img_reg_array_44_9_imag;
  reg        [17:0]   img_reg_array_44_10_real;
  reg        [17:0]   img_reg_array_44_10_imag;
  reg        [17:0]   img_reg_array_44_11_real;
  reg        [17:0]   img_reg_array_44_11_imag;
  reg        [17:0]   img_reg_array_44_12_real;
  reg        [17:0]   img_reg_array_44_12_imag;
  reg        [17:0]   img_reg_array_44_13_real;
  reg        [17:0]   img_reg_array_44_13_imag;
  reg        [17:0]   img_reg_array_44_14_real;
  reg        [17:0]   img_reg_array_44_14_imag;
  reg        [17:0]   img_reg_array_44_15_real;
  reg        [17:0]   img_reg_array_44_15_imag;
  reg        [17:0]   img_reg_array_44_16_real;
  reg        [17:0]   img_reg_array_44_16_imag;
  reg        [17:0]   img_reg_array_44_17_real;
  reg        [17:0]   img_reg_array_44_17_imag;
  reg        [17:0]   img_reg_array_44_18_real;
  reg        [17:0]   img_reg_array_44_18_imag;
  reg        [17:0]   img_reg_array_44_19_real;
  reg        [17:0]   img_reg_array_44_19_imag;
  reg        [17:0]   img_reg_array_44_20_real;
  reg        [17:0]   img_reg_array_44_20_imag;
  reg        [17:0]   img_reg_array_44_21_real;
  reg        [17:0]   img_reg_array_44_21_imag;
  reg        [17:0]   img_reg_array_44_22_real;
  reg        [17:0]   img_reg_array_44_22_imag;
  reg        [17:0]   img_reg_array_44_23_real;
  reg        [17:0]   img_reg_array_44_23_imag;
  reg        [17:0]   img_reg_array_44_24_real;
  reg        [17:0]   img_reg_array_44_24_imag;
  reg        [17:0]   img_reg_array_44_25_real;
  reg        [17:0]   img_reg_array_44_25_imag;
  reg        [17:0]   img_reg_array_44_26_real;
  reg        [17:0]   img_reg_array_44_26_imag;
  reg        [17:0]   img_reg_array_44_27_real;
  reg        [17:0]   img_reg_array_44_27_imag;
  reg        [17:0]   img_reg_array_44_28_real;
  reg        [17:0]   img_reg_array_44_28_imag;
  reg        [17:0]   img_reg_array_44_29_real;
  reg        [17:0]   img_reg_array_44_29_imag;
  reg        [17:0]   img_reg_array_44_30_real;
  reg        [17:0]   img_reg_array_44_30_imag;
  reg        [17:0]   img_reg_array_44_31_real;
  reg        [17:0]   img_reg_array_44_31_imag;
  reg        [17:0]   img_reg_array_44_32_real;
  reg        [17:0]   img_reg_array_44_32_imag;
  reg        [17:0]   img_reg_array_44_33_real;
  reg        [17:0]   img_reg_array_44_33_imag;
  reg        [17:0]   img_reg_array_44_34_real;
  reg        [17:0]   img_reg_array_44_34_imag;
  reg        [17:0]   img_reg_array_44_35_real;
  reg        [17:0]   img_reg_array_44_35_imag;
  reg        [17:0]   img_reg_array_44_36_real;
  reg        [17:0]   img_reg_array_44_36_imag;
  reg        [17:0]   img_reg_array_44_37_real;
  reg        [17:0]   img_reg_array_44_37_imag;
  reg        [17:0]   img_reg_array_44_38_real;
  reg        [17:0]   img_reg_array_44_38_imag;
  reg        [17:0]   img_reg_array_44_39_real;
  reg        [17:0]   img_reg_array_44_39_imag;
  reg        [17:0]   img_reg_array_44_40_real;
  reg        [17:0]   img_reg_array_44_40_imag;
  reg        [17:0]   img_reg_array_44_41_real;
  reg        [17:0]   img_reg_array_44_41_imag;
  reg        [17:0]   img_reg_array_44_42_real;
  reg        [17:0]   img_reg_array_44_42_imag;
  reg        [17:0]   img_reg_array_44_43_real;
  reg        [17:0]   img_reg_array_44_43_imag;
  reg        [17:0]   img_reg_array_44_44_real;
  reg        [17:0]   img_reg_array_44_44_imag;
  reg        [17:0]   img_reg_array_44_45_real;
  reg        [17:0]   img_reg_array_44_45_imag;
  reg        [17:0]   img_reg_array_44_46_real;
  reg        [17:0]   img_reg_array_44_46_imag;
  reg        [17:0]   img_reg_array_44_47_real;
  reg        [17:0]   img_reg_array_44_47_imag;
  reg        [17:0]   img_reg_array_44_48_real;
  reg        [17:0]   img_reg_array_44_48_imag;
  reg        [17:0]   img_reg_array_44_49_real;
  reg        [17:0]   img_reg_array_44_49_imag;
  reg        [17:0]   img_reg_array_44_50_real;
  reg        [17:0]   img_reg_array_44_50_imag;
  reg        [17:0]   img_reg_array_44_51_real;
  reg        [17:0]   img_reg_array_44_51_imag;
  reg        [17:0]   img_reg_array_44_52_real;
  reg        [17:0]   img_reg_array_44_52_imag;
  reg        [17:0]   img_reg_array_44_53_real;
  reg        [17:0]   img_reg_array_44_53_imag;
  reg        [17:0]   img_reg_array_44_54_real;
  reg        [17:0]   img_reg_array_44_54_imag;
  reg        [17:0]   img_reg_array_44_55_real;
  reg        [17:0]   img_reg_array_44_55_imag;
  reg        [17:0]   img_reg_array_44_56_real;
  reg        [17:0]   img_reg_array_44_56_imag;
  reg        [17:0]   img_reg_array_44_57_real;
  reg        [17:0]   img_reg_array_44_57_imag;
  reg        [17:0]   img_reg_array_44_58_real;
  reg        [17:0]   img_reg_array_44_58_imag;
  reg        [17:0]   img_reg_array_44_59_real;
  reg        [17:0]   img_reg_array_44_59_imag;
  reg        [17:0]   img_reg_array_44_60_real;
  reg        [17:0]   img_reg_array_44_60_imag;
  reg        [17:0]   img_reg_array_44_61_real;
  reg        [17:0]   img_reg_array_44_61_imag;
  reg        [17:0]   img_reg_array_44_62_real;
  reg        [17:0]   img_reg_array_44_62_imag;
  reg        [17:0]   img_reg_array_44_63_real;
  reg        [17:0]   img_reg_array_44_63_imag;
  reg        [17:0]   img_reg_array_45_0_real;
  reg        [17:0]   img_reg_array_45_0_imag;
  reg        [17:0]   img_reg_array_45_1_real;
  reg        [17:0]   img_reg_array_45_1_imag;
  reg        [17:0]   img_reg_array_45_2_real;
  reg        [17:0]   img_reg_array_45_2_imag;
  reg        [17:0]   img_reg_array_45_3_real;
  reg        [17:0]   img_reg_array_45_3_imag;
  reg        [17:0]   img_reg_array_45_4_real;
  reg        [17:0]   img_reg_array_45_4_imag;
  reg        [17:0]   img_reg_array_45_5_real;
  reg        [17:0]   img_reg_array_45_5_imag;
  reg        [17:0]   img_reg_array_45_6_real;
  reg        [17:0]   img_reg_array_45_6_imag;
  reg        [17:0]   img_reg_array_45_7_real;
  reg        [17:0]   img_reg_array_45_7_imag;
  reg        [17:0]   img_reg_array_45_8_real;
  reg        [17:0]   img_reg_array_45_8_imag;
  reg        [17:0]   img_reg_array_45_9_real;
  reg        [17:0]   img_reg_array_45_9_imag;
  reg        [17:0]   img_reg_array_45_10_real;
  reg        [17:0]   img_reg_array_45_10_imag;
  reg        [17:0]   img_reg_array_45_11_real;
  reg        [17:0]   img_reg_array_45_11_imag;
  reg        [17:0]   img_reg_array_45_12_real;
  reg        [17:0]   img_reg_array_45_12_imag;
  reg        [17:0]   img_reg_array_45_13_real;
  reg        [17:0]   img_reg_array_45_13_imag;
  reg        [17:0]   img_reg_array_45_14_real;
  reg        [17:0]   img_reg_array_45_14_imag;
  reg        [17:0]   img_reg_array_45_15_real;
  reg        [17:0]   img_reg_array_45_15_imag;
  reg        [17:0]   img_reg_array_45_16_real;
  reg        [17:0]   img_reg_array_45_16_imag;
  reg        [17:0]   img_reg_array_45_17_real;
  reg        [17:0]   img_reg_array_45_17_imag;
  reg        [17:0]   img_reg_array_45_18_real;
  reg        [17:0]   img_reg_array_45_18_imag;
  reg        [17:0]   img_reg_array_45_19_real;
  reg        [17:0]   img_reg_array_45_19_imag;
  reg        [17:0]   img_reg_array_45_20_real;
  reg        [17:0]   img_reg_array_45_20_imag;
  reg        [17:0]   img_reg_array_45_21_real;
  reg        [17:0]   img_reg_array_45_21_imag;
  reg        [17:0]   img_reg_array_45_22_real;
  reg        [17:0]   img_reg_array_45_22_imag;
  reg        [17:0]   img_reg_array_45_23_real;
  reg        [17:0]   img_reg_array_45_23_imag;
  reg        [17:0]   img_reg_array_45_24_real;
  reg        [17:0]   img_reg_array_45_24_imag;
  reg        [17:0]   img_reg_array_45_25_real;
  reg        [17:0]   img_reg_array_45_25_imag;
  reg        [17:0]   img_reg_array_45_26_real;
  reg        [17:0]   img_reg_array_45_26_imag;
  reg        [17:0]   img_reg_array_45_27_real;
  reg        [17:0]   img_reg_array_45_27_imag;
  reg        [17:0]   img_reg_array_45_28_real;
  reg        [17:0]   img_reg_array_45_28_imag;
  reg        [17:0]   img_reg_array_45_29_real;
  reg        [17:0]   img_reg_array_45_29_imag;
  reg        [17:0]   img_reg_array_45_30_real;
  reg        [17:0]   img_reg_array_45_30_imag;
  reg        [17:0]   img_reg_array_45_31_real;
  reg        [17:0]   img_reg_array_45_31_imag;
  reg        [17:0]   img_reg_array_45_32_real;
  reg        [17:0]   img_reg_array_45_32_imag;
  reg        [17:0]   img_reg_array_45_33_real;
  reg        [17:0]   img_reg_array_45_33_imag;
  reg        [17:0]   img_reg_array_45_34_real;
  reg        [17:0]   img_reg_array_45_34_imag;
  reg        [17:0]   img_reg_array_45_35_real;
  reg        [17:0]   img_reg_array_45_35_imag;
  reg        [17:0]   img_reg_array_45_36_real;
  reg        [17:0]   img_reg_array_45_36_imag;
  reg        [17:0]   img_reg_array_45_37_real;
  reg        [17:0]   img_reg_array_45_37_imag;
  reg        [17:0]   img_reg_array_45_38_real;
  reg        [17:0]   img_reg_array_45_38_imag;
  reg        [17:0]   img_reg_array_45_39_real;
  reg        [17:0]   img_reg_array_45_39_imag;
  reg        [17:0]   img_reg_array_45_40_real;
  reg        [17:0]   img_reg_array_45_40_imag;
  reg        [17:0]   img_reg_array_45_41_real;
  reg        [17:0]   img_reg_array_45_41_imag;
  reg        [17:0]   img_reg_array_45_42_real;
  reg        [17:0]   img_reg_array_45_42_imag;
  reg        [17:0]   img_reg_array_45_43_real;
  reg        [17:0]   img_reg_array_45_43_imag;
  reg        [17:0]   img_reg_array_45_44_real;
  reg        [17:0]   img_reg_array_45_44_imag;
  reg        [17:0]   img_reg_array_45_45_real;
  reg        [17:0]   img_reg_array_45_45_imag;
  reg        [17:0]   img_reg_array_45_46_real;
  reg        [17:0]   img_reg_array_45_46_imag;
  reg        [17:0]   img_reg_array_45_47_real;
  reg        [17:0]   img_reg_array_45_47_imag;
  reg        [17:0]   img_reg_array_45_48_real;
  reg        [17:0]   img_reg_array_45_48_imag;
  reg        [17:0]   img_reg_array_45_49_real;
  reg        [17:0]   img_reg_array_45_49_imag;
  reg        [17:0]   img_reg_array_45_50_real;
  reg        [17:0]   img_reg_array_45_50_imag;
  reg        [17:0]   img_reg_array_45_51_real;
  reg        [17:0]   img_reg_array_45_51_imag;
  reg        [17:0]   img_reg_array_45_52_real;
  reg        [17:0]   img_reg_array_45_52_imag;
  reg        [17:0]   img_reg_array_45_53_real;
  reg        [17:0]   img_reg_array_45_53_imag;
  reg        [17:0]   img_reg_array_45_54_real;
  reg        [17:0]   img_reg_array_45_54_imag;
  reg        [17:0]   img_reg_array_45_55_real;
  reg        [17:0]   img_reg_array_45_55_imag;
  reg        [17:0]   img_reg_array_45_56_real;
  reg        [17:0]   img_reg_array_45_56_imag;
  reg        [17:0]   img_reg_array_45_57_real;
  reg        [17:0]   img_reg_array_45_57_imag;
  reg        [17:0]   img_reg_array_45_58_real;
  reg        [17:0]   img_reg_array_45_58_imag;
  reg        [17:0]   img_reg_array_45_59_real;
  reg        [17:0]   img_reg_array_45_59_imag;
  reg        [17:0]   img_reg_array_45_60_real;
  reg        [17:0]   img_reg_array_45_60_imag;
  reg        [17:0]   img_reg_array_45_61_real;
  reg        [17:0]   img_reg_array_45_61_imag;
  reg        [17:0]   img_reg_array_45_62_real;
  reg        [17:0]   img_reg_array_45_62_imag;
  reg        [17:0]   img_reg_array_45_63_real;
  reg        [17:0]   img_reg_array_45_63_imag;
  reg        [17:0]   img_reg_array_46_0_real;
  reg        [17:0]   img_reg_array_46_0_imag;
  reg        [17:0]   img_reg_array_46_1_real;
  reg        [17:0]   img_reg_array_46_1_imag;
  reg        [17:0]   img_reg_array_46_2_real;
  reg        [17:0]   img_reg_array_46_2_imag;
  reg        [17:0]   img_reg_array_46_3_real;
  reg        [17:0]   img_reg_array_46_3_imag;
  reg        [17:0]   img_reg_array_46_4_real;
  reg        [17:0]   img_reg_array_46_4_imag;
  reg        [17:0]   img_reg_array_46_5_real;
  reg        [17:0]   img_reg_array_46_5_imag;
  reg        [17:0]   img_reg_array_46_6_real;
  reg        [17:0]   img_reg_array_46_6_imag;
  reg        [17:0]   img_reg_array_46_7_real;
  reg        [17:0]   img_reg_array_46_7_imag;
  reg        [17:0]   img_reg_array_46_8_real;
  reg        [17:0]   img_reg_array_46_8_imag;
  reg        [17:0]   img_reg_array_46_9_real;
  reg        [17:0]   img_reg_array_46_9_imag;
  reg        [17:0]   img_reg_array_46_10_real;
  reg        [17:0]   img_reg_array_46_10_imag;
  reg        [17:0]   img_reg_array_46_11_real;
  reg        [17:0]   img_reg_array_46_11_imag;
  reg        [17:0]   img_reg_array_46_12_real;
  reg        [17:0]   img_reg_array_46_12_imag;
  reg        [17:0]   img_reg_array_46_13_real;
  reg        [17:0]   img_reg_array_46_13_imag;
  reg        [17:0]   img_reg_array_46_14_real;
  reg        [17:0]   img_reg_array_46_14_imag;
  reg        [17:0]   img_reg_array_46_15_real;
  reg        [17:0]   img_reg_array_46_15_imag;
  reg        [17:0]   img_reg_array_46_16_real;
  reg        [17:0]   img_reg_array_46_16_imag;
  reg        [17:0]   img_reg_array_46_17_real;
  reg        [17:0]   img_reg_array_46_17_imag;
  reg        [17:0]   img_reg_array_46_18_real;
  reg        [17:0]   img_reg_array_46_18_imag;
  reg        [17:0]   img_reg_array_46_19_real;
  reg        [17:0]   img_reg_array_46_19_imag;
  reg        [17:0]   img_reg_array_46_20_real;
  reg        [17:0]   img_reg_array_46_20_imag;
  reg        [17:0]   img_reg_array_46_21_real;
  reg        [17:0]   img_reg_array_46_21_imag;
  reg        [17:0]   img_reg_array_46_22_real;
  reg        [17:0]   img_reg_array_46_22_imag;
  reg        [17:0]   img_reg_array_46_23_real;
  reg        [17:0]   img_reg_array_46_23_imag;
  reg        [17:0]   img_reg_array_46_24_real;
  reg        [17:0]   img_reg_array_46_24_imag;
  reg        [17:0]   img_reg_array_46_25_real;
  reg        [17:0]   img_reg_array_46_25_imag;
  reg        [17:0]   img_reg_array_46_26_real;
  reg        [17:0]   img_reg_array_46_26_imag;
  reg        [17:0]   img_reg_array_46_27_real;
  reg        [17:0]   img_reg_array_46_27_imag;
  reg        [17:0]   img_reg_array_46_28_real;
  reg        [17:0]   img_reg_array_46_28_imag;
  reg        [17:0]   img_reg_array_46_29_real;
  reg        [17:0]   img_reg_array_46_29_imag;
  reg        [17:0]   img_reg_array_46_30_real;
  reg        [17:0]   img_reg_array_46_30_imag;
  reg        [17:0]   img_reg_array_46_31_real;
  reg        [17:0]   img_reg_array_46_31_imag;
  reg        [17:0]   img_reg_array_46_32_real;
  reg        [17:0]   img_reg_array_46_32_imag;
  reg        [17:0]   img_reg_array_46_33_real;
  reg        [17:0]   img_reg_array_46_33_imag;
  reg        [17:0]   img_reg_array_46_34_real;
  reg        [17:0]   img_reg_array_46_34_imag;
  reg        [17:0]   img_reg_array_46_35_real;
  reg        [17:0]   img_reg_array_46_35_imag;
  reg        [17:0]   img_reg_array_46_36_real;
  reg        [17:0]   img_reg_array_46_36_imag;
  reg        [17:0]   img_reg_array_46_37_real;
  reg        [17:0]   img_reg_array_46_37_imag;
  reg        [17:0]   img_reg_array_46_38_real;
  reg        [17:0]   img_reg_array_46_38_imag;
  reg        [17:0]   img_reg_array_46_39_real;
  reg        [17:0]   img_reg_array_46_39_imag;
  reg        [17:0]   img_reg_array_46_40_real;
  reg        [17:0]   img_reg_array_46_40_imag;
  reg        [17:0]   img_reg_array_46_41_real;
  reg        [17:0]   img_reg_array_46_41_imag;
  reg        [17:0]   img_reg_array_46_42_real;
  reg        [17:0]   img_reg_array_46_42_imag;
  reg        [17:0]   img_reg_array_46_43_real;
  reg        [17:0]   img_reg_array_46_43_imag;
  reg        [17:0]   img_reg_array_46_44_real;
  reg        [17:0]   img_reg_array_46_44_imag;
  reg        [17:0]   img_reg_array_46_45_real;
  reg        [17:0]   img_reg_array_46_45_imag;
  reg        [17:0]   img_reg_array_46_46_real;
  reg        [17:0]   img_reg_array_46_46_imag;
  reg        [17:0]   img_reg_array_46_47_real;
  reg        [17:0]   img_reg_array_46_47_imag;
  reg        [17:0]   img_reg_array_46_48_real;
  reg        [17:0]   img_reg_array_46_48_imag;
  reg        [17:0]   img_reg_array_46_49_real;
  reg        [17:0]   img_reg_array_46_49_imag;
  reg        [17:0]   img_reg_array_46_50_real;
  reg        [17:0]   img_reg_array_46_50_imag;
  reg        [17:0]   img_reg_array_46_51_real;
  reg        [17:0]   img_reg_array_46_51_imag;
  reg        [17:0]   img_reg_array_46_52_real;
  reg        [17:0]   img_reg_array_46_52_imag;
  reg        [17:0]   img_reg_array_46_53_real;
  reg        [17:0]   img_reg_array_46_53_imag;
  reg        [17:0]   img_reg_array_46_54_real;
  reg        [17:0]   img_reg_array_46_54_imag;
  reg        [17:0]   img_reg_array_46_55_real;
  reg        [17:0]   img_reg_array_46_55_imag;
  reg        [17:0]   img_reg_array_46_56_real;
  reg        [17:0]   img_reg_array_46_56_imag;
  reg        [17:0]   img_reg_array_46_57_real;
  reg        [17:0]   img_reg_array_46_57_imag;
  reg        [17:0]   img_reg_array_46_58_real;
  reg        [17:0]   img_reg_array_46_58_imag;
  reg        [17:0]   img_reg_array_46_59_real;
  reg        [17:0]   img_reg_array_46_59_imag;
  reg        [17:0]   img_reg_array_46_60_real;
  reg        [17:0]   img_reg_array_46_60_imag;
  reg        [17:0]   img_reg_array_46_61_real;
  reg        [17:0]   img_reg_array_46_61_imag;
  reg        [17:0]   img_reg_array_46_62_real;
  reg        [17:0]   img_reg_array_46_62_imag;
  reg        [17:0]   img_reg_array_46_63_real;
  reg        [17:0]   img_reg_array_46_63_imag;
  reg        [17:0]   img_reg_array_47_0_real;
  reg        [17:0]   img_reg_array_47_0_imag;
  reg        [17:0]   img_reg_array_47_1_real;
  reg        [17:0]   img_reg_array_47_1_imag;
  reg        [17:0]   img_reg_array_47_2_real;
  reg        [17:0]   img_reg_array_47_2_imag;
  reg        [17:0]   img_reg_array_47_3_real;
  reg        [17:0]   img_reg_array_47_3_imag;
  reg        [17:0]   img_reg_array_47_4_real;
  reg        [17:0]   img_reg_array_47_4_imag;
  reg        [17:0]   img_reg_array_47_5_real;
  reg        [17:0]   img_reg_array_47_5_imag;
  reg        [17:0]   img_reg_array_47_6_real;
  reg        [17:0]   img_reg_array_47_6_imag;
  reg        [17:0]   img_reg_array_47_7_real;
  reg        [17:0]   img_reg_array_47_7_imag;
  reg        [17:0]   img_reg_array_47_8_real;
  reg        [17:0]   img_reg_array_47_8_imag;
  reg        [17:0]   img_reg_array_47_9_real;
  reg        [17:0]   img_reg_array_47_9_imag;
  reg        [17:0]   img_reg_array_47_10_real;
  reg        [17:0]   img_reg_array_47_10_imag;
  reg        [17:0]   img_reg_array_47_11_real;
  reg        [17:0]   img_reg_array_47_11_imag;
  reg        [17:0]   img_reg_array_47_12_real;
  reg        [17:0]   img_reg_array_47_12_imag;
  reg        [17:0]   img_reg_array_47_13_real;
  reg        [17:0]   img_reg_array_47_13_imag;
  reg        [17:0]   img_reg_array_47_14_real;
  reg        [17:0]   img_reg_array_47_14_imag;
  reg        [17:0]   img_reg_array_47_15_real;
  reg        [17:0]   img_reg_array_47_15_imag;
  reg        [17:0]   img_reg_array_47_16_real;
  reg        [17:0]   img_reg_array_47_16_imag;
  reg        [17:0]   img_reg_array_47_17_real;
  reg        [17:0]   img_reg_array_47_17_imag;
  reg        [17:0]   img_reg_array_47_18_real;
  reg        [17:0]   img_reg_array_47_18_imag;
  reg        [17:0]   img_reg_array_47_19_real;
  reg        [17:0]   img_reg_array_47_19_imag;
  reg        [17:0]   img_reg_array_47_20_real;
  reg        [17:0]   img_reg_array_47_20_imag;
  reg        [17:0]   img_reg_array_47_21_real;
  reg        [17:0]   img_reg_array_47_21_imag;
  reg        [17:0]   img_reg_array_47_22_real;
  reg        [17:0]   img_reg_array_47_22_imag;
  reg        [17:0]   img_reg_array_47_23_real;
  reg        [17:0]   img_reg_array_47_23_imag;
  reg        [17:0]   img_reg_array_47_24_real;
  reg        [17:0]   img_reg_array_47_24_imag;
  reg        [17:0]   img_reg_array_47_25_real;
  reg        [17:0]   img_reg_array_47_25_imag;
  reg        [17:0]   img_reg_array_47_26_real;
  reg        [17:0]   img_reg_array_47_26_imag;
  reg        [17:0]   img_reg_array_47_27_real;
  reg        [17:0]   img_reg_array_47_27_imag;
  reg        [17:0]   img_reg_array_47_28_real;
  reg        [17:0]   img_reg_array_47_28_imag;
  reg        [17:0]   img_reg_array_47_29_real;
  reg        [17:0]   img_reg_array_47_29_imag;
  reg        [17:0]   img_reg_array_47_30_real;
  reg        [17:0]   img_reg_array_47_30_imag;
  reg        [17:0]   img_reg_array_47_31_real;
  reg        [17:0]   img_reg_array_47_31_imag;
  reg        [17:0]   img_reg_array_47_32_real;
  reg        [17:0]   img_reg_array_47_32_imag;
  reg        [17:0]   img_reg_array_47_33_real;
  reg        [17:0]   img_reg_array_47_33_imag;
  reg        [17:0]   img_reg_array_47_34_real;
  reg        [17:0]   img_reg_array_47_34_imag;
  reg        [17:0]   img_reg_array_47_35_real;
  reg        [17:0]   img_reg_array_47_35_imag;
  reg        [17:0]   img_reg_array_47_36_real;
  reg        [17:0]   img_reg_array_47_36_imag;
  reg        [17:0]   img_reg_array_47_37_real;
  reg        [17:0]   img_reg_array_47_37_imag;
  reg        [17:0]   img_reg_array_47_38_real;
  reg        [17:0]   img_reg_array_47_38_imag;
  reg        [17:0]   img_reg_array_47_39_real;
  reg        [17:0]   img_reg_array_47_39_imag;
  reg        [17:0]   img_reg_array_47_40_real;
  reg        [17:0]   img_reg_array_47_40_imag;
  reg        [17:0]   img_reg_array_47_41_real;
  reg        [17:0]   img_reg_array_47_41_imag;
  reg        [17:0]   img_reg_array_47_42_real;
  reg        [17:0]   img_reg_array_47_42_imag;
  reg        [17:0]   img_reg_array_47_43_real;
  reg        [17:0]   img_reg_array_47_43_imag;
  reg        [17:0]   img_reg_array_47_44_real;
  reg        [17:0]   img_reg_array_47_44_imag;
  reg        [17:0]   img_reg_array_47_45_real;
  reg        [17:0]   img_reg_array_47_45_imag;
  reg        [17:0]   img_reg_array_47_46_real;
  reg        [17:0]   img_reg_array_47_46_imag;
  reg        [17:0]   img_reg_array_47_47_real;
  reg        [17:0]   img_reg_array_47_47_imag;
  reg        [17:0]   img_reg_array_47_48_real;
  reg        [17:0]   img_reg_array_47_48_imag;
  reg        [17:0]   img_reg_array_47_49_real;
  reg        [17:0]   img_reg_array_47_49_imag;
  reg        [17:0]   img_reg_array_47_50_real;
  reg        [17:0]   img_reg_array_47_50_imag;
  reg        [17:0]   img_reg_array_47_51_real;
  reg        [17:0]   img_reg_array_47_51_imag;
  reg        [17:0]   img_reg_array_47_52_real;
  reg        [17:0]   img_reg_array_47_52_imag;
  reg        [17:0]   img_reg_array_47_53_real;
  reg        [17:0]   img_reg_array_47_53_imag;
  reg        [17:0]   img_reg_array_47_54_real;
  reg        [17:0]   img_reg_array_47_54_imag;
  reg        [17:0]   img_reg_array_47_55_real;
  reg        [17:0]   img_reg_array_47_55_imag;
  reg        [17:0]   img_reg_array_47_56_real;
  reg        [17:0]   img_reg_array_47_56_imag;
  reg        [17:0]   img_reg_array_47_57_real;
  reg        [17:0]   img_reg_array_47_57_imag;
  reg        [17:0]   img_reg_array_47_58_real;
  reg        [17:0]   img_reg_array_47_58_imag;
  reg        [17:0]   img_reg_array_47_59_real;
  reg        [17:0]   img_reg_array_47_59_imag;
  reg        [17:0]   img_reg_array_47_60_real;
  reg        [17:0]   img_reg_array_47_60_imag;
  reg        [17:0]   img_reg_array_47_61_real;
  reg        [17:0]   img_reg_array_47_61_imag;
  reg        [17:0]   img_reg_array_47_62_real;
  reg        [17:0]   img_reg_array_47_62_imag;
  reg        [17:0]   img_reg_array_47_63_real;
  reg        [17:0]   img_reg_array_47_63_imag;
  reg        [17:0]   img_reg_array_48_0_real;
  reg        [17:0]   img_reg_array_48_0_imag;
  reg        [17:0]   img_reg_array_48_1_real;
  reg        [17:0]   img_reg_array_48_1_imag;
  reg        [17:0]   img_reg_array_48_2_real;
  reg        [17:0]   img_reg_array_48_2_imag;
  reg        [17:0]   img_reg_array_48_3_real;
  reg        [17:0]   img_reg_array_48_3_imag;
  reg        [17:0]   img_reg_array_48_4_real;
  reg        [17:0]   img_reg_array_48_4_imag;
  reg        [17:0]   img_reg_array_48_5_real;
  reg        [17:0]   img_reg_array_48_5_imag;
  reg        [17:0]   img_reg_array_48_6_real;
  reg        [17:0]   img_reg_array_48_6_imag;
  reg        [17:0]   img_reg_array_48_7_real;
  reg        [17:0]   img_reg_array_48_7_imag;
  reg        [17:0]   img_reg_array_48_8_real;
  reg        [17:0]   img_reg_array_48_8_imag;
  reg        [17:0]   img_reg_array_48_9_real;
  reg        [17:0]   img_reg_array_48_9_imag;
  reg        [17:0]   img_reg_array_48_10_real;
  reg        [17:0]   img_reg_array_48_10_imag;
  reg        [17:0]   img_reg_array_48_11_real;
  reg        [17:0]   img_reg_array_48_11_imag;
  reg        [17:0]   img_reg_array_48_12_real;
  reg        [17:0]   img_reg_array_48_12_imag;
  reg        [17:0]   img_reg_array_48_13_real;
  reg        [17:0]   img_reg_array_48_13_imag;
  reg        [17:0]   img_reg_array_48_14_real;
  reg        [17:0]   img_reg_array_48_14_imag;
  reg        [17:0]   img_reg_array_48_15_real;
  reg        [17:0]   img_reg_array_48_15_imag;
  reg        [17:0]   img_reg_array_48_16_real;
  reg        [17:0]   img_reg_array_48_16_imag;
  reg        [17:0]   img_reg_array_48_17_real;
  reg        [17:0]   img_reg_array_48_17_imag;
  reg        [17:0]   img_reg_array_48_18_real;
  reg        [17:0]   img_reg_array_48_18_imag;
  reg        [17:0]   img_reg_array_48_19_real;
  reg        [17:0]   img_reg_array_48_19_imag;
  reg        [17:0]   img_reg_array_48_20_real;
  reg        [17:0]   img_reg_array_48_20_imag;
  reg        [17:0]   img_reg_array_48_21_real;
  reg        [17:0]   img_reg_array_48_21_imag;
  reg        [17:0]   img_reg_array_48_22_real;
  reg        [17:0]   img_reg_array_48_22_imag;
  reg        [17:0]   img_reg_array_48_23_real;
  reg        [17:0]   img_reg_array_48_23_imag;
  reg        [17:0]   img_reg_array_48_24_real;
  reg        [17:0]   img_reg_array_48_24_imag;
  reg        [17:0]   img_reg_array_48_25_real;
  reg        [17:0]   img_reg_array_48_25_imag;
  reg        [17:0]   img_reg_array_48_26_real;
  reg        [17:0]   img_reg_array_48_26_imag;
  reg        [17:0]   img_reg_array_48_27_real;
  reg        [17:0]   img_reg_array_48_27_imag;
  reg        [17:0]   img_reg_array_48_28_real;
  reg        [17:0]   img_reg_array_48_28_imag;
  reg        [17:0]   img_reg_array_48_29_real;
  reg        [17:0]   img_reg_array_48_29_imag;
  reg        [17:0]   img_reg_array_48_30_real;
  reg        [17:0]   img_reg_array_48_30_imag;
  reg        [17:0]   img_reg_array_48_31_real;
  reg        [17:0]   img_reg_array_48_31_imag;
  reg        [17:0]   img_reg_array_48_32_real;
  reg        [17:0]   img_reg_array_48_32_imag;
  reg        [17:0]   img_reg_array_48_33_real;
  reg        [17:0]   img_reg_array_48_33_imag;
  reg        [17:0]   img_reg_array_48_34_real;
  reg        [17:0]   img_reg_array_48_34_imag;
  reg        [17:0]   img_reg_array_48_35_real;
  reg        [17:0]   img_reg_array_48_35_imag;
  reg        [17:0]   img_reg_array_48_36_real;
  reg        [17:0]   img_reg_array_48_36_imag;
  reg        [17:0]   img_reg_array_48_37_real;
  reg        [17:0]   img_reg_array_48_37_imag;
  reg        [17:0]   img_reg_array_48_38_real;
  reg        [17:0]   img_reg_array_48_38_imag;
  reg        [17:0]   img_reg_array_48_39_real;
  reg        [17:0]   img_reg_array_48_39_imag;
  reg        [17:0]   img_reg_array_48_40_real;
  reg        [17:0]   img_reg_array_48_40_imag;
  reg        [17:0]   img_reg_array_48_41_real;
  reg        [17:0]   img_reg_array_48_41_imag;
  reg        [17:0]   img_reg_array_48_42_real;
  reg        [17:0]   img_reg_array_48_42_imag;
  reg        [17:0]   img_reg_array_48_43_real;
  reg        [17:0]   img_reg_array_48_43_imag;
  reg        [17:0]   img_reg_array_48_44_real;
  reg        [17:0]   img_reg_array_48_44_imag;
  reg        [17:0]   img_reg_array_48_45_real;
  reg        [17:0]   img_reg_array_48_45_imag;
  reg        [17:0]   img_reg_array_48_46_real;
  reg        [17:0]   img_reg_array_48_46_imag;
  reg        [17:0]   img_reg_array_48_47_real;
  reg        [17:0]   img_reg_array_48_47_imag;
  reg        [17:0]   img_reg_array_48_48_real;
  reg        [17:0]   img_reg_array_48_48_imag;
  reg        [17:0]   img_reg_array_48_49_real;
  reg        [17:0]   img_reg_array_48_49_imag;
  reg        [17:0]   img_reg_array_48_50_real;
  reg        [17:0]   img_reg_array_48_50_imag;
  reg        [17:0]   img_reg_array_48_51_real;
  reg        [17:0]   img_reg_array_48_51_imag;
  reg        [17:0]   img_reg_array_48_52_real;
  reg        [17:0]   img_reg_array_48_52_imag;
  reg        [17:0]   img_reg_array_48_53_real;
  reg        [17:0]   img_reg_array_48_53_imag;
  reg        [17:0]   img_reg_array_48_54_real;
  reg        [17:0]   img_reg_array_48_54_imag;
  reg        [17:0]   img_reg_array_48_55_real;
  reg        [17:0]   img_reg_array_48_55_imag;
  reg        [17:0]   img_reg_array_48_56_real;
  reg        [17:0]   img_reg_array_48_56_imag;
  reg        [17:0]   img_reg_array_48_57_real;
  reg        [17:0]   img_reg_array_48_57_imag;
  reg        [17:0]   img_reg_array_48_58_real;
  reg        [17:0]   img_reg_array_48_58_imag;
  reg        [17:0]   img_reg_array_48_59_real;
  reg        [17:0]   img_reg_array_48_59_imag;
  reg        [17:0]   img_reg_array_48_60_real;
  reg        [17:0]   img_reg_array_48_60_imag;
  reg        [17:0]   img_reg_array_48_61_real;
  reg        [17:0]   img_reg_array_48_61_imag;
  reg        [17:0]   img_reg_array_48_62_real;
  reg        [17:0]   img_reg_array_48_62_imag;
  reg        [17:0]   img_reg_array_48_63_real;
  reg        [17:0]   img_reg_array_48_63_imag;
  reg        [17:0]   img_reg_array_49_0_real;
  reg        [17:0]   img_reg_array_49_0_imag;
  reg        [17:0]   img_reg_array_49_1_real;
  reg        [17:0]   img_reg_array_49_1_imag;
  reg        [17:0]   img_reg_array_49_2_real;
  reg        [17:0]   img_reg_array_49_2_imag;
  reg        [17:0]   img_reg_array_49_3_real;
  reg        [17:0]   img_reg_array_49_3_imag;
  reg        [17:0]   img_reg_array_49_4_real;
  reg        [17:0]   img_reg_array_49_4_imag;
  reg        [17:0]   img_reg_array_49_5_real;
  reg        [17:0]   img_reg_array_49_5_imag;
  reg        [17:0]   img_reg_array_49_6_real;
  reg        [17:0]   img_reg_array_49_6_imag;
  reg        [17:0]   img_reg_array_49_7_real;
  reg        [17:0]   img_reg_array_49_7_imag;
  reg        [17:0]   img_reg_array_49_8_real;
  reg        [17:0]   img_reg_array_49_8_imag;
  reg        [17:0]   img_reg_array_49_9_real;
  reg        [17:0]   img_reg_array_49_9_imag;
  reg        [17:0]   img_reg_array_49_10_real;
  reg        [17:0]   img_reg_array_49_10_imag;
  reg        [17:0]   img_reg_array_49_11_real;
  reg        [17:0]   img_reg_array_49_11_imag;
  reg        [17:0]   img_reg_array_49_12_real;
  reg        [17:0]   img_reg_array_49_12_imag;
  reg        [17:0]   img_reg_array_49_13_real;
  reg        [17:0]   img_reg_array_49_13_imag;
  reg        [17:0]   img_reg_array_49_14_real;
  reg        [17:0]   img_reg_array_49_14_imag;
  reg        [17:0]   img_reg_array_49_15_real;
  reg        [17:0]   img_reg_array_49_15_imag;
  reg        [17:0]   img_reg_array_49_16_real;
  reg        [17:0]   img_reg_array_49_16_imag;
  reg        [17:0]   img_reg_array_49_17_real;
  reg        [17:0]   img_reg_array_49_17_imag;
  reg        [17:0]   img_reg_array_49_18_real;
  reg        [17:0]   img_reg_array_49_18_imag;
  reg        [17:0]   img_reg_array_49_19_real;
  reg        [17:0]   img_reg_array_49_19_imag;
  reg        [17:0]   img_reg_array_49_20_real;
  reg        [17:0]   img_reg_array_49_20_imag;
  reg        [17:0]   img_reg_array_49_21_real;
  reg        [17:0]   img_reg_array_49_21_imag;
  reg        [17:0]   img_reg_array_49_22_real;
  reg        [17:0]   img_reg_array_49_22_imag;
  reg        [17:0]   img_reg_array_49_23_real;
  reg        [17:0]   img_reg_array_49_23_imag;
  reg        [17:0]   img_reg_array_49_24_real;
  reg        [17:0]   img_reg_array_49_24_imag;
  reg        [17:0]   img_reg_array_49_25_real;
  reg        [17:0]   img_reg_array_49_25_imag;
  reg        [17:0]   img_reg_array_49_26_real;
  reg        [17:0]   img_reg_array_49_26_imag;
  reg        [17:0]   img_reg_array_49_27_real;
  reg        [17:0]   img_reg_array_49_27_imag;
  reg        [17:0]   img_reg_array_49_28_real;
  reg        [17:0]   img_reg_array_49_28_imag;
  reg        [17:0]   img_reg_array_49_29_real;
  reg        [17:0]   img_reg_array_49_29_imag;
  reg        [17:0]   img_reg_array_49_30_real;
  reg        [17:0]   img_reg_array_49_30_imag;
  reg        [17:0]   img_reg_array_49_31_real;
  reg        [17:0]   img_reg_array_49_31_imag;
  reg        [17:0]   img_reg_array_49_32_real;
  reg        [17:0]   img_reg_array_49_32_imag;
  reg        [17:0]   img_reg_array_49_33_real;
  reg        [17:0]   img_reg_array_49_33_imag;
  reg        [17:0]   img_reg_array_49_34_real;
  reg        [17:0]   img_reg_array_49_34_imag;
  reg        [17:0]   img_reg_array_49_35_real;
  reg        [17:0]   img_reg_array_49_35_imag;
  reg        [17:0]   img_reg_array_49_36_real;
  reg        [17:0]   img_reg_array_49_36_imag;
  reg        [17:0]   img_reg_array_49_37_real;
  reg        [17:0]   img_reg_array_49_37_imag;
  reg        [17:0]   img_reg_array_49_38_real;
  reg        [17:0]   img_reg_array_49_38_imag;
  reg        [17:0]   img_reg_array_49_39_real;
  reg        [17:0]   img_reg_array_49_39_imag;
  reg        [17:0]   img_reg_array_49_40_real;
  reg        [17:0]   img_reg_array_49_40_imag;
  reg        [17:0]   img_reg_array_49_41_real;
  reg        [17:0]   img_reg_array_49_41_imag;
  reg        [17:0]   img_reg_array_49_42_real;
  reg        [17:0]   img_reg_array_49_42_imag;
  reg        [17:0]   img_reg_array_49_43_real;
  reg        [17:0]   img_reg_array_49_43_imag;
  reg        [17:0]   img_reg_array_49_44_real;
  reg        [17:0]   img_reg_array_49_44_imag;
  reg        [17:0]   img_reg_array_49_45_real;
  reg        [17:0]   img_reg_array_49_45_imag;
  reg        [17:0]   img_reg_array_49_46_real;
  reg        [17:0]   img_reg_array_49_46_imag;
  reg        [17:0]   img_reg_array_49_47_real;
  reg        [17:0]   img_reg_array_49_47_imag;
  reg        [17:0]   img_reg_array_49_48_real;
  reg        [17:0]   img_reg_array_49_48_imag;
  reg        [17:0]   img_reg_array_49_49_real;
  reg        [17:0]   img_reg_array_49_49_imag;
  reg        [17:0]   img_reg_array_49_50_real;
  reg        [17:0]   img_reg_array_49_50_imag;
  reg        [17:0]   img_reg_array_49_51_real;
  reg        [17:0]   img_reg_array_49_51_imag;
  reg        [17:0]   img_reg_array_49_52_real;
  reg        [17:0]   img_reg_array_49_52_imag;
  reg        [17:0]   img_reg_array_49_53_real;
  reg        [17:0]   img_reg_array_49_53_imag;
  reg        [17:0]   img_reg_array_49_54_real;
  reg        [17:0]   img_reg_array_49_54_imag;
  reg        [17:0]   img_reg_array_49_55_real;
  reg        [17:0]   img_reg_array_49_55_imag;
  reg        [17:0]   img_reg_array_49_56_real;
  reg        [17:0]   img_reg_array_49_56_imag;
  reg        [17:0]   img_reg_array_49_57_real;
  reg        [17:0]   img_reg_array_49_57_imag;
  reg        [17:0]   img_reg_array_49_58_real;
  reg        [17:0]   img_reg_array_49_58_imag;
  reg        [17:0]   img_reg_array_49_59_real;
  reg        [17:0]   img_reg_array_49_59_imag;
  reg        [17:0]   img_reg_array_49_60_real;
  reg        [17:0]   img_reg_array_49_60_imag;
  reg        [17:0]   img_reg_array_49_61_real;
  reg        [17:0]   img_reg_array_49_61_imag;
  reg        [17:0]   img_reg_array_49_62_real;
  reg        [17:0]   img_reg_array_49_62_imag;
  reg        [17:0]   img_reg_array_49_63_real;
  reg        [17:0]   img_reg_array_49_63_imag;
  reg        [17:0]   img_reg_array_50_0_real;
  reg        [17:0]   img_reg_array_50_0_imag;
  reg        [17:0]   img_reg_array_50_1_real;
  reg        [17:0]   img_reg_array_50_1_imag;
  reg        [17:0]   img_reg_array_50_2_real;
  reg        [17:0]   img_reg_array_50_2_imag;
  reg        [17:0]   img_reg_array_50_3_real;
  reg        [17:0]   img_reg_array_50_3_imag;
  reg        [17:0]   img_reg_array_50_4_real;
  reg        [17:0]   img_reg_array_50_4_imag;
  reg        [17:0]   img_reg_array_50_5_real;
  reg        [17:0]   img_reg_array_50_5_imag;
  reg        [17:0]   img_reg_array_50_6_real;
  reg        [17:0]   img_reg_array_50_6_imag;
  reg        [17:0]   img_reg_array_50_7_real;
  reg        [17:0]   img_reg_array_50_7_imag;
  reg        [17:0]   img_reg_array_50_8_real;
  reg        [17:0]   img_reg_array_50_8_imag;
  reg        [17:0]   img_reg_array_50_9_real;
  reg        [17:0]   img_reg_array_50_9_imag;
  reg        [17:0]   img_reg_array_50_10_real;
  reg        [17:0]   img_reg_array_50_10_imag;
  reg        [17:0]   img_reg_array_50_11_real;
  reg        [17:0]   img_reg_array_50_11_imag;
  reg        [17:0]   img_reg_array_50_12_real;
  reg        [17:0]   img_reg_array_50_12_imag;
  reg        [17:0]   img_reg_array_50_13_real;
  reg        [17:0]   img_reg_array_50_13_imag;
  reg        [17:0]   img_reg_array_50_14_real;
  reg        [17:0]   img_reg_array_50_14_imag;
  reg        [17:0]   img_reg_array_50_15_real;
  reg        [17:0]   img_reg_array_50_15_imag;
  reg        [17:0]   img_reg_array_50_16_real;
  reg        [17:0]   img_reg_array_50_16_imag;
  reg        [17:0]   img_reg_array_50_17_real;
  reg        [17:0]   img_reg_array_50_17_imag;
  reg        [17:0]   img_reg_array_50_18_real;
  reg        [17:0]   img_reg_array_50_18_imag;
  reg        [17:0]   img_reg_array_50_19_real;
  reg        [17:0]   img_reg_array_50_19_imag;
  reg        [17:0]   img_reg_array_50_20_real;
  reg        [17:0]   img_reg_array_50_20_imag;
  reg        [17:0]   img_reg_array_50_21_real;
  reg        [17:0]   img_reg_array_50_21_imag;
  reg        [17:0]   img_reg_array_50_22_real;
  reg        [17:0]   img_reg_array_50_22_imag;
  reg        [17:0]   img_reg_array_50_23_real;
  reg        [17:0]   img_reg_array_50_23_imag;
  reg        [17:0]   img_reg_array_50_24_real;
  reg        [17:0]   img_reg_array_50_24_imag;
  reg        [17:0]   img_reg_array_50_25_real;
  reg        [17:0]   img_reg_array_50_25_imag;
  reg        [17:0]   img_reg_array_50_26_real;
  reg        [17:0]   img_reg_array_50_26_imag;
  reg        [17:0]   img_reg_array_50_27_real;
  reg        [17:0]   img_reg_array_50_27_imag;
  reg        [17:0]   img_reg_array_50_28_real;
  reg        [17:0]   img_reg_array_50_28_imag;
  reg        [17:0]   img_reg_array_50_29_real;
  reg        [17:0]   img_reg_array_50_29_imag;
  reg        [17:0]   img_reg_array_50_30_real;
  reg        [17:0]   img_reg_array_50_30_imag;
  reg        [17:0]   img_reg_array_50_31_real;
  reg        [17:0]   img_reg_array_50_31_imag;
  reg        [17:0]   img_reg_array_50_32_real;
  reg        [17:0]   img_reg_array_50_32_imag;
  reg        [17:0]   img_reg_array_50_33_real;
  reg        [17:0]   img_reg_array_50_33_imag;
  reg        [17:0]   img_reg_array_50_34_real;
  reg        [17:0]   img_reg_array_50_34_imag;
  reg        [17:0]   img_reg_array_50_35_real;
  reg        [17:0]   img_reg_array_50_35_imag;
  reg        [17:0]   img_reg_array_50_36_real;
  reg        [17:0]   img_reg_array_50_36_imag;
  reg        [17:0]   img_reg_array_50_37_real;
  reg        [17:0]   img_reg_array_50_37_imag;
  reg        [17:0]   img_reg_array_50_38_real;
  reg        [17:0]   img_reg_array_50_38_imag;
  reg        [17:0]   img_reg_array_50_39_real;
  reg        [17:0]   img_reg_array_50_39_imag;
  reg        [17:0]   img_reg_array_50_40_real;
  reg        [17:0]   img_reg_array_50_40_imag;
  reg        [17:0]   img_reg_array_50_41_real;
  reg        [17:0]   img_reg_array_50_41_imag;
  reg        [17:0]   img_reg_array_50_42_real;
  reg        [17:0]   img_reg_array_50_42_imag;
  reg        [17:0]   img_reg_array_50_43_real;
  reg        [17:0]   img_reg_array_50_43_imag;
  reg        [17:0]   img_reg_array_50_44_real;
  reg        [17:0]   img_reg_array_50_44_imag;
  reg        [17:0]   img_reg_array_50_45_real;
  reg        [17:0]   img_reg_array_50_45_imag;
  reg        [17:0]   img_reg_array_50_46_real;
  reg        [17:0]   img_reg_array_50_46_imag;
  reg        [17:0]   img_reg_array_50_47_real;
  reg        [17:0]   img_reg_array_50_47_imag;
  reg        [17:0]   img_reg_array_50_48_real;
  reg        [17:0]   img_reg_array_50_48_imag;
  reg        [17:0]   img_reg_array_50_49_real;
  reg        [17:0]   img_reg_array_50_49_imag;
  reg        [17:0]   img_reg_array_50_50_real;
  reg        [17:0]   img_reg_array_50_50_imag;
  reg        [17:0]   img_reg_array_50_51_real;
  reg        [17:0]   img_reg_array_50_51_imag;
  reg        [17:0]   img_reg_array_50_52_real;
  reg        [17:0]   img_reg_array_50_52_imag;
  reg        [17:0]   img_reg_array_50_53_real;
  reg        [17:0]   img_reg_array_50_53_imag;
  reg        [17:0]   img_reg_array_50_54_real;
  reg        [17:0]   img_reg_array_50_54_imag;
  reg        [17:0]   img_reg_array_50_55_real;
  reg        [17:0]   img_reg_array_50_55_imag;
  reg        [17:0]   img_reg_array_50_56_real;
  reg        [17:0]   img_reg_array_50_56_imag;
  reg        [17:0]   img_reg_array_50_57_real;
  reg        [17:0]   img_reg_array_50_57_imag;
  reg        [17:0]   img_reg_array_50_58_real;
  reg        [17:0]   img_reg_array_50_58_imag;
  reg        [17:0]   img_reg_array_50_59_real;
  reg        [17:0]   img_reg_array_50_59_imag;
  reg        [17:0]   img_reg_array_50_60_real;
  reg        [17:0]   img_reg_array_50_60_imag;
  reg        [17:0]   img_reg_array_50_61_real;
  reg        [17:0]   img_reg_array_50_61_imag;
  reg        [17:0]   img_reg_array_50_62_real;
  reg        [17:0]   img_reg_array_50_62_imag;
  reg        [17:0]   img_reg_array_50_63_real;
  reg        [17:0]   img_reg_array_50_63_imag;
  reg        [17:0]   img_reg_array_51_0_real;
  reg        [17:0]   img_reg_array_51_0_imag;
  reg        [17:0]   img_reg_array_51_1_real;
  reg        [17:0]   img_reg_array_51_1_imag;
  reg        [17:0]   img_reg_array_51_2_real;
  reg        [17:0]   img_reg_array_51_2_imag;
  reg        [17:0]   img_reg_array_51_3_real;
  reg        [17:0]   img_reg_array_51_3_imag;
  reg        [17:0]   img_reg_array_51_4_real;
  reg        [17:0]   img_reg_array_51_4_imag;
  reg        [17:0]   img_reg_array_51_5_real;
  reg        [17:0]   img_reg_array_51_5_imag;
  reg        [17:0]   img_reg_array_51_6_real;
  reg        [17:0]   img_reg_array_51_6_imag;
  reg        [17:0]   img_reg_array_51_7_real;
  reg        [17:0]   img_reg_array_51_7_imag;
  reg        [17:0]   img_reg_array_51_8_real;
  reg        [17:0]   img_reg_array_51_8_imag;
  reg        [17:0]   img_reg_array_51_9_real;
  reg        [17:0]   img_reg_array_51_9_imag;
  reg        [17:0]   img_reg_array_51_10_real;
  reg        [17:0]   img_reg_array_51_10_imag;
  reg        [17:0]   img_reg_array_51_11_real;
  reg        [17:0]   img_reg_array_51_11_imag;
  reg        [17:0]   img_reg_array_51_12_real;
  reg        [17:0]   img_reg_array_51_12_imag;
  reg        [17:0]   img_reg_array_51_13_real;
  reg        [17:0]   img_reg_array_51_13_imag;
  reg        [17:0]   img_reg_array_51_14_real;
  reg        [17:0]   img_reg_array_51_14_imag;
  reg        [17:0]   img_reg_array_51_15_real;
  reg        [17:0]   img_reg_array_51_15_imag;
  reg        [17:0]   img_reg_array_51_16_real;
  reg        [17:0]   img_reg_array_51_16_imag;
  reg        [17:0]   img_reg_array_51_17_real;
  reg        [17:0]   img_reg_array_51_17_imag;
  reg        [17:0]   img_reg_array_51_18_real;
  reg        [17:0]   img_reg_array_51_18_imag;
  reg        [17:0]   img_reg_array_51_19_real;
  reg        [17:0]   img_reg_array_51_19_imag;
  reg        [17:0]   img_reg_array_51_20_real;
  reg        [17:0]   img_reg_array_51_20_imag;
  reg        [17:0]   img_reg_array_51_21_real;
  reg        [17:0]   img_reg_array_51_21_imag;
  reg        [17:0]   img_reg_array_51_22_real;
  reg        [17:0]   img_reg_array_51_22_imag;
  reg        [17:0]   img_reg_array_51_23_real;
  reg        [17:0]   img_reg_array_51_23_imag;
  reg        [17:0]   img_reg_array_51_24_real;
  reg        [17:0]   img_reg_array_51_24_imag;
  reg        [17:0]   img_reg_array_51_25_real;
  reg        [17:0]   img_reg_array_51_25_imag;
  reg        [17:0]   img_reg_array_51_26_real;
  reg        [17:0]   img_reg_array_51_26_imag;
  reg        [17:0]   img_reg_array_51_27_real;
  reg        [17:0]   img_reg_array_51_27_imag;
  reg        [17:0]   img_reg_array_51_28_real;
  reg        [17:0]   img_reg_array_51_28_imag;
  reg        [17:0]   img_reg_array_51_29_real;
  reg        [17:0]   img_reg_array_51_29_imag;
  reg        [17:0]   img_reg_array_51_30_real;
  reg        [17:0]   img_reg_array_51_30_imag;
  reg        [17:0]   img_reg_array_51_31_real;
  reg        [17:0]   img_reg_array_51_31_imag;
  reg        [17:0]   img_reg_array_51_32_real;
  reg        [17:0]   img_reg_array_51_32_imag;
  reg        [17:0]   img_reg_array_51_33_real;
  reg        [17:0]   img_reg_array_51_33_imag;
  reg        [17:0]   img_reg_array_51_34_real;
  reg        [17:0]   img_reg_array_51_34_imag;
  reg        [17:0]   img_reg_array_51_35_real;
  reg        [17:0]   img_reg_array_51_35_imag;
  reg        [17:0]   img_reg_array_51_36_real;
  reg        [17:0]   img_reg_array_51_36_imag;
  reg        [17:0]   img_reg_array_51_37_real;
  reg        [17:0]   img_reg_array_51_37_imag;
  reg        [17:0]   img_reg_array_51_38_real;
  reg        [17:0]   img_reg_array_51_38_imag;
  reg        [17:0]   img_reg_array_51_39_real;
  reg        [17:0]   img_reg_array_51_39_imag;
  reg        [17:0]   img_reg_array_51_40_real;
  reg        [17:0]   img_reg_array_51_40_imag;
  reg        [17:0]   img_reg_array_51_41_real;
  reg        [17:0]   img_reg_array_51_41_imag;
  reg        [17:0]   img_reg_array_51_42_real;
  reg        [17:0]   img_reg_array_51_42_imag;
  reg        [17:0]   img_reg_array_51_43_real;
  reg        [17:0]   img_reg_array_51_43_imag;
  reg        [17:0]   img_reg_array_51_44_real;
  reg        [17:0]   img_reg_array_51_44_imag;
  reg        [17:0]   img_reg_array_51_45_real;
  reg        [17:0]   img_reg_array_51_45_imag;
  reg        [17:0]   img_reg_array_51_46_real;
  reg        [17:0]   img_reg_array_51_46_imag;
  reg        [17:0]   img_reg_array_51_47_real;
  reg        [17:0]   img_reg_array_51_47_imag;
  reg        [17:0]   img_reg_array_51_48_real;
  reg        [17:0]   img_reg_array_51_48_imag;
  reg        [17:0]   img_reg_array_51_49_real;
  reg        [17:0]   img_reg_array_51_49_imag;
  reg        [17:0]   img_reg_array_51_50_real;
  reg        [17:0]   img_reg_array_51_50_imag;
  reg        [17:0]   img_reg_array_51_51_real;
  reg        [17:0]   img_reg_array_51_51_imag;
  reg        [17:0]   img_reg_array_51_52_real;
  reg        [17:0]   img_reg_array_51_52_imag;
  reg        [17:0]   img_reg_array_51_53_real;
  reg        [17:0]   img_reg_array_51_53_imag;
  reg        [17:0]   img_reg_array_51_54_real;
  reg        [17:0]   img_reg_array_51_54_imag;
  reg        [17:0]   img_reg_array_51_55_real;
  reg        [17:0]   img_reg_array_51_55_imag;
  reg        [17:0]   img_reg_array_51_56_real;
  reg        [17:0]   img_reg_array_51_56_imag;
  reg        [17:0]   img_reg_array_51_57_real;
  reg        [17:0]   img_reg_array_51_57_imag;
  reg        [17:0]   img_reg_array_51_58_real;
  reg        [17:0]   img_reg_array_51_58_imag;
  reg        [17:0]   img_reg_array_51_59_real;
  reg        [17:0]   img_reg_array_51_59_imag;
  reg        [17:0]   img_reg_array_51_60_real;
  reg        [17:0]   img_reg_array_51_60_imag;
  reg        [17:0]   img_reg_array_51_61_real;
  reg        [17:0]   img_reg_array_51_61_imag;
  reg        [17:0]   img_reg_array_51_62_real;
  reg        [17:0]   img_reg_array_51_62_imag;
  reg        [17:0]   img_reg_array_51_63_real;
  reg        [17:0]   img_reg_array_51_63_imag;
  reg        [17:0]   img_reg_array_52_0_real;
  reg        [17:0]   img_reg_array_52_0_imag;
  reg        [17:0]   img_reg_array_52_1_real;
  reg        [17:0]   img_reg_array_52_1_imag;
  reg        [17:0]   img_reg_array_52_2_real;
  reg        [17:0]   img_reg_array_52_2_imag;
  reg        [17:0]   img_reg_array_52_3_real;
  reg        [17:0]   img_reg_array_52_3_imag;
  reg        [17:0]   img_reg_array_52_4_real;
  reg        [17:0]   img_reg_array_52_4_imag;
  reg        [17:0]   img_reg_array_52_5_real;
  reg        [17:0]   img_reg_array_52_5_imag;
  reg        [17:0]   img_reg_array_52_6_real;
  reg        [17:0]   img_reg_array_52_6_imag;
  reg        [17:0]   img_reg_array_52_7_real;
  reg        [17:0]   img_reg_array_52_7_imag;
  reg        [17:0]   img_reg_array_52_8_real;
  reg        [17:0]   img_reg_array_52_8_imag;
  reg        [17:0]   img_reg_array_52_9_real;
  reg        [17:0]   img_reg_array_52_9_imag;
  reg        [17:0]   img_reg_array_52_10_real;
  reg        [17:0]   img_reg_array_52_10_imag;
  reg        [17:0]   img_reg_array_52_11_real;
  reg        [17:0]   img_reg_array_52_11_imag;
  reg        [17:0]   img_reg_array_52_12_real;
  reg        [17:0]   img_reg_array_52_12_imag;
  reg        [17:0]   img_reg_array_52_13_real;
  reg        [17:0]   img_reg_array_52_13_imag;
  reg        [17:0]   img_reg_array_52_14_real;
  reg        [17:0]   img_reg_array_52_14_imag;
  reg        [17:0]   img_reg_array_52_15_real;
  reg        [17:0]   img_reg_array_52_15_imag;
  reg        [17:0]   img_reg_array_52_16_real;
  reg        [17:0]   img_reg_array_52_16_imag;
  reg        [17:0]   img_reg_array_52_17_real;
  reg        [17:0]   img_reg_array_52_17_imag;
  reg        [17:0]   img_reg_array_52_18_real;
  reg        [17:0]   img_reg_array_52_18_imag;
  reg        [17:0]   img_reg_array_52_19_real;
  reg        [17:0]   img_reg_array_52_19_imag;
  reg        [17:0]   img_reg_array_52_20_real;
  reg        [17:0]   img_reg_array_52_20_imag;
  reg        [17:0]   img_reg_array_52_21_real;
  reg        [17:0]   img_reg_array_52_21_imag;
  reg        [17:0]   img_reg_array_52_22_real;
  reg        [17:0]   img_reg_array_52_22_imag;
  reg        [17:0]   img_reg_array_52_23_real;
  reg        [17:0]   img_reg_array_52_23_imag;
  reg        [17:0]   img_reg_array_52_24_real;
  reg        [17:0]   img_reg_array_52_24_imag;
  reg        [17:0]   img_reg_array_52_25_real;
  reg        [17:0]   img_reg_array_52_25_imag;
  reg        [17:0]   img_reg_array_52_26_real;
  reg        [17:0]   img_reg_array_52_26_imag;
  reg        [17:0]   img_reg_array_52_27_real;
  reg        [17:0]   img_reg_array_52_27_imag;
  reg        [17:0]   img_reg_array_52_28_real;
  reg        [17:0]   img_reg_array_52_28_imag;
  reg        [17:0]   img_reg_array_52_29_real;
  reg        [17:0]   img_reg_array_52_29_imag;
  reg        [17:0]   img_reg_array_52_30_real;
  reg        [17:0]   img_reg_array_52_30_imag;
  reg        [17:0]   img_reg_array_52_31_real;
  reg        [17:0]   img_reg_array_52_31_imag;
  reg        [17:0]   img_reg_array_52_32_real;
  reg        [17:0]   img_reg_array_52_32_imag;
  reg        [17:0]   img_reg_array_52_33_real;
  reg        [17:0]   img_reg_array_52_33_imag;
  reg        [17:0]   img_reg_array_52_34_real;
  reg        [17:0]   img_reg_array_52_34_imag;
  reg        [17:0]   img_reg_array_52_35_real;
  reg        [17:0]   img_reg_array_52_35_imag;
  reg        [17:0]   img_reg_array_52_36_real;
  reg        [17:0]   img_reg_array_52_36_imag;
  reg        [17:0]   img_reg_array_52_37_real;
  reg        [17:0]   img_reg_array_52_37_imag;
  reg        [17:0]   img_reg_array_52_38_real;
  reg        [17:0]   img_reg_array_52_38_imag;
  reg        [17:0]   img_reg_array_52_39_real;
  reg        [17:0]   img_reg_array_52_39_imag;
  reg        [17:0]   img_reg_array_52_40_real;
  reg        [17:0]   img_reg_array_52_40_imag;
  reg        [17:0]   img_reg_array_52_41_real;
  reg        [17:0]   img_reg_array_52_41_imag;
  reg        [17:0]   img_reg_array_52_42_real;
  reg        [17:0]   img_reg_array_52_42_imag;
  reg        [17:0]   img_reg_array_52_43_real;
  reg        [17:0]   img_reg_array_52_43_imag;
  reg        [17:0]   img_reg_array_52_44_real;
  reg        [17:0]   img_reg_array_52_44_imag;
  reg        [17:0]   img_reg_array_52_45_real;
  reg        [17:0]   img_reg_array_52_45_imag;
  reg        [17:0]   img_reg_array_52_46_real;
  reg        [17:0]   img_reg_array_52_46_imag;
  reg        [17:0]   img_reg_array_52_47_real;
  reg        [17:0]   img_reg_array_52_47_imag;
  reg        [17:0]   img_reg_array_52_48_real;
  reg        [17:0]   img_reg_array_52_48_imag;
  reg        [17:0]   img_reg_array_52_49_real;
  reg        [17:0]   img_reg_array_52_49_imag;
  reg        [17:0]   img_reg_array_52_50_real;
  reg        [17:0]   img_reg_array_52_50_imag;
  reg        [17:0]   img_reg_array_52_51_real;
  reg        [17:0]   img_reg_array_52_51_imag;
  reg        [17:0]   img_reg_array_52_52_real;
  reg        [17:0]   img_reg_array_52_52_imag;
  reg        [17:0]   img_reg_array_52_53_real;
  reg        [17:0]   img_reg_array_52_53_imag;
  reg        [17:0]   img_reg_array_52_54_real;
  reg        [17:0]   img_reg_array_52_54_imag;
  reg        [17:0]   img_reg_array_52_55_real;
  reg        [17:0]   img_reg_array_52_55_imag;
  reg        [17:0]   img_reg_array_52_56_real;
  reg        [17:0]   img_reg_array_52_56_imag;
  reg        [17:0]   img_reg_array_52_57_real;
  reg        [17:0]   img_reg_array_52_57_imag;
  reg        [17:0]   img_reg_array_52_58_real;
  reg        [17:0]   img_reg_array_52_58_imag;
  reg        [17:0]   img_reg_array_52_59_real;
  reg        [17:0]   img_reg_array_52_59_imag;
  reg        [17:0]   img_reg_array_52_60_real;
  reg        [17:0]   img_reg_array_52_60_imag;
  reg        [17:0]   img_reg_array_52_61_real;
  reg        [17:0]   img_reg_array_52_61_imag;
  reg        [17:0]   img_reg_array_52_62_real;
  reg        [17:0]   img_reg_array_52_62_imag;
  reg        [17:0]   img_reg_array_52_63_real;
  reg        [17:0]   img_reg_array_52_63_imag;
  reg        [17:0]   img_reg_array_53_0_real;
  reg        [17:0]   img_reg_array_53_0_imag;
  reg        [17:0]   img_reg_array_53_1_real;
  reg        [17:0]   img_reg_array_53_1_imag;
  reg        [17:0]   img_reg_array_53_2_real;
  reg        [17:0]   img_reg_array_53_2_imag;
  reg        [17:0]   img_reg_array_53_3_real;
  reg        [17:0]   img_reg_array_53_3_imag;
  reg        [17:0]   img_reg_array_53_4_real;
  reg        [17:0]   img_reg_array_53_4_imag;
  reg        [17:0]   img_reg_array_53_5_real;
  reg        [17:0]   img_reg_array_53_5_imag;
  reg        [17:0]   img_reg_array_53_6_real;
  reg        [17:0]   img_reg_array_53_6_imag;
  reg        [17:0]   img_reg_array_53_7_real;
  reg        [17:0]   img_reg_array_53_7_imag;
  reg        [17:0]   img_reg_array_53_8_real;
  reg        [17:0]   img_reg_array_53_8_imag;
  reg        [17:0]   img_reg_array_53_9_real;
  reg        [17:0]   img_reg_array_53_9_imag;
  reg        [17:0]   img_reg_array_53_10_real;
  reg        [17:0]   img_reg_array_53_10_imag;
  reg        [17:0]   img_reg_array_53_11_real;
  reg        [17:0]   img_reg_array_53_11_imag;
  reg        [17:0]   img_reg_array_53_12_real;
  reg        [17:0]   img_reg_array_53_12_imag;
  reg        [17:0]   img_reg_array_53_13_real;
  reg        [17:0]   img_reg_array_53_13_imag;
  reg        [17:0]   img_reg_array_53_14_real;
  reg        [17:0]   img_reg_array_53_14_imag;
  reg        [17:0]   img_reg_array_53_15_real;
  reg        [17:0]   img_reg_array_53_15_imag;
  reg        [17:0]   img_reg_array_53_16_real;
  reg        [17:0]   img_reg_array_53_16_imag;
  reg        [17:0]   img_reg_array_53_17_real;
  reg        [17:0]   img_reg_array_53_17_imag;
  reg        [17:0]   img_reg_array_53_18_real;
  reg        [17:0]   img_reg_array_53_18_imag;
  reg        [17:0]   img_reg_array_53_19_real;
  reg        [17:0]   img_reg_array_53_19_imag;
  reg        [17:0]   img_reg_array_53_20_real;
  reg        [17:0]   img_reg_array_53_20_imag;
  reg        [17:0]   img_reg_array_53_21_real;
  reg        [17:0]   img_reg_array_53_21_imag;
  reg        [17:0]   img_reg_array_53_22_real;
  reg        [17:0]   img_reg_array_53_22_imag;
  reg        [17:0]   img_reg_array_53_23_real;
  reg        [17:0]   img_reg_array_53_23_imag;
  reg        [17:0]   img_reg_array_53_24_real;
  reg        [17:0]   img_reg_array_53_24_imag;
  reg        [17:0]   img_reg_array_53_25_real;
  reg        [17:0]   img_reg_array_53_25_imag;
  reg        [17:0]   img_reg_array_53_26_real;
  reg        [17:0]   img_reg_array_53_26_imag;
  reg        [17:0]   img_reg_array_53_27_real;
  reg        [17:0]   img_reg_array_53_27_imag;
  reg        [17:0]   img_reg_array_53_28_real;
  reg        [17:0]   img_reg_array_53_28_imag;
  reg        [17:0]   img_reg_array_53_29_real;
  reg        [17:0]   img_reg_array_53_29_imag;
  reg        [17:0]   img_reg_array_53_30_real;
  reg        [17:0]   img_reg_array_53_30_imag;
  reg        [17:0]   img_reg_array_53_31_real;
  reg        [17:0]   img_reg_array_53_31_imag;
  reg        [17:0]   img_reg_array_53_32_real;
  reg        [17:0]   img_reg_array_53_32_imag;
  reg        [17:0]   img_reg_array_53_33_real;
  reg        [17:0]   img_reg_array_53_33_imag;
  reg        [17:0]   img_reg_array_53_34_real;
  reg        [17:0]   img_reg_array_53_34_imag;
  reg        [17:0]   img_reg_array_53_35_real;
  reg        [17:0]   img_reg_array_53_35_imag;
  reg        [17:0]   img_reg_array_53_36_real;
  reg        [17:0]   img_reg_array_53_36_imag;
  reg        [17:0]   img_reg_array_53_37_real;
  reg        [17:0]   img_reg_array_53_37_imag;
  reg        [17:0]   img_reg_array_53_38_real;
  reg        [17:0]   img_reg_array_53_38_imag;
  reg        [17:0]   img_reg_array_53_39_real;
  reg        [17:0]   img_reg_array_53_39_imag;
  reg        [17:0]   img_reg_array_53_40_real;
  reg        [17:0]   img_reg_array_53_40_imag;
  reg        [17:0]   img_reg_array_53_41_real;
  reg        [17:0]   img_reg_array_53_41_imag;
  reg        [17:0]   img_reg_array_53_42_real;
  reg        [17:0]   img_reg_array_53_42_imag;
  reg        [17:0]   img_reg_array_53_43_real;
  reg        [17:0]   img_reg_array_53_43_imag;
  reg        [17:0]   img_reg_array_53_44_real;
  reg        [17:0]   img_reg_array_53_44_imag;
  reg        [17:0]   img_reg_array_53_45_real;
  reg        [17:0]   img_reg_array_53_45_imag;
  reg        [17:0]   img_reg_array_53_46_real;
  reg        [17:0]   img_reg_array_53_46_imag;
  reg        [17:0]   img_reg_array_53_47_real;
  reg        [17:0]   img_reg_array_53_47_imag;
  reg        [17:0]   img_reg_array_53_48_real;
  reg        [17:0]   img_reg_array_53_48_imag;
  reg        [17:0]   img_reg_array_53_49_real;
  reg        [17:0]   img_reg_array_53_49_imag;
  reg        [17:0]   img_reg_array_53_50_real;
  reg        [17:0]   img_reg_array_53_50_imag;
  reg        [17:0]   img_reg_array_53_51_real;
  reg        [17:0]   img_reg_array_53_51_imag;
  reg        [17:0]   img_reg_array_53_52_real;
  reg        [17:0]   img_reg_array_53_52_imag;
  reg        [17:0]   img_reg_array_53_53_real;
  reg        [17:0]   img_reg_array_53_53_imag;
  reg        [17:0]   img_reg_array_53_54_real;
  reg        [17:0]   img_reg_array_53_54_imag;
  reg        [17:0]   img_reg_array_53_55_real;
  reg        [17:0]   img_reg_array_53_55_imag;
  reg        [17:0]   img_reg_array_53_56_real;
  reg        [17:0]   img_reg_array_53_56_imag;
  reg        [17:0]   img_reg_array_53_57_real;
  reg        [17:0]   img_reg_array_53_57_imag;
  reg        [17:0]   img_reg_array_53_58_real;
  reg        [17:0]   img_reg_array_53_58_imag;
  reg        [17:0]   img_reg_array_53_59_real;
  reg        [17:0]   img_reg_array_53_59_imag;
  reg        [17:0]   img_reg_array_53_60_real;
  reg        [17:0]   img_reg_array_53_60_imag;
  reg        [17:0]   img_reg_array_53_61_real;
  reg        [17:0]   img_reg_array_53_61_imag;
  reg        [17:0]   img_reg_array_53_62_real;
  reg        [17:0]   img_reg_array_53_62_imag;
  reg        [17:0]   img_reg_array_53_63_real;
  reg        [17:0]   img_reg_array_53_63_imag;
  reg        [17:0]   img_reg_array_54_0_real;
  reg        [17:0]   img_reg_array_54_0_imag;
  reg        [17:0]   img_reg_array_54_1_real;
  reg        [17:0]   img_reg_array_54_1_imag;
  reg        [17:0]   img_reg_array_54_2_real;
  reg        [17:0]   img_reg_array_54_2_imag;
  reg        [17:0]   img_reg_array_54_3_real;
  reg        [17:0]   img_reg_array_54_3_imag;
  reg        [17:0]   img_reg_array_54_4_real;
  reg        [17:0]   img_reg_array_54_4_imag;
  reg        [17:0]   img_reg_array_54_5_real;
  reg        [17:0]   img_reg_array_54_5_imag;
  reg        [17:0]   img_reg_array_54_6_real;
  reg        [17:0]   img_reg_array_54_6_imag;
  reg        [17:0]   img_reg_array_54_7_real;
  reg        [17:0]   img_reg_array_54_7_imag;
  reg        [17:0]   img_reg_array_54_8_real;
  reg        [17:0]   img_reg_array_54_8_imag;
  reg        [17:0]   img_reg_array_54_9_real;
  reg        [17:0]   img_reg_array_54_9_imag;
  reg        [17:0]   img_reg_array_54_10_real;
  reg        [17:0]   img_reg_array_54_10_imag;
  reg        [17:0]   img_reg_array_54_11_real;
  reg        [17:0]   img_reg_array_54_11_imag;
  reg        [17:0]   img_reg_array_54_12_real;
  reg        [17:0]   img_reg_array_54_12_imag;
  reg        [17:0]   img_reg_array_54_13_real;
  reg        [17:0]   img_reg_array_54_13_imag;
  reg        [17:0]   img_reg_array_54_14_real;
  reg        [17:0]   img_reg_array_54_14_imag;
  reg        [17:0]   img_reg_array_54_15_real;
  reg        [17:0]   img_reg_array_54_15_imag;
  reg        [17:0]   img_reg_array_54_16_real;
  reg        [17:0]   img_reg_array_54_16_imag;
  reg        [17:0]   img_reg_array_54_17_real;
  reg        [17:0]   img_reg_array_54_17_imag;
  reg        [17:0]   img_reg_array_54_18_real;
  reg        [17:0]   img_reg_array_54_18_imag;
  reg        [17:0]   img_reg_array_54_19_real;
  reg        [17:0]   img_reg_array_54_19_imag;
  reg        [17:0]   img_reg_array_54_20_real;
  reg        [17:0]   img_reg_array_54_20_imag;
  reg        [17:0]   img_reg_array_54_21_real;
  reg        [17:0]   img_reg_array_54_21_imag;
  reg        [17:0]   img_reg_array_54_22_real;
  reg        [17:0]   img_reg_array_54_22_imag;
  reg        [17:0]   img_reg_array_54_23_real;
  reg        [17:0]   img_reg_array_54_23_imag;
  reg        [17:0]   img_reg_array_54_24_real;
  reg        [17:0]   img_reg_array_54_24_imag;
  reg        [17:0]   img_reg_array_54_25_real;
  reg        [17:0]   img_reg_array_54_25_imag;
  reg        [17:0]   img_reg_array_54_26_real;
  reg        [17:0]   img_reg_array_54_26_imag;
  reg        [17:0]   img_reg_array_54_27_real;
  reg        [17:0]   img_reg_array_54_27_imag;
  reg        [17:0]   img_reg_array_54_28_real;
  reg        [17:0]   img_reg_array_54_28_imag;
  reg        [17:0]   img_reg_array_54_29_real;
  reg        [17:0]   img_reg_array_54_29_imag;
  reg        [17:0]   img_reg_array_54_30_real;
  reg        [17:0]   img_reg_array_54_30_imag;
  reg        [17:0]   img_reg_array_54_31_real;
  reg        [17:0]   img_reg_array_54_31_imag;
  reg        [17:0]   img_reg_array_54_32_real;
  reg        [17:0]   img_reg_array_54_32_imag;
  reg        [17:0]   img_reg_array_54_33_real;
  reg        [17:0]   img_reg_array_54_33_imag;
  reg        [17:0]   img_reg_array_54_34_real;
  reg        [17:0]   img_reg_array_54_34_imag;
  reg        [17:0]   img_reg_array_54_35_real;
  reg        [17:0]   img_reg_array_54_35_imag;
  reg        [17:0]   img_reg_array_54_36_real;
  reg        [17:0]   img_reg_array_54_36_imag;
  reg        [17:0]   img_reg_array_54_37_real;
  reg        [17:0]   img_reg_array_54_37_imag;
  reg        [17:0]   img_reg_array_54_38_real;
  reg        [17:0]   img_reg_array_54_38_imag;
  reg        [17:0]   img_reg_array_54_39_real;
  reg        [17:0]   img_reg_array_54_39_imag;
  reg        [17:0]   img_reg_array_54_40_real;
  reg        [17:0]   img_reg_array_54_40_imag;
  reg        [17:0]   img_reg_array_54_41_real;
  reg        [17:0]   img_reg_array_54_41_imag;
  reg        [17:0]   img_reg_array_54_42_real;
  reg        [17:0]   img_reg_array_54_42_imag;
  reg        [17:0]   img_reg_array_54_43_real;
  reg        [17:0]   img_reg_array_54_43_imag;
  reg        [17:0]   img_reg_array_54_44_real;
  reg        [17:0]   img_reg_array_54_44_imag;
  reg        [17:0]   img_reg_array_54_45_real;
  reg        [17:0]   img_reg_array_54_45_imag;
  reg        [17:0]   img_reg_array_54_46_real;
  reg        [17:0]   img_reg_array_54_46_imag;
  reg        [17:0]   img_reg_array_54_47_real;
  reg        [17:0]   img_reg_array_54_47_imag;
  reg        [17:0]   img_reg_array_54_48_real;
  reg        [17:0]   img_reg_array_54_48_imag;
  reg        [17:0]   img_reg_array_54_49_real;
  reg        [17:0]   img_reg_array_54_49_imag;
  reg        [17:0]   img_reg_array_54_50_real;
  reg        [17:0]   img_reg_array_54_50_imag;
  reg        [17:0]   img_reg_array_54_51_real;
  reg        [17:0]   img_reg_array_54_51_imag;
  reg        [17:0]   img_reg_array_54_52_real;
  reg        [17:0]   img_reg_array_54_52_imag;
  reg        [17:0]   img_reg_array_54_53_real;
  reg        [17:0]   img_reg_array_54_53_imag;
  reg        [17:0]   img_reg_array_54_54_real;
  reg        [17:0]   img_reg_array_54_54_imag;
  reg        [17:0]   img_reg_array_54_55_real;
  reg        [17:0]   img_reg_array_54_55_imag;
  reg        [17:0]   img_reg_array_54_56_real;
  reg        [17:0]   img_reg_array_54_56_imag;
  reg        [17:0]   img_reg_array_54_57_real;
  reg        [17:0]   img_reg_array_54_57_imag;
  reg        [17:0]   img_reg_array_54_58_real;
  reg        [17:0]   img_reg_array_54_58_imag;
  reg        [17:0]   img_reg_array_54_59_real;
  reg        [17:0]   img_reg_array_54_59_imag;
  reg        [17:0]   img_reg_array_54_60_real;
  reg        [17:0]   img_reg_array_54_60_imag;
  reg        [17:0]   img_reg_array_54_61_real;
  reg        [17:0]   img_reg_array_54_61_imag;
  reg        [17:0]   img_reg_array_54_62_real;
  reg        [17:0]   img_reg_array_54_62_imag;
  reg        [17:0]   img_reg_array_54_63_real;
  reg        [17:0]   img_reg_array_54_63_imag;
  reg        [17:0]   img_reg_array_55_0_real;
  reg        [17:0]   img_reg_array_55_0_imag;
  reg        [17:0]   img_reg_array_55_1_real;
  reg        [17:0]   img_reg_array_55_1_imag;
  reg        [17:0]   img_reg_array_55_2_real;
  reg        [17:0]   img_reg_array_55_2_imag;
  reg        [17:0]   img_reg_array_55_3_real;
  reg        [17:0]   img_reg_array_55_3_imag;
  reg        [17:0]   img_reg_array_55_4_real;
  reg        [17:0]   img_reg_array_55_4_imag;
  reg        [17:0]   img_reg_array_55_5_real;
  reg        [17:0]   img_reg_array_55_5_imag;
  reg        [17:0]   img_reg_array_55_6_real;
  reg        [17:0]   img_reg_array_55_6_imag;
  reg        [17:0]   img_reg_array_55_7_real;
  reg        [17:0]   img_reg_array_55_7_imag;
  reg        [17:0]   img_reg_array_55_8_real;
  reg        [17:0]   img_reg_array_55_8_imag;
  reg        [17:0]   img_reg_array_55_9_real;
  reg        [17:0]   img_reg_array_55_9_imag;
  reg        [17:0]   img_reg_array_55_10_real;
  reg        [17:0]   img_reg_array_55_10_imag;
  reg        [17:0]   img_reg_array_55_11_real;
  reg        [17:0]   img_reg_array_55_11_imag;
  reg        [17:0]   img_reg_array_55_12_real;
  reg        [17:0]   img_reg_array_55_12_imag;
  reg        [17:0]   img_reg_array_55_13_real;
  reg        [17:0]   img_reg_array_55_13_imag;
  reg        [17:0]   img_reg_array_55_14_real;
  reg        [17:0]   img_reg_array_55_14_imag;
  reg        [17:0]   img_reg_array_55_15_real;
  reg        [17:0]   img_reg_array_55_15_imag;
  reg        [17:0]   img_reg_array_55_16_real;
  reg        [17:0]   img_reg_array_55_16_imag;
  reg        [17:0]   img_reg_array_55_17_real;
  reg        [17:0]   img_reg_array_55_17_imag;
  reg        [17:0]   img_reg_array_55_18_real;
  reg        [17:0]   img_reg_array_55_18_imag;
  reg        [17:0]   img_reg_array_55_19_real;
  reg        [17:0]   img_reg_array_55_19_imag;
  reg        [17:0]   img_reg_array_55_20_real;
  reg        [17:0]   img_reg_array_55_20_imag;
  reg        [17:0]   img_reg_array_55_21_real;
  reg        [17:0]   img_reg_array_55_21_imag;
  reg        [17:0]   img_reg_array_55_22_real;
  reg        [17:0]   img_reg_array_55_22_imag;
  reg        [17:0]   img_reg_array_55_23_real;
  reg        [17:0]   img_reg_array_55_23_imag;
  reg        [17:0]   img_reg_array_55_24_real;
  reg        [17:0]   img_reg_array_55_24_imag;
  reg        [17:0]   img_reg_array_55_25_real;
  reg        [17:0]   img_reg_array_55_25_imag;
  reg        [17:0]   img_reg_array_55_26_real;
  reg        [17:0]   img_reg_array_55_26_imag;
  reg        [17:0]   img_reg_array_55_27_real;
  reg        [17:0]   img_reg_array_55_27_imag;
  reg        [17:0]   img_reg_array_55_28_real;
  reg        [17:0]   img_reg_array_55_28_imag;
  reg        [17:0]   img_reg_array_55_29_real;
  reg        [17:0]   img_reg_array_55_29_imag;
  reg        [17:0]   img_reg_array_55_30_real;
  reg        [17:0]   img_reg_array_55_30_imag;
  reg        [17:0]   img_reg_array_55_31_real;
  reg        [17:0]   img_reg_array_55_31_imag;
  reg        [17:0]   img_reg_array_55_32_real;
  reg        [17:0]   img_reg_array_55_32_imag;
  reg        [17:0]   img_reg_array_55_33_real;
  reg        [17:0]   img_reg_array_55_33_imag;
  reg        [17:0]   img_reg_array_55_34_real;
  reg        [17:0]   img_reg_array_55_34_imag;
  reg        [17:0]   img_reg_array_55_35_real;
  reg        [17:0]   img_reg_array_55_35_imag;
  reg        [17:0]   img_reg_array_55_36_real;
  reg        [17:0]   img_reg_array_55_36_imag;
  reg        [17:0]   img_reg_array_55_37_real;
  reg        [17:0]   img_reg_array_55_37_imag;
  reg        [17:0]   img_reg_array_55_38_real;
  reg        [17:0]   img_reg_array_55_38_imag;
  reg        [17:0]   img_reg_array_55_39_real;
  reg        [17:0]   img_reg_array_55_39_imag;
  reg        [17:0]   img_reg_array_55_40_real;
  reg        [17:0]   img_reg_array_55_40_imag;
  reg        [17:0]   img_reg_array_55_41_real;
  reg        [17:0]   img_reg_array_55_41_imag;
  reg        [17:0]   img_reg_array_55_42_real;
  reg        [17:0]   img_reg_array_55_42_imag;
  reg        [17:0]   img_reg_array_55_43_real;
  reg        [17:0]   img_reg_array_55_43_imag;
  reg        [17:0]   img_reg_array_55_44_real;
  reg        [17:0]   img_reg_array_55_44_imag;
  reg        [17:0]   img_reg_array_55_45_real;
  reg        [17:0]   img_reg_array_55_45_imag;
  reg        [17:0]   img_reg_array_55_46_real;
  reg        [17:0]   img_reg_array_55_46_imag;
  reg        [17:0]   img_reg_array_55_47_real;
  reg        [17:0]   img_reg_array_55_47_imag;
  reg        [17:0]   img_reg_array_55_48_real;
  reg        [17:0]   img_reg_array_55_48_imag;
  reg        [17:0]   img_reg_array_55_49_real;
  reg        [17:0]   img_reg_array_55_49_imag;
  reg        [17:0]   img_reg_array_55_50_real;
  reg        [17:0]   img_reg_array_55_50_imag;
  reg        [17:0]   img_reg_array_55_51_real;
  reg        [17:0]   img_reg_array_55_51_imag;
  reg        [17:0]   img_reg_array_55_52_real;
  reg        [17:0]   img_reg_array_55_52_imag;
  reg        [17:0]   img_reg_array_55_53_real;
  reg        [17:0]   img_reg_array_55_53_imag;
  reg        [17:0]   img_reg_array_55_54_real;
  reg        [17:0]   img_reg_array_55_54_imag;
  reg        [17:0]   img_reg_array_55_55_real;
  reg        [17:0]   img_reg_array_55_55_imag;
  reg        [17:0]   img_reg_array_55_56_real;
  reg        [17:0]   img_reg_array_55_56_imag;
  reg        [17:0]   img_reg_array_55_57_real;
  reg        [17:0]   img_reg_array_55_57_imag;
  reg        [17:0]   img_reg_array_55_58_real;
  reg        [17:0]   img_reg_array_55_58_imag;
  reg        [17:0]   img_reg_array_55_59_real;
  reg        [17:0]   img_reg_array_55_59_imag;
  reg        [17:0]   img_reg_array_55_60_real;
  reg        [17:0]   img_reg_array_55_60_imag;
  reg        [17:0]   img_reg_array_55_61_real;
  reg        [17:0]   img_reg_array_55_61_imag;
  reg        [17:0]   img_reg_array_55_62_real;
  reg        [17:0]   img_reg_array_55_62_imag;
  reg        [17:0]   img_reg_array_55_63_real;
  reg        [17:0]   img_reg_array_55_63_imag;
  reg        [17:0]   img_reg_array_56_0_real;
  reg        [17:0]   img_reg_array_56_0_imag;
  reg        [17:0]   img_reg_array_56_1_real;
  reg        [17:0]   img_reg_array_56_1_imag;
  reg        [17:0]   img_reg_array_56_2_real;
  reg        [17:0]   img_reg_array_56_2_imag;
  reg        [17:0]   img_reg_array_56_3_real;
  reg        [17:0]   img_reg_array_56_3_imag;
  reg        [17:0]   img_reg_array_56_4_real;
  reg        [17:0]   img_reg_array_56_4_imag;
  reg        [17:0]   img_reg_array_56_5_real;
  reg        [17:0]   img_reg_array_56_5_imag;
  reg        [17:0]   img_reg_array_56_6_real;
  reg        [17:0]   img_reg_array_56_6_imag;
  reg        [17:0]   img_reg_array_56_7_real;
  reg        [17:0]   img_reg_array_56_7_imag;
  reg        [17:0]   img_reg_array_56_8_real;
  reg        [17:0]   img_reg_array_56_8_imag;
  reg        [17:0]   img_reg_array_56_9_real;
  reg        [17:0]   img_reg_array_56_9_imag;
  reg        [17:0]   img_reg_array_56_10_real;
  reg        [17:0]   img_reg_array_56_10_imag;
  reg        [17:0]   img_reg_array_56_11_real;
  reg        [17:0]   img_reg_array_56_11_imag;
  reg        [17:0]   img_reg_array_56_12_real;
  reg        [17:0]   img_reg_array_56_12_imag;
  reg        [17:0]   img_reg_array_56_13_real;
  reg        [17:0]   img_reg_array_56_13_imag;
  reg        [17:0]   img_reg_array_56_14_real;
  reg        [17:0]   img_reg_array_56_14_imag;
  reg        [17:0]   img_reg_array_56_15_real;
  reg        [17:0]   img_reg_array_56_15_imag;
  reg        [17:0]   img_reg_array_56_16_real;
  reg        [17:0]   img_reg_array_56_16_imag;
  reg        [17:0]   img_reg_array_56_17_real;
  reg        [17:0]   img_reg_array_56_17_imag;
  reg        [17:0]   img_reg_array_56_18_real;
  reg        [17:0]   img_reg_array_56_18_imag;
  reg        [17:0]   img_reg_array_56_19_real;
  reg        [17:0]   img_reg_array_56_19_imag;
  reg        [17:0]   img_reg_array_56_20_real;
  reg        [17:0]   img_reg_array_56_20_imag;
  reg        [17:0]   img_reg_array_56_21_real;
  reg        [17:0]   img_reg_array_56_21_imag;
  reg        [17:0]   img_reg_array_56_22_real;
  reg        [17:0]   img_reg_array_56_22_imag;
  reg        [17:0]   img_reg_array_56_23_real;
  reg        [17:0]   img_reg_array_56_23_imag;
  reg        [17:0]   img_reg_array_56_24_real;
  reg        [17:0]   img_reg_array_56_24_imag;
  reg        [17:0]   img_reg_array_56_25_real;
  reg        [17:0]   img_reg_array_56_25_imag;
  reg        [17:0]   img_reg_array_56_26_real;
  reg        [17:0]   img_reg_array_56_26_imag;
  reg        [17:0]   img_reg_array_56_27_real;
  reg        [17:0]   img_reg_array_56_27_imag;
  reg        [17:0]   img_reg_array_56_28_real;
  reg        [17:0]   img_reg_array_56_28_imag;
  reg        [17:0]   img_reg_array_56_29_real;
  reg        [17:0]   img_reg_array_56_29_imag;
  reg        [17:0]   img_reg_array_56_30_real;
  reg        [17:0]   img_reg_array_56_30_imag;
  reg        [17:0]   img_reg_array_56_31_real;
  reg        [17:0]   img_reg_array_56_31_imag;
  reg        [17:0]   img_reg_array_56_32_real;
  reg        [17:0]   img_reg_array_56_32_imag;
  reg        [17:0]   img_reg_array_56_33_real;
  reg        [17:0]   img_reg_array_56_33_imag;
  reg        [17:0]   img_reg_array_56_34_real;
  reg        [17:0]   img_reg_array_56_34_imag;
  reg        [17:0]   img_reg_array_56_35_real;
  reg        [17:0]   img_reg_array_56_35_imag;
  reg        [17:0]   img_reg_array_56_36_real;
  reg        [17:0]   img_reg_array_56_36_imag;
  reg        [17:0]   img_reg_array_56_37_real;
  reg        [17:0]   img_reg_array_56_37_imag;
  reg        [17:0]   img_reg_array_56_38_real;
  reg        [17:0]   img_reg_array_56_38_imag;
  reg        [17:0]   img_reg_array_56_39_real;
  reg        [17:0]   img_reg_array_56_39_imag;
  reg        [17:0]   img_reg_array_56_40_real;
  reg        [17:0]   img_reg_array_56_40_imag;
  reg        [17:0]   img_reg_array_56_41_real;
  reg        [17:0]   img_reg_array_56_41_imag;
  reg        [17:0]   img_reg_array_56_42_real;
  reg        [17:0]   img_reg_array_56_42_imag;
  reg        [17:0]   img_reg_array_56_43_real;
  reg        [17:0]   img_reg_array_56_43_imag;
  reg        [17:0]   img_reg_array_56_44_real;
  reg        [17:0]   img_reg_array_56_44_imag;
  reg        [17:0]   img_reg_array_56_45_real;
  reg        [17:0]   img_reg_array_56_45_imag;
  reg        [17:0]   img_reg_array_56_46_real;
  reg        [17:0]   img_reg_array_56_46_imag;
  reg        [17:0]   img_reg_array_56_47_real;
  reg        [17:0]   img_reg_array_56_47_imag;
  reg        [17:0]   img_reg_array_56_48_real;
  reg        [17:0]   img_reg_array_56_48_imag;
  reg        [17:0]   img_reg_array_56_49_real;
  reg        [17:0]   img_reg_array_56_49_imag;
  reg        [17:0]   img_reg_array_56_50_real;
  reg        [17:0]   img_reg_array_56_50_imag;
  reg        [17:0]   img_reg_array_56_51_real;
  reg        [17:0]   img_reg_array_56_51_imag;
  reg        [17:0]   img_reg_array_56_52_real;
  reg        [17:0]   img_reg_array_56_52_imag;
  reg        [17:0]   img_reg_array_56_53_real;
  reg        [17:0]   img_reg_array_56_53_imag;
  reg        [17:0]   img_reg_array_56_54_real;
  reg        [17:0]   img_reg_array_56_54_imag;
  reg        [17:0]   img_reg_array_56_55_real;
  reg        [17:0]   img_reg_array_56_55_imag;
  reg        [17:0]   img_reg_array_56_56_real;
  reg        [17:0]   img_reg_array_56_56_imag;
  reg        [17:0]   img_reg_array_56_57_real;
  reg        [17:0]   img_reg_array_56_57_imag;
  reg        [17:0]   img_reg_array_56_58_real;
  reg        [17:0]   img_reg_array_56_58_imag;
  reg        [17:0]   img_reg_array_56_59_real;
  reg        [17:0]   img_reg_array_56_59_imag;
  reg        [17:0]   img_reg_array_56_60_real;
  reg        [17:0]   img_reg_array_56_60_imag;
  reg        [17:0]   img_reg_array_56_61_real;
  reg        [17:0]   img_reg_array_56_61_imag;
  reg        [17:0]   img_reg_array_56_62_real;
  reg        [17:0]   img_reg_array_56_62_imag;
  reg        [17:0]   img_reg_array_56_63_real;
  reg        [17:0]   img_reg_array_56_63_imag;
  reg        [17:0]   img_reg_array_57_0_real;
  reg        [17:0]   img_reg_array_57_0_imag;
  reg        [17:0]   img_reg_array_57_1_real;
  reg        [17:0]   img_reg_array_57_1_imag;
  reg        [17:0]   img_reg_array_57_2_real;
  reg        [17:0]   img_reg_array_57_2_imag;
  reg        [17:0]   img_reg_array_57_3_real;
  reg        [17:0]   img_reg_array_57_3_imag;
  reg        [17:0]   img_reg_array_57_4_real;
  reg        [17:0]   img_reg_array_57_4_imag;
  reg        [17:0]   img_reg_array_57_5_real;
  reg        [17:0]   img_reg_array_57_5_imag;
  reg        [17:0]   img_reg_array_57_6_real;
  reg        [17:0]   img_reg_array_57_6_imag;
  reg        [17:0]   img_reg_array_57_7_real;
  reg        [17:0]   img_reg_array_57_7_imag;
  reg        [17:0]   img_reg_array_57_8_real;
  reg        [17:0]   img_reg_array_57_8_imag;
  reg        [17:0]   img_reg_array_57_9_real;
  reg        [17:0]   img_reg_array_57_9_imag;
  reg        [17:0]   img_reg_array_57_10_real;
  reg        [17:0]   img_reg_array_57_10_imag;
  reg        [17:0]   img_reg_array_57_11_real;
  reg        [17:0]   img_reg_array_57_11_imag;
  reg        [17:0]   img_reg_array_57_12_real;
  reg        [17:0]   img_reg_array_57_12_imag;
  reg        [17:0]   img_reg_array_57_13_real;
  reg        [17:0]   img_reg_array_57_13_imag;
  reg        [17:0]   img_reg_array_57_14_real;
  reg        [17:0]   img_reg_array_57_14_imag;
  reg        [17:0]   img_reg_array_57_15_real;
  reg        [17:0]   img_reg_array_57_15_imag;
  reg        [17:0]   img_reg_array_57_16_real;
  reg        [17:0]   img_reg_array_57_16_imag;
  reg        [17:0]   img_reg_array_57_17_real;
  reg        [17:0]   img_reg_array_57_17_imag;
  reg        [17:0]   img_reg_array_57_18_real;
  reg        [17:0]   img_reg_array_57_18_imag;
  reg        [17:0]   img_reg_array_57_19_real;
  reg        [17:0]   img_reg_array_57_19_imag;
  reg        [17:0]   img_reg_array_57_20_real;
  reg        [17:0]   img_reg_array_57_20_imag;
  reg        [17:0]   img_reg_array_57_21_real;
  reg        [17:0]   img_reg_array_57_21_imag;
  reg        [17:0]   img_reg_array_57_22_real;
  reg        [17:0]   img_reg_array_57_22_imag;
  reg        [17:0]   img_reg_array_57_23_real;
  reg        [17:0]   img_reg_array_57_23_imag;
  reg        [17:0]   img_reg_array_57_24_real;
  reg        [17:0]   img_reg_array_57_24_imag;
  reg        [17:0]   img_reg_array_57_25_real;
  reg        [17:0]   img_reg_array_57_25_imag;
  reg        [17:0]   img_reg_array_57_26_real;
  reg        [17:0]   img_reg_array_57_26_imag;
  reg        [17:0]   img_reg_array_57_27_real;
  reg        [17:0]   img_reg_array_57_27_imag;
  reg        [17:0]   img_reg_array_57_28_real;
  reg        [17:0]   img_reg_array_57_28_imag;
  reg        [17:0]   img_reg_array_57_29_real;
  reg        [17:0]   img_reg_array_57_29_imag;
  reg        [17:0]   img_reg_array_57_30_real;
  reg        [17:0]   img_reg_array_57_30_imag;
  reg        [17:0]   img_reg_array_57_31_real;
  reg        [17:0]   img_reg_array_57_31_imag;
  reg        [17:0]   img_reg_array_57_32_real;
  reg        [17:0]   img_reg_array_57_32_imag;
  reg        [17:0]   img_reg_array_57_33_real;
  reg        [17:0]   img_reg_array_57_33_imag;
  reg        [17:0]   img_reg_array_57_34_real;
  reg        [17:0]   img_reg_array_57_34_imag;
  reg        [17:0]   img_reg_array_57_35_real;
  reg        [17:0]   img_reg_array_57_35_imag;
  reg        [17:0]   img_reg_array_57_36_real;
  reg        [17:0]   img_reg_array_57_36_imag;
  reg        [17:0]   img_reg_array_57_37_real;
  reg        [17:0]   img_reg_array_57_37_imag;
  reg        [17:0]   img_reg_array_57_38_real;
  reg        [17:0]   img_reg_array_57_38_imag;
  reg        [17:0]   img_reg_array_57_39_real;
  reg        [17:0]   img_reg_array_57_39_imag;
  reg        [17:0]   img_reg_array_57_40_real;
  reg        [17:0]   img_reg_array_57_40_imag;
  reg        [17:0]   img_reg_array_57_41_real;
  reg        [17:0]   img_reg_array_57_41_imag;
  reg        [17:0]   img_reg_array_57_42_real;
  reg        [17:0]   img_reg_array_57_42_imag;
  reg        [17:0]   img_reg_array_57_43_real;
  reg        [17:0]   img_reg_array_57_43_imag;
  reg        [17:0]   img_reg_array_57_44_real;
  reg        [17:0]   img_reg_array_57_44_imag;
  reg        [17:0]   img_reg_array_57_45_real;
  reg        [17:0]   img_reg_array_57_45_imag;
  reg        [17:0]   img_reg_array_57_46_real;
  reg        [17:0]   img_reg_array_57_46_imag;
  reg        [17:0]   img_reg_array_57_47_real;
  reg        [17:0]   img_reg_array_57_47_imag;
  reg        [17:0]   img_reg_array_57_48_real;
  reg        [17:0]   img_reg_array_57_48_imag;
  reg        [17:0]   img_reg_array_57_49_real;
  reg        [17:0]   img_reg_array_57_49_imag;
  reg        [17:0]   img_reg_array_57_50_real;
  reg        [17:0]   img_reg_array_57_50_imag;
  reg        [17:0]   img_reg_array_57_51_real;
  reg        [17:0]   img_reg_array_57_51_imag;
  reg        [17:0]   img_reg_array_57_52_real;
  reg        [17:0]   img_reg_array_57_52_imag;
  reg        [17:0]   img_reg_array_57_53_real;
  reg        [17:0]   img_reg_array_57_53_imag;
  reg        [17:0]   img_reg_array_57_54_real;
  reg        [17:0]   img_reg_array_57_54_imag;
  reg        [17:0]   img_reg_array_57_55_real;
  reg        [17:0]   img_reg_array_57_55_imag;
  reg        [17:0]   img_reg_array_57_56_real;
  reg        [17:0]   img_reg_array_57_56_imag;
  reg        [17:0]   img_reg_array_57_57_real;
  reg        [17:0]   img_reg_array_57_57_imag;
  reg        [17:0]   img_reg_array_57_58_real;
  reg        [17:0]   img_reg_array_57_58_imag;
  reg        [17:0]   img_reg_array_57_59_real;
  reg        [17:0]   img_reg_array_57_59_imag;
  reg        [17:0]   img_reg_array_57_60_real;
  reg        [17:0]   img_reg_array_57_60_imag;
  reg        [17:0]   img_reg_array_57_61_real;
  reg        [17:0]   img_reg_array_57_61_imag;
  reg        [17:0]   img_reg_array_57_62_real;
  reg        [17:0]   img_reg_array_57_62_imag;
  reg        [17:0]   img_reg_array_57_63_real;
  reg        [17:0]   img_reg_array_57_63_imag;
  reg        [17:0]   img_reg_array_58_0_real;
  reg        [17:0]   img_reg_array_58_0_imag;
  reg        [17:0]   img_reg_array_58_1_real;
  reg        [17:0]   img_reg_array_58_1_imag;
  reg        [17:0]   img_reg_array_58_2_real;
  reg        [17:0]   img_reg_array_58_2_imag;
  reg        [17:0]   img_reg_array_58_3_real;
  reg        [17:0]   img_reg_array_58_3_imag;
  reg        [17:0]   img_reg_array_58_4_real;
  reg        [17:0]   img_reg_array_58_4_imag;
  reg        [17:0]   img_reg_array_58_5_real;
  reg        [17:0]   img_reg_array_58_5_imag;
  reg        [17:0]   img_reg_array_58_6_real;
  reg        [17:0]   img_reg_array_58_6_imag;
  reg        [17:0]   img_reg_array_58_7_real;
  reg        [17:0]   img_reg_array_58_7_imag;
  reg        [17:0]   img_reg_array_58_8_real;
  reg        [17:0]   img_reg_array_58_8_imag;
  reg        [17:0]   img_reg_array_58_9_real;
  reg        [17:0]   img_reg_array_58_9_imag;
  reg        [17:0]   img_reg_array_58_10_real;
  reg        [17:0]   img_reg_array_58_10_imag;
  reg        [17:0]   img_reg_array_58_11_real;
  reg        [17:0]   img_reg_array_58_11_imag;
  reg        [17:0]   img_reg_array_58_12_real;
  reg        [17:0]   img_reg_array_58_12_imag;
  reg        [17:0]   img_reg_array_58_13_real;
  reg        [17:0]   img_reg_array_58_13_imag;
  reg        [17:0]   img_reg_array_58_14_real;
  reg        [17:0]   img_reg_array_58_14_imag;
  reg        [17:0]   img_reg_array_58_15_real;
  reg        [17:0]   img_reg_array_58_15_imag;
  reg        [17:0]   img_reg_array_58_16_real;
  reg        [17:0]   img_reg_array_58_16_imag;
  reg        [17:0]   img_reg_array_58_17_real;
  reg        [17:0]   img_reg_array_58_17_imag;
  reg        [17:0]   img_reg_array_58_18_real;
  reg        [17:0]   img_reg_array_58_18_imag;
  reg        [17:0]   img_reg_array_58_19_real;
  reg        [17:0]   img_reg_array_58_19_imag;
  reg        [17:0]   img_reg_array_58_20_real;
  reg        [17:0]   img_reg_array_58_20_imag;
  reg        [17:0]   img_reg_array_58_21_real;
  reg        [17:0]   img_reg_array_58_21_imag;
  reg        [17:0]   img_reg_array_58_22_real;
  reg        [17:0]   img_reg_array_58_22_imag;
  reg        [17:0]   img_reg_array_58_23_real;
  reg        [17:0]   img_reg_array_58_23_imag;
  reg        [17:0]   img_reg_array_58_24_real;
  reg        [17:0]   img_reg_array_58_24_imag;
  reg        [17:0]   img_reg_array_58_25_real;
  reg        [17:0]   img_reg_array_58_25_imag;
  reg        [17:0]   img_reg_array_58_26_real;
  reg        [17:0]   img_reg_array_58_26_imag;
  reg        [17:0]   img_reg_array_58_27_real;
  reg        [17:0]   img_reg_array_58_27_imag;
  reg        [17:0]   img_reg_array_58_28_real;
  reg        [17:0]   img_reg_array_58_28_imag;
  reg        [17:0]   img_reg_array_58_29_real;
  reg        [17:0]   img_reg_array_58_29_imag;
  reg        [17:0]   img_reg_array_58_30_real;
  reg        [17:0]   img_reg_array_58_30_imag;
  reg        [17:0]   img_reg_array_58_31_real;
  reg        [17:0]   img_reg_array_58_31_imag;
  reg        [17:0]   img_reg_array_58_32_real;
  reg        [17:0]   img_reg_array_58_32_imag;
  reg        [17:0]   img_reg_array_58_33_real;
  reg        [17:0]   img_reg_array_58_33_imag;
  reg        [17:0]   img_reg_array_58_34_real;
  reg        [17:0]   img_reg_array_58_34_imag;
  reg        [17:0]   img_reg_array_58_35_real;
  reg        [17:0]   img_reg_array_58_35_imag;
  reg        [17:0]   img_reg_array_58_36_real;
  reg        [17:0]   img_reg_array_58_36_imag;
  reg        [17:0]   img_reg_array_58_37_real;
  reg        [17:0]   img_reg_array_58_37_imag;
  reg        [17:0]   img_reg_array_58_38_real;
  reg        [17:0]   img_reg_array_58_38_imag;
  reg        [17:0]   img_reg_array_58_39_real;
  reg        [17:0]   img_reg_array_58_39_imag;
  reg        [17:0]   img_reg_array_58_40_real;
  reg        [17:0]   img_reg_array_58_40_imag;
  reg        [17:0]   img_reg_array_58_41_real;
  reg        [17:0]   img_reg_array_58_41_imag;
  reg        [17:0]   img_reg_array_58_42_real;
  reg        [17:0]   img_reg_array_58_42_imag;
  reg        [17:0]   img_reg_array_58_43_real;
  reg        [17:0]   img_reg_array_58_43_imag;
  reg        [17:0]   img_reg_array_58_44_real;
  reg        [17:0]   img_reg_array_58_44_imag;
  reg        [17:0]   img_reg_array_58_45_real;
  reg        [17:0]   img_reg_array_58_45_imag;
  reg        [17:0]   img_reg_array_58_46_real;
  reg        [17:0]   img_reg_array_58_46_imag;
  reg        [17:0]   img_reg_array_58_47_real;
  reg        [17:0]   img_reg_array_58_47_imag;
  reg        [17:0]   img_reg_array_58_48_real;
  reg        [17:0]   img_reg_array_58_48_imag;
  reg        [17:0]   img_reg_array_58_49_real;
  reg        [17:0]   img_reg_array_58_49_imag;
  reg        [17:0]   img_reg_array_58_50_real;
  reg        [17:0]   img_reg_array_58_50_imag;
  reg        [17:0]   img_reg_array_58_51_real;
  reg        [17:0]   img_reg_array_58_51_imag;
  reg        [17:0]   img_reg_array_58_52_real;
  reg        [17:0]   img_reg_array_58_52_imag;
  reg        [17:0]   img_reg_array_58_53_real;
  reg        [17:0]   img_reg_array_58_53_imag;
  reg        [17:0]   img_reg_array_58_54_real;
  reg        [17:0]   img_reg_array_58_54_imag;
  reg        [17:0]   img_reg_array_58_55_real;
  reg        [17:0]   img_reg_array_58_55_imag;
  reg        [17:0]   img_reg_array_58_56_real;
  reg        [17:0]   img_reg_array_58_56_imag;
  reg        [17:0]   img_reg_array_58_57_real;
  reg        [17:0]   img_reg_array_58_57_imag;
  reg        [17:0]   img_reg_array_58_58_real;
  reg        [17:0]   img_reg_array_58_58_imag;
  reg        [17:0]   img_reg_array_58_59_real;
  reg        [17:0]   img_reg_array_58_59_imag;
  reg        [17:0]   img_reg_array_58_60_real;
  reg        [17:0]   img_reg_array_58_60_imag;
  reg        [17:0]   img_reg_array_58_61_real;
  reg        [17:0]   img_reg_array_58_61_imag;
  reg        [17:0]   img_reg_array_58_62_real;
  reg        [17:0]   img_reg_array_58_62_imag;
  reg        [17:0]   img_reg_array_58_63_real;
  reg        [17:0]   img_reg_array_58_63_imag;
  reg        [17:0]   img_reg_array_59_0_real;
  reg        [17:0]   img_reg_array_59_0_imag;
  reg        [17:0]   img_reg_array_59_1_real;
  reg        [17:0]   img_reg_array_59_1_imag;
  reg        [17:0]   img_reg_array_59_2_real;
  reg        [17:0]   img_reg_array_59_2_imag;
  reg        [17:0]   img_reg_array_59_3_real;
  reg        [17:0]   img_reg_array_59_3_imag;
  reg        [17:0]   img_reg_array_59_4_real;
  reg        [17:0]   img_reg_array_59_4_imag;
  reg        [17:0]   img_reg_array_59_5_real;
  reg        [17:0]   img_reg_array_59_5_imag;
  reg        [17:0]   img_reg_array_59_6_real;
  reg        [17:0]   img_reg_array_59_6_imag;
  reg        [17:0]   img_reg_array_59_7_real;
  reg        [17:0]   img_reg_array_59_7_imag;
  reg        [17:0]   img_reg_array_59_8_real;
  reg        [17:0]   img_reg_array_59_8_imag;
  reg        [17:0]   img_reg_array_59_9_real;
  reg        [17:0]   img_reg_array_59_9_imag;
  reg        [17:0]   img_reg_array_59_10_real;
  reg        [17:0]   img_reg_array_59_10_imag;
  reg        [17:0]   img_reg_array_59_11_real;
  reg        [17:0]   img_reg_array_59_11_imag;
  reg        [17:0]   img_reg_array_59_12_real;
  reg        [17:0]   img_reg_array_59_12_imag;
  reg        [17:0]   img_reg_array_59_13_real;
  reg        [17:0]   img_reg_array_59_13_imag;
  reg        [17:0]   img_reg_array_59_14_real;
  reg        [17:0]   img_reg_array_59_14_imag;
  reg        [17:0]   img_reg_array_59_15_real;
  reg        [17:0]   img_reg_array_59_15_imag;
  reg        [17:0]   img_reg_array_59_16_real;
  reg        [17:0]   img_reg_array_59_16_imag;
  reg        [17:0]   img_reg_array_59_17_real;
  reg        [17:0]   img_reg_array_59_17_imag;
  reg        [17:0]   img_reg_array_59_18_real;
  reg        [17:0]   img_reg_array_59_18_imag;
  reg        [17:0]   img_reg_array_59_19_real;
  reg        [17:0]   img_reg_array_59_19_imag;
  reg        [17:0]   img_reg_array_59_20_real;
  reg        [17:0]   img_reg_array_59_20_imag;
  reg        [17:0]   img_reg_array_59_21_real;
  reg        [17:0]   img_reg_array_59_21_imag;
  reg        [17:0]   img_reg_array_59_22_real;
  reg        [17:0]   img_reg_array_59_22_imag;
  reg        [17:0]   img_reg_array_59_23_real;
  reg        [17:0]   img_reg_array_59_23_imag;
  reg        [17:0]   img_reg_array_59_24_real;
  reg        [17:0]   img_reg_array_59_24_imag;
  reg        [17:0]   img_reg_array_59_25_real;
  reg        [17:0]   img_reg_array_59_25_imag;
  reg        [17:0]   img_reg_array_59_26_real;
  reg        [17:0]   img_reg_array_59_26_imag;
  reg        [17:0]   img_reg_array_59_27_real;
  reg        [17:0]   img_reg_array_59_27_imag;
  reg        [17:0]   img_reg_array_59_28_real;
  reg        [17:0]   img_reg_array_59_28_imag;
  reg        [17:0]   img_reg_array_59_29_real;
  reg        [17:0]   img_reg_array_59_29_imag;
  reg        [17:0]   img_reg_array_59_30_real;
  reg        [17:0]   img_reg_array_59_30_imag;
  reg        [17:0]   img_reg_array_59_31_real;
  reg        [17:0]   img_reg_array_59_31_imag;
  reg        [17:0]   img_reg_array_59_32_real;
  reg        [17:0]   img_reg_array_59_32_imag;
  reg        [17:0]   img_reg_array_59_33_real;
  reg        [17:0]   img_reg_array_59_33_imag;
  reg        [17:0]   img_reg_array_59_34_real;
  reg        [17:0]   img_reg_array_59_34_imag;
  reg        [17:0]   img_reg_array_59_35_real;
  reg        [17:0]   img_reg_array_59_35_imag;
  reg        [17:0]   img_reg_array_59_36_real;
  reg        [17:0]   img_reg_array_59_36_imag;
  reg        [17:0]   img_reg_array_59_37_real;
  reg        [17:0]   img_reg_array_59_37_imag;
  reg        [17:0]   img_reg_array_59_38_real;
  reg        [17:0]   img_reg_array_59_38_imag;
  reg        [17:0]   img_reg_array_59_39_real;
  reg        [17:0]   img_reg_array_59_39_imag;
  reg        [17:0]   img_reg_array_59_40_real;
  reg        [17:0]   img_reg_array_59_40_imag;
  reg        [17:0]   img_reg_array_59_41_real;
  reg        [17:0]   img_reg_array_59_41_imag;
  reg        [17:0]   img_reg_array_59_42_real;
  reg        [17:0]   img_reg_array_59_42_imag;
  reg        [17:0]   img_reg_array_59_43_real;
  reg        [17:0]   img_reg_array_59_43_imag;
  reg        [17:0]   img_reg_array_59_44_real;
  reg        [17:0]   img_reg_array_59_44_imag;
  reg        [17:0]   img_reg_array_59_45_real;
  reg        [17:0]   img_reg_array_59_45_imag;
  reg        [17:0]   img_reg_array_59_46_real;
  reg        [17:0]   img_reg_array_59_46_imag;
  reg        [17:0]   img_reg_array_59_47_real;
  reg        [17:0]   img_reg_array_59_47_imag;
  reg        [17:0]   img_reg_array_59_48_real;
  reg        [17:0]   img_reg_array_59_48_imag;
  reg        [17:0]   img_reg_array_59_49_real;
  reg        [17:0]   img_reg_array_59_49_imag;
  reg        [17:0]   img_reg_array_59_50_real;
  reg        [17:0]   img_reg_array_59_50_imag;
  reg        [17:0]   img_reg_array_59_51_real;
  reg        [17:0]   img_reg_array_59_51_imag;
  reg        [17:0]   img_reg_array_59_52_real;
  reg        [17:0]   img_reg_array_59_52_imag;
  reg        [17:0]   img_reg_array_59_53_real;
  reg        [17:0]   img_reg_array_59_53_imag;
  reg        [17:0]   img_reg_array_59_54_real;
  reg        [17:0]   img_reg_array_59_54_imag;
  reg        [17:0]   img_reg_array_59_55_real;
  reg        [17:0]   img_reg_array_59_55_imag;
  reg        [17:0]   img_reg_array_59_56_real;
  reg        [17:0]   img_reg_array_59_56_imag;
  reg        [17:0]   img_reg_array_59_57_real;
  reg        [17:0]   img_reg_array_59_57_imag;
  reg        [17:0]   img_reg_array_59_58_real;
  reg        [17:0]   img_reg_array_59_58_imag;
  reg        [17:0]   img_reg_array_59_59_real;
  reg        [17:0]   img_reg_array_59_59_imag;
  reg        [17:0]   img_reg_array_59_60_real;
  reg        [17:0]   img_reg_array_59_60_imag;
  reg        [17:0]   img_reg_array_59_61_real;
  reg        [17:0]   img_reg_array_59_61_imag;
  reg        [17:0]   img_reg_array_59_62_real;
  reg        [17:0]   img_reg_array_59_62_imag;
  reg        [17:0]   img_reg_array_59_63_real;
  reg        [17:0]   img_reg_array_59_63_imag;
  reg        [17:0]   img_reg_array_60_0_real;
  reg        [17:0]   img_reg_array_60_0_imag;
  reg        [17:0]   img_reg_array_60_1_real;
  reg        [17:0]   img_reg_array_60_1_imag;
  reg        [17:0]   img_reg_array_60_2_real;
  reg        [17:0]   img_reg_array_60_2_imag;
  reg        [17:0]   img_reg_array_60_3_real;
  reg        [17:0]   img_reg_array_60_3_imag;
  reg        [17:0]   img_reg_array_60_4_real;
  reg        [17:0]   img_reg_array_60_4_imag;
  reg        [17:0]   img_reg_array_60_5_real;
  reg        [17:0]   img_reg_array_60_5_imag;
  reg        [17:0]   img_reg_array_60_6_real;
  reg        [17:0]   img_reg_array_60_6_imag;
  reg        [17:0]   img_reg_array_60_7_real;
  reg        [17:0]   img_reg_array_60_7_imag;
  reg        [17:0]   img_reg_array_60_8_real;
  reg        [17:0]   img_reg_array_60_8_imag;
  reg        [17:0]   img_reg_array_60_9_real;
  reg        [17:0]   img_reg_array_60_9_imag;
  reg        [17:0]   img_reg_array_60_10_real;
  reg        [17:0]   img_reg_array_60_10_imag;
  reg        [17:0]   img_reg_array_60_11_real;
  reg        [17:0]   img_reg_array_60_11_imag;
  reg        [17:0]   img_reg_array_60_12_real;
  reg        [17:0]   img_reg_array_60_12_imag;
  reg        [17:0]   img_reg_array_60_13_real;
  reg        [17:0]   img_reg_array_60_13_imag;
  reg        [17:0]   img_reg_array_60_14_real;
  reg        [17:0]   img_reg_array_60_14_imag;
  reg        [17:0]   img_reg_array_60_15_real;
  reg        [17:0]   img_reg_array_60_15_imag;
  reg        [17:0]   img_reg_array_60_16_real;
  reg        [17:0]   img_reg_array_60_16_imag;
  reg        [17:0]   img_reg_array_60_17_real;
  reg        [17:0]   img_reg_array_60_17_imag;
  reg        [17:0]   img_reg_array_60_18_real;
  reg        [17:0]   img_reg_array_60_18_imag;
  reg        [17:0]   img_reg_array_60_19_real;
  reg        [17:0]   img_reg_array_60_19_imag;
  reg        [17:0]   img_reg_array_60_20_real;
  reg        [17:0]   img_reg_array_60_20_imag;
  reg        [17:0]   img_reg_array_60_21_real;
  reg        [17:0]   img_reg_array_60_21_imag;
  reg        [17:0]   img_reg_array_60_22_real;
  reg        [17:0]   img_reg_array_60_22_imag;
  reg        [17:0]   img_reg_array_60_23_real;
  reg        [17:0]   img_reg_array_60_23_imag;
  reg        [17:0]   img_reg_array_60_24_real;
  reg        [17:0]   img_reg_array_60_24_imag;
  reg        [17:0]   img_reg_array_60_25_real;
  reg        [17:0]   img_reg_array_60_25_imag;
  reg        [17:0]   img_reg_array_60_26_real;
  reg        [17:0]   img_reg_array_60_26_imag;
  reg        [17:0]   img_reg_array_60_27_real;
  reg        [17:0]   img_reg_array_60_27_imag;
  reg        [17:0]   img_reg_array_60_28_real;
  reg        [17:0]   img_reg_array_60_28_imag;
  reg        [17:0]   img_reg_array_60_29_real;
  reg        [17:0]   img_reg_array_60_29_imag;
  reg        [17:0]   img_reg_array_60_30_real;
  reg        [17:0]   img_reg_array_60_30_imag;
  reg        [17:0]   img_reg_array_60_31_real;
  reg        [17:0]   img_reg_array_60_31_imag;
  reg        [17:0]   img_reg_array_60_32_real;
  reg        [17:0]   img_reg_array_60_32_imag;
  reg        [17:0]   img_reg_array_60_33_real;
  reg        [17:0]   img_reg_array_60_33_imag;
  reg        [17:0]   img_reg_array_60_34_real;
  reg        [17:0]   img_reg_array_60_34_imag;
  reg        [17:0]   img_reg_array_60_35_real;
  reg        [17:0]   img_reg_array_60_35_imag;
  reg        [17:0]   img_reg_array_60_36_real;
  reg        [17:0]   img_reg_array_60_36_imag;
  reg        [17:0]   img_reg_array_60_37_real;
  reg        [17:0]   img_reg_array_60_37_imag;
  reg        [17:0]   img_reg_array_60_38_real;
  reg        [17:0]   img_reg_array_60_38_imag;
  reg        [17:0]   img_reg_array_60_39_real;
  reg        [17:0]   img_reg_array_60_39_imag;
  reg        [17:0]   img_reg_array_60_40_real;
  reg        [17:0]   img_reg_array_60_40_imag;
  reg        [17:0]   img_reg_array_60_41_real;
  reg        [17:0]   img_reg_array_60_41_imag;
  reg        [17:0]   img_reg_array_60_42_real;
  reg        [17:0]   img_reg_array_60_42_imag;
  reg        [17:0]   img_reg_array_60_43_real;
  reg        [17:0]   img_reg_array_60_43_imag;
  reg        [17:0]   img_reg_array_60_44_real;
  reg        [17:0]   img_reg_array_60_44_imag;
  reg        [17:0]   img_reg_array_60_45_real;
  reg        [17:0]   img_reg_array_60_45_imag;
  reg        [17:0]   img_reg_array_60_46_real;
  reg        [17:0]   img_reg_array_60_46_imag;
  reg        [17:0]   img_reg_array_60_47_real;
  reg        [17:0]   img_reg_array_60_47_imag;
  reg        [17:0]   img_reg_array_60_48_real;
  reg        [17:0]   img_reg_array_60_48_imag;
  reg        [17:0]   img_reg_array_60_49_real;
  reg        [17:0]   img_reg_array_60_49_imag;
  reg        [17:0]   img_reg_array_60_50_real;
  reg        [17:0]   img_reg_array_60_50_imag;
  reg        [17:0]   img_reg_array_60_51_real;
  reg        [17:0]   img_reg_array_60_51_imag;
  reg        [17:0]   img_reg_array_60_52_real;
  reg        [17:0]   img_reg_array_60_52_imag;
  reg        [17:0]   img_reg_array_60_53_real;
  reg        [17:0]   img_reg_array_60_53_imag;
  reg        [17:0]   img_reg_array_60_54_real;
  reg        [17:0]   img_reg_array_60_54_imag;
  reg        [17:0]   img_reg_array_60_55_real;
  reg        [17:0]   img_reg_array_60_55_imag;
  reg        [17:0]   img_reg_array_60_56_real;
  reg        [17:0]   img_reg_array_60_56_imag;
  reg        [17:0]   img_reg_array_60_57_real;
  reg        [17:0]   img_reg_array_60_57_imag;
  reg        [17:0]   img_reg_array_60_58_real;
  reg        [17:0]   img_reg_array_60_58_imag;
  reg        [17:0]   img_reg_array_60_59_real;
  reg        [17:0]   img_reg_array_60_59_imag;
  reg        [17:0]   img_reg_array_60_60_real;
  reg        [17:0]   img_reg_array_60_60_imag;
  reg        [17:0]   img_reg_array_60_61_real;
  reg        [17:0]   img_reg_array_60_61_imag;
  reg        [17:0]   img_reg_array_60_62_real;
  reg        [17:0]   img_reg_array_60_62_imag;
  reg        [17:0]   img_reg_array_60_63_real;
  reg        [17:0]   img_reg_array_60_63_imag;
  reg        [17:0]   img_reg_array_61_0_real;
  reg        [17:0]   img_reg_array_61_0_imag;
  reg        [17:0]   img_reg_array_61_1_real;
  reg        [17:0]   img_reg_array_61_1_imag;
  reg        [17:0]   img_reg_array_61_2_real;
  reg        [17:0]   img_reg_array_61_2_imag;
  reg        [17:0]   img_reg_array_61_3_real;
  reg        [17:0]   img_reg_array_61_3_imag;
  reg        [17:0]   img_reg_array_61_4_real;
  reg        [17:0]   img_reg_array_61_4_imag;
  reg        [17:0]   img_reg_array_61_5_real;
  reg        [17:0]   img_reg_array_61_5_imag;
  reg        [17:0]   img_reg_array_61_6_real;
  reg        [17:0]   img_reg_array_61_6_imag;
  reg        [17:0]   img_reg_array_61_7_real;
  reg        [17:0]   img_reg_array_61_7_imag;
  reg        [17:0]   img_reg_array_61_8_real;
  reg        [17:0]   img_reg_array_61_8_imag;
  reg        [17:0]   img_reg_array_61_9_real;
  reg        [17:0]   img_reg_array_61_9_imag;
  reg        [17:0]   img_reg_array_61_10_real;
  reg        [17:0]   img_reg_array_61_10_imag;
  reg        [17:0]   img_reg_array_61_11_real;
  reg        [17:0]   img_reg_array_61_11_imag;
  reg        [17:0]   img_reg_array_61_12_real;
  reg        [17:0]   img_reg_array_61_12_imag;
  reg        [17:0]   img_reg_array_61_13_real;
  reg        [17:0]   img_reg_array_61_13_imag;
  reg        [17:0]   img_reg_array_61_14_real;
  reg        [17:0]   img_reg_array_61_14_imag;
  reg        [17:0]   img_reg_array_61_15_real;
  reg        [17:0]   img_reg_array_61_15_imag;
  reg        [17:0]   img_reg_array_61_16_real;
  reg        [17:0]   img_reg_array_61_16_imag;
  reg        [17:0]   img_reg_array_61_17_real;
  reg        [17:0]   img_reg_array_61_17_imag;
  reg        [17:0]   img_reg_array_61_18_real;
  reg        [17:0]   img_reg_array_61_18_imag;
  reg        [17:0]   img_reg_array_61_19_real;
  reg        [17:0]   img_reg_array_61_19_imag;
  reg        [17:0]   img_reg_array_61_20_real;
  reg        [17:0]   img_reg_array_61_20_imag;
  reg        [17:0]   img_reg_array_61_21_real;
  reg        [17:0]   img_reg_array_61_21_imag;
  reg        [17:0]   img_reg_array_61_22_real;
  reg        [17:0]   img_reg_array_61_22_imag;
  reg        [17:0]   img_reg_array_61_23_real;
  reg        [17:0]   img_reg_array_61_23_imag;
  reg        [17:0]   img_reg_array_61_24_real;
  reg        [17:0]   img_reg_array_61_24_imag;
  reg        [17:0]   img_reg_array_61_25_real;
  reg        [17:0]   img_reg_array_61_25_imag;
  reg        [17:0]   img_reg_array_61_26_real;
  reg        [17:0]   img_reg_array_61_26_imag;
  reg        [17:0]   img_reg_array_61_27_real;
  reg        [17:0]   img_reg_array_61_27_imag;
  reg        [17:0]   img_reg_array_61_28_real;
  reg        [17:0]   img_reg_array_61_28_imag;
  reg        [17:0]   img_reg_array_61_29_real;
  reg        [17:0]   img_reg_array_61_29_imag;
  reg        [17:0]   img_reg_array_61_30_real;
  reg        [17:0]   img_reg_array_61_30_imag;
  reg        [17:0]   img_reg_array_61_31_real;
  reg        [17:0]   img_reg_array_61_31_imag;
  reg        [17:0]   img_reg_array_61_32_real;
  reg        [17:0]   img_reg_array_61_32_imag;
  reg        [17:0]   img_reg_array_61_33_real;
  reg        [17:0]   img_reg_array_61_33_imag;
  reg        [17:0]   img_reg_array_61_34_real;
  reg        [17:0]   img_reg_array_61_34_imag;
  reg        [17:0]   img_reg_array_61_35_real;
  reg        [17:0]   img_reg_array_61_35_imag;
  reg        [17:0]   img_reg_array_61_36_real;
  reg        [17:0]   img_reg_array_61_36_imag;
  reg        [17:0]   img_reg_array_61_37_real;
  reg        [17:0]   img_reg_array_61_37_imag;
  reg        [17:0]   img_reg_array_61_38_real;
  reg        [17:0]   img_reg_array_61_38_imag;
  reg        [17:0]   img_reg_array_61_39_real;
  reg        [17:0]   img_reg_array_61_39_imag;
  reg        [17:0]   img_reg_array_61_40_real;
  reg        [17:0]   img_reg_array_61_40_imag;
  reg        [17:0]   img_reg_array_61_41_real;
  reg        [17:0]   img_reg_array_61_41_imag;
  reg        [17:0]   img_reg_array_61_42_real;
  reg        [17:0]   img_reg_array_61_42_imag;
  reg        [17:0]   img_reg_array_61_43_real;
  reg        [17:0]   img_reg_array_61_43_imag;
  reg        [17:0]   img_reg_array_61_44_real;
  reg        [17:0]   img_reg_array_61_44_imag;
  reg        [17:0]   img_reg_array_61_45_real;
  reg        [17:0]   img_reg_array_61_45_imag;
  reg        [17:0]   img_reg_array_61_46_real;
  reg        [17:0]   img_reg_array_61_46_imag;
  reg        [17:0]   img_reg_array_61_47_real;
  reg        [17:0]   img_reg_array_61_47_imag;
  reg        [17:0]   img_reg_array_61_48_real;
  reg        [17:0]   img_reg_array_61_48_imag;
  reg        [17:0]   img_reg_array_61_49_real;
  reg        [17:0]   img_reg_array_61_49_imag;
  reg        [17:0]   img_reg_array_61_50_real;
  reg        [17:0]   img_reg_array_61_50_imag;
  reg        [17:0]   img_reg_array_61_51_real;
  reg        [17:0]   img_reg_array_61_51_imag;
  reg        [17:0]   img_reg_array_61_52_real;
  reg        [17:0]   img_reg_array_61_52_imag;
  reg        [17:0]   img_reg_array_61_53_real;
  reg        [17:0]   img_reg_array_61_53_imag;
  reg        [17:0]   img_reg_array_61_54_real;
  reg        [17:0]   img_reg_array_61_54_imag;
  reg        [17:0]   img_reg_array_61_55_real;
  reg        [17:0]   img_reg_array_61_55_imag;
  reg        [17:0]   img_reg_array_61_56_real;
  reg        [17:0]   img_reg_array_61_56_imag;
  reg        [17:0]   img_reg_array_61_57_real;
  reg        [17:0]   img_reg_array_61_57_imag;
  reg        [17:0]   img_reg_array_61_58_real;
  reg        [17:0]   img_reg_array_61_58_imag;
  reg        [17:0]   img_reg_array_61_59_real;
  reg        [17:0]   img_reg_array_61_59_imag;
  reg        [17:0]   img_reg_array_61_60_real;
  reg        [17:0]   img_reg_array_61_60_imag;
  reg        [17:0]   img_reg_array_61_61_real;
  reg        [17:0]   img_reg_array_61_61_imag;
  reg        [17:0]   img_reg_array_61_62_real;
  reg        [17:0]   img_reg_array_61_62_imag;
  reg        [17:0]   img_reg_array_61_63_real;
  reg        [17:0]   img_reg_array_61_63_imag;
  reg        [17:0]   img_reg_array_62_0_real;
  reg        [17:0]   img_reg_array_62_0_imag;
  reg        [17:0]   img_reg_array_62_1_real;
  reg        [17:0]   img_reg_array_62_1_imag;
  reg        [17:0]   img_reg_array_62_2_real;
  reg        [17:0]   img_reg_array_62_2_imag;
  reg        [17:0]   img_reg_array_62_3_real;
  reg        [17:0]   img_reg_array_62_3_imag;
  reg        [17:0]   img_reg_array_62_4_real;
  reg        [17:0]   img_reg_array_62_4_imag;
  reg        [17:0]   img_reg_array_62_5_real;
  reg        [17:0]   img_reg_array_62_5_imag;
  reg        [17:0]   img_reg_array_62_6_real;
  reg        [17:0]   img_reg_array_62_6_imag;
  reg        [17:0]   img_reg_array_62_7_real;
  reg        [17:0]   img_reg_array_62_7_imag;
  reg        [17:0]   img_reg_array_62_8_real;
  reg        [17:0]   img_reg_array_62_8_imag;
  reg        [17:0]   img_reg_array_62_9_real;
  reg        [17:0]   img_reg_array_62_9_imag;
  reg        [17:0]   img_reg_array_62_10_real;
  reg        [17:0]   img_reg_array_62_10_imag;
  reg        [17:0]   img_reg_array_62_11_real;
  reg        [17:0]   img_reg_array_62_11_imag;
  reg        [17:0]   img_reg_array_62_12_real;
  reg        [17:0]   img_reg_array_62_12_imag;
  reg        [17:0]   img_reg_array_62_13_real;
  reg        [17:0]   img_reg_array_62_13_imag;
  reg        [17:0]   img_reg_array_62_14_real;
  reg        [17:0]   img_reg_array_62_14_imag;
  reg        [17:0]   img_reg_array_62_15_real;
  reg        [17:0]   img_reg_array_62_15_imag;
  reg        [17:0]   img_reg_array_62_16_real;
  reg        [17:0]   img_reg_array_62_16_imag;
  reg        [17:0]   img_reg_array_62_17_real;
  reg        [17:0]   img_reg_array_62_17_imag;
  reg        [17:0]   img_reg_array_62_18_real;
  reg        [17:0]   img_reg_array_62_18_imag;
  reg        [17:0]   img_reg_array_62_19_real;
  reg        [17:0]   img_reg_array_62_19_imag;
  reg        [17:0]   img_reg_array_62_20_real;
  reg        [17:0]   img_reg_array_62_20_imag;
  reg        [17:0]   img_reg_array_62_21_real;
  reg        [17:0]   img_reg_array_62_21_imag;
  reg        [17:0]   img_reg_array_62_22_real;
  reg        [17:0]   img_reg_array_62_22_imag;
  reg        [17:0]   img_reg_array_62_23_real;
  reg        [17:0]   img_reg_array_62_23_imag;
  reg        [17:0]   img_reg_array_62_24_real;
  reg        [17:0]   img_reg_array_62_24_imag;
  reg        [17:0]   img_reg_array_62_25_real;
  reg        [17:0]   img_reg_array_62_25_imag;
  reg        [17:0]   img_reg_array_62_26_real;
  reg        [17:0]   img_reg_array_62_26_imag;
  reg        [17:0]   img_reg_array_62_27_real;
  reg        [17:0]   img_reg_array_62_27_imag;
  reg        [17:0]   img_reg_array_62_28_real;
  reg        [17:0]   img_reg_array_62_28_imag;
  reg        [17:0]   img_reg_array_62_29_real;
  reg        [17:0]   img_reg_array_62_29_imag;
  reg        [17:0]   img_reg_array_62_30_real;
  reg        [17:0]   img_reg_array_62_30_imag;
  reg        [17:0]   img_reg_array_62_31_real;
  reg        [17:0]   img_reg_array_62_31_imag;
  reg        [17:0]   img_reg_array_62_32_real;
  reg        [17:0]   img_reg_array_62_32_imag;
  reg        [17:0]   img_reg_array_62_33_real;
  reg        [17:0]   img_reg_array_62_33_imag;
  reg        [17:0]   img_reg_array_62_34_real;
  reg        [17:0]   img_reg_array_62_34_imag;
  reg        [17:0]   img_reg_array_62_35_real;
  reg        [17:0]   img_reg_array_62_35_imag;
  reg        [17:0]   img_reg_array_62_36_real;
  reg        [17:0]   img_reg_array_62_36_imag;
  reg        [17:0]   img_reg_array_62_37_real;
  reg        [17:0]   img_reg_array_62_37_imag;
  reg        [17:0]   img_reg_array_62_38_real;
  reg        [17:0]   img_reg_array_62_38_imag;
  reg        [17:0]   img_reg_array_62_39_real;
  reg        [17:0]   img_reg_array_62_39_imag;
  reg        [17:0]   img_reg_array_62_40_real;
  reg        [17:0]   img_reg_array_62_40_imag;
  reg        [17:0]   img_reg_array_62_41_real;
  reg        [17:0]   img_reg_array_62_41_imag;
  reg        [17:0]   img_reg_array_62_42_real;
  reg        [17:0]   img_reg_array_62_42_imag;
  reg        [17:0]   img_reg_array_62_43_real;
  reg        [17:0]   img_reg_array_62_43_imag;
  reg        [17:0]   img_reg_array_62_44_real;
  reg        [17:0]   img_reg_array_62_44_imag;
  reg        [17:0]   img_reg_array_62_45_real;
  reg        [17:0]   img_reg_array_62_45_imag;
  reg        [17:0]   img_reg_array_62_46_real;
  reg        [17:0]   img_reg_array_62_46_imag;
  reg        [17:0]   img_reg_array_62_47_real;
  reg        [17:0]   img_reg_array_62_47_imag;
  reg        [17:0]   img_reg_array_62_48_real;
  reg        [17:0]   img_reg_array_62_48_imag;
  reg        [17:0]   img_reg_array_62_49_real;
  reg        [17:0]   img_reg_array_62_49_imag;
  reg        [17:0]   img_reg_array_62_50_real;
  reg        [17:0]   img_reg_array_62_50_imag;
  reg        [17:0]   img_reg_array_62_51_real;
  reg        [17:0]   img_reg_array_62_51_imag;
  reg        [17:0]   img_reg_array_62_52_real;
  reg        [17:0]   img_reg_array_62_52_imag;
  reg        [17:0]   img_reg_array_62_53_real;
  reg        [17:0]   img_reg_array_62_53_imag;
  reg        [17:0]   img_reg_array_62_54_real;
  reg        [17:0]   img_reg_array_62_54_imag;
  reg        [17:0]   img_reg_array_62_55_real;
  reg        [17:0]   img_reg_array_62_55_imag;
  reg        [17:0]   img_reg_array_62_56_real;
  reg        [17:0]   img_reg_array_62_56_imag;
  reg        [17:0]   img_reg_array_62_57_real;
  reg        [17:0]   img_reg_array_62_57_imag;
  reg        [17:0]   img_reg_array_62_58_real;
  reg        [17:0]   img_reg_array_62_58_imag;
  reg        [17:0]   img_reg_array_62_59_real;
  reg        [17:0]   img_reg_array_62_59_imag;
  reg        [17:0]   img_reg_array_62_60_real;
  reg        [17:0]   img_reg_array_62_60_imag;
  reg        [17:0]   img_reg_array_62_61_real;
  reg        [17:0]   img_reg_array_62_61_imag;
  reg        [17:0]   img_reg_array_62_62_real;
  reg        [17:0]   img_reg_array_62_62_imag;
  reg        [17:0]   img_reg_array_62_63_real;
  reg        [17:0]   img_reg_array_62_63_imag;
  reg        [17:0]   img_reg_array_63_0_real;
  reg        [17:0]   img_reg_array_63_0_imag;
  reg        [17:0]   img_reg_array_63_1_real;
  reg        [17:0]   img_reg_array_63_1_imag;
  reg        [17:0]   img_reg_array_63_2_real;
  reg        [17:0]   img_reg_array_63_2_imag;
  reg        [17:0]   img_reg_array_63_3_real;
  reg        [17:0]   img_reg_array_63_3_imag;
  reg        [17:0]   img_reg_array_63_4_real;
  reg        [17:0]   img_reg_array_63_4_imag;
  reg        [17:0]   img_reg_array_63_5_real;
  reg        [17:0]   img_reg_array_63_5_imag;
  reg        [17:0]   img_reg_array_63_6_real;
  reg        [17:0]   img_reg_array_63_6_imag;
  reg        [17:0]   img_reg_array_63_7_real;
  reg        [17:0]   img_reg_array_63_7_imag;
  reg        [17:0]   img_reg_array_63_8_real;
  reg        [17:0]   img_reg_array_63_8_imag;
  reg        [17:0]   img_reg_array_63_9_real;
  reg        [17:0]   img_reg_array_63_9_imag;
  reg        [17:0]   img_reg_array_63_10_real;
  reg        [17:0]   img_reg_array_63_10_imag;
  reg        [17:0]   img_reg_array_63_11_real;
  reg        [17:0]   img_reg_array_63_11_imag;
  reg        [17:0]   img_reg_array_63_12_real;
  reg        [17:0]   img_reg_array_63_12_imag;
  reg        [17:0]   img_reg_array_63_13_real;
  reg        [17:0]   img_reg_array_63_13_imag;
  reg        [17:0]   img_reg_array_63_14_real;
  reg        [17:0]   img_reg_array_63_14_imag;
  reg        [17:0]   img_reg_array_63_15_real;
  reg        [17:0]   img_reg_array_63_15_imag;
  reg        [17:0]   img_reg_array_63_16_real;
  reg        [17:0]   img_reg_array_63_16_imag;
  reg        [17:0]   img_reg_array_63_17_real;
  reg        [17:0]   img_reg_array_63_17_imag;
  reg        [17:0]   img_reg_array_63_18_real;
  reg        [17:0]   img_reg_array_63_18_imag;
  reg        [17:0]   img_reg_array_63_19_real;
  reg        [17:0]   img_reg_array_63_19_imag;
  reg        [17:0]   img_reg_array_63_20_real;
  reg        [17:0]   img_reg_array_63_20_imag;
  reg        [17:0]   img_reg_array_63_21_real;
  reg        [17:0]   img_reg_array_63_21_imag;
  reg        [17:0]   img_reg_array_63_22_real;
  reg        [17:0]   img_reg_array_63_22_imag;
  reg        [17:0]   img_reg_array_63_23_real;
  reg        [17:0]   img_reg_array_63_23_imag;
  reg        [17:0]   img_reg_array_63_24_real;
  reg        [17:0]   img_reg_array_63_24_imag;
  reg        [17:0]   img_reg_array_63_25_real;
  reg        [17:0]   img_reg_array_63_25_imag;
  reg        [17:0]   img_reg_array_63_26_real;
  reg        [17:0]   img_reg_array_63_26_imag;
  reg        [17:0]   img_reg_array_63_27_real;
  reg        [17:0]   img_reg_array_63_27_imag;
  reg        [17:0]   img_reg_array_63_28_real;
  reg        [17:0]   img_reg_array_63_28_imag;
  reg        [17:0]   img_reg_array_63_29_real;
  reg        [17:0]   img_reg_array_63_29_imag;
  reg        [17:0]   img_reg_array_63_30_real;
  reg        [17:0]   img_reg_array_63_30_imag;
  reg        [17:0]   img_reg_array_63_31_real;
  reg        [17:0]   img_reg_array_63_31_imag;
  reg        [17:0]   img_reg_array_63_32_real;
  reg        [17:0]   img_reg_array_63_32_imag;
  reg        [17:0]   img_reg_array_63_33_real;
  reg        [17:0]   img_reg_array_63_33_imag;
  reg        [17:0]   img_reg_array_63_34_real;
  reg        [17:0]   img_reg_array_63_34_imag;
  reg        [17:0]   img_reg_array_63_35_real;
  reg        [17:0]   img_reg_array_63_35_imag;
  reg        [17:0]   img_reg_array_63_36_real;
  reg        [17:0]   img_reg_array_63_36_imag;
  reg        [17:0]   img_reg_array_63_37_real;
  reg        [17:0]   img_reg_array_63_37_imag;
  reg        [17:0]   img_reg_array_63_38_real;
  reg        [17:0]   img_reg_array_63_38_imag;
  reg        [17:0]   img_reg_array_63_39_real;
  reg        [17:0]   img_reg_array_63_39_imag;
  reg        [17:0]   img_reg_array_63_40_real;
  reg        [17:0]   img_reg_array_63_40_imag;
  reg        [17:0]   img_reg_array_63_41_real;
  reg        [17:0]   img_reg_array_63_41_imag;
  reg        [17:0]   img_reg_array_63_42_real;
  reg        [17:0]   img_reg_array_63_42_imag;
  reg        [17:0]   img_reg_array_63_43_real;
  reg        [17:0]   img_reg_array_63_43_imag;
  reg        [17:0]   img_reg_array_63_44_real;
  reg        [17:0]   img_reg_array_63_44_imag;
  reg        [17:0]   img_reg_array_63_45_real;
  reg        [17:0]   img_reg_array_63_45_imag;
  reg        [17:0]   img_reg_array_63_46_real;
  reg        [17:0]   img_reg_array_63_46_imag;
  reg        [17:0]   img_reg_array_63_47_real;
  reg        [17:0]   img_reg_array_63_47_imag;
  reg        [17:0]   img_reg_array_63_48_real;
  reg        [17:0]   img_reg_array_63_48_imag;
  reg        [17:0]   img_reg_array_63_49_real;
  reg        [17:0]   img_reg_array_63_49_imag;
  reg        [17:0]   img_reg_array_63_50_real;
  reg        [17:0]   img_reg_array_63_50_imag;
  reg        [17:0]   img_reg_array_63_51_real;
  reg        [17:0]   img_reg_array_63_51_imag;
  reg        [17:0]   img_reg_array_63_52_real;
  reg        [17:0]   img_reg_array_63_52_imag;
  reg        [17:0]   img_reg_array_63_53_real;
  reg        [17:0]   img_reg_array_63_53_imag;
  reg        [17:0]   img_reg_array_63_54_real;
  reg        [17:0]   img_reg_array_63_54_imag;
  reg        [17:0]   img_reg_array_63_55_real;
  reg        [17:0]   img_reg_array_63_55_imag;
  reg        [17:0]   img_reg_array_63_56_real;
  reg        [17:0]   img_reg_array_63_56_imag;
  reg        [17:0]   img_reg_array_63_57_real;
  reg        [17:0]   img_reg_array_63_57_imag;
  reg        [17:0]   img_reg_array_63_58_real;
  reg        [17:0]   img_reg_array_63_58_imag;
  reg        [17:0]   img_reg_array_63_59_real;
  reg        [17:0]   img_reg_array_63_59_imag;
  reg        [17:0]   img_reg_array_63_60_real;
  reg        [17:0]   img_reg_array_63_60_imag;
  reg        [17:0]   img_reg_array_63_61_real;
  reg        [17:0]   img_reg_array_63_61_imag;
  reg        [17:0]   img_reg_array_63_62_real;
  reg        [17:0]   img_reg_array_63_62_imag;
  reg        [17:0]   img_reg_array_63_63_real;
  reg        [17:0]   img_reg_array_63_63_imag;
  reg                 row_addr_willIncrement;
  wire                row_addr_willClear;
  reg        [5:0]    row_addr_valueNext;
  reg        [5:0]    row_addr_value;
  wire                row_addr_willOverflowIfInc;
  wire                row_addr_willOverflow;
  wire       [63:0]   _zz_1;
  wire                _zz_2;
  wire                _zz_3;
  wire                _zz_4;
  wire                _zz_5;
  wire                _zz_6;
  wire                _zz_7;
  wire                _zz_8;
  wire                _zz_9;
  wire                _zz_10;
  wire                _zz_11;
  wire                _zz_12;
  wire                _zz_13;
  wire                _zz_14;
  wire                _zz_15;
  wire                _zz_16;
  wire                _zz_17;
  wire                _zz_18;
  wire                _zz_19;
  wire                _zz_20;
  wire                _zz_21;
  wire                _zz_22;
  wire                _zz_23;
  wire                _zz_24;
  wire                _zz_25;
  wire                _zz_26;
  wire                _zz_27;
  wire                _zz_28;
  wire                _zz_29;
  wire                _zz_30;
  wire                _zz_31;
  wire                _zz_32;
  wire                _zz_33;
  wire                _zz_34;
  wire                _zz_35;
  wire                _zz_36;
  wire                _zz_37;
  wire                _zz_38;
  wire                _zz_39;
  wire                _zz_40;
  wire                _zz_41;
  wire                _zz_42;
  wire                _zz_43;
  wire                _zz_44;
  wire                _zz_45;
  wire                _zz_46;
  wire                _zz_47;
  wire                _zz_48;
  wire                _zz_49;
  wire                _zz_50;
  wire                _zz_51;
  wire                _zz_52;
  wire                _zz_53;
  wire                _zz_54;
  wire                _zz_55;
  wire                _zz_56;
  wire                _zz_57;
  wire                _zz_58;
  wire                _zz_59;
  wire                _zz_60;
  wire                _zz_61;
  wire                _zz_62;
  wire                _zz_63;
  wire                _zz_64;
  wire                _zz_65;
  wire       [17:0]   _zz_66;
  wire       [17:0]   _zz_67;
  wire       [17:0]   _zz_68;
  wire       [17:0]   _zz_69;
  wire       [17:0]   _zz_70;
  wire       [17:0]   _zz_71;
  wire       [17:0]   _zz_72;
  wire       [17:0]   _zz_73;
  wire       [17:0]   _zz_74;
  wire       [17:0]   _zz_75;
  wire       [17:0]   _zz_76;
  wire       [17:0]   _zz_77;
  wire       [17:0]   _zz_78;
  wire       [17:0]   _zz_79;
  wire       [17:0]   _zz_80;
  wire       [17:0]   _zz_81;
  wire       [17:0]   _zz_82;
  wire       [17:0]   _zz_83;
  wire       [17:0]   _zz_84;
  wire       [17:0]   _zz_85;
  wire       [17:0]   _zz_86;
  wire       [17:0]   _zz_87;
  wire       [17:0]   _zz_88;
  wire       [17:0]   _zz_89;
  wire       [17:0]   _zz_90;
  wire       [17:0]   _zz_91;
  wire       [17:0]   _zz_92;
  wire       [17:0]   _zz_93;
  wire       [17:0]   _zz_94;
  wire       [17:0]   _zz_95;
  wire       [17:0]   _zz_96;
  wire       [17:0]   _zz_97;
  wire       [17:0]   _zz_98;
  wire       [17:0]   _zz_99;
  wire       [17:0]   _zz_100;
  wire       [17:0]   _zz_101;
  wire       [17:0]   _zz_102;
  wire       [17:0]   _zz_103;
  wire       [17:0]   _zz_104;
  wire       [17:0]   _zz_105;
  wire       [17:0]   _zz_106;
  wire       [17:0]   _zz_107;
  wire       [17:0]   _zz_108;
  wire       [17:0]   _zz_109;
  wire       [17:0]   _zz_110;
  wire       [17:0]   _zz_111;
  wire       [17:0]   _zz_112;
  wire       [17:0]   _zz_113;
  wire       [17:0]   _zz_114;
  wire       [17:0]   _zz_115;
  wire       [17:0]   _zz_116;
  wire       [17:0]   _zz_117;
  wire       [17:0]   _zz_118;
  wire       [17:0]   _zz_119;
  wire       [17:0]   _zz_120;
  wire       [17:0]   _zz_121;
  wire       [17:0]   _zz_122;
  wire       [17:0]   _zz_123;
  wire       [17:0]   _zz_124;
  wire       [17:0]   _zz_125;
  wire       [17:0]   _zz_126;
  wire       [17:0]   _zz_127;
  wire       [17:0]   _zz_128;
  wire       [17:0]   _zz_129;
  wire       [17:0]   _zz_130;
  wire       [17:0]   _zz_131;
  wire       [17:0]   _zz_132;
  wire       [17:0]   _zz_133;
  wire       [17:0]   _zz_134;
  wire       [17:0]   _zz_135;
  wire       [17:0]   _zz_136;
  wire       [17:0]   _zz_137;
  wire       [17:0]   _zz_138;
  wire       [17:0]   _zz_139;
  wire       [17:0]   _zz_140;
  wire       [17:0]   _zz_141;
  wire       [17:0]   _zz_142;
  wire       [17:0]   _zz_143;
  wire       [17:0]   _zz_144;
  wire       [17:0]   _zz_145;
  wire       [17:0]   _zz_146;
  wire       [17:0]   _zz_147;
  wire       [17:0]   _zz_148;
  wire       [17:0]   _zz_149;
  wire       [17:0]   _zz_150;
  wire       [17:0]   _zz_151;
  wire       [17:0]   _zz_152;
  wire       [17:0]   _zz_153;
  wire       [17:0]   _zz_154;
  wire       [17:0]   _zz_155;
  wire       [17:0]   _zz_156;
  wire       [17:0]   _zz_157;
  wire       [17:0]   _zz_158;
  wire       [17:0]   _zz_159;
  wire       [17:0]   _zz_160;
  wire       [17:0]   _zz_161;
  wire       [17:0]   _zz_162;
  wire       [17:0]   _zz_163;
  wire       [17:0]   _zz_164;
  wire       [17:0]   _zz_165;
  wire       [17:0]   _zz_166;
  wire       [17:0]   _zz_167;
  wire       [17:0]   _zz_168;
  wire       [17:0]   _zz_169;
  wire       [17:0]   _zz_170;
  wire       [17:0]   _zz_171;
  wire       [17:0]   _zz_172;
  wire       [17:0]   _zz_173;
  wire       [17:0]   _zz_174;
  wire       [17:0]   _zz_175;
  wire       [17:0]   _zz_176;
  wire       [17:0]   _zz_177;
  wire       [17:0]   _zz_178;
  wire       [17:0]   _zz_179;
  wire       [17:0]   _zz_180;
  wire       [17:0]   _zz_181;
  wire       [17:0]   _zz_182;
  wire       [17:0]   _zz_183;
  wire       [17:0]   _zz_184;
  wire       [17:0]   _zz_185;
  wire       [17:0]   _zz_186;
  wire       [17:0]   _zz_187;
  wire       [17:0]   _zz_188;
  wire       [17:0]   _zz_189;
  wire       [17:0]   _zz_190;
  wire       [17:0]   _zz_191;
  wire       [17:0]   _zz_192;
  wire       [17:0]   _zz_193;
  reg                 null_cnt_willIncrement;
  wire                null_cnt_willClear;
  reg        [5:0]    null_cnt_valueNext;
  reg        [5:0]    null_cnt_value;
  wire                null_cnt_willOverflowIfInc;
  wire                null_cnt_willOverflow;
  reg                 null_cond_period_minus_1;
  wire                null_cond_period;
  reg        [5:0]    col_addr;
  wire                fft_col_in_valid;
  wire       [17:0]   fft_col_in_payload_0_real;
  wire       [17:0]   fft_col_in_payload_0_imag;
  wire       [17:0]   fft_col_in_payload_1_real;
  wire       [17:0]   fft_col_in_payload_1_imag;
  wire       [17:0]   fft_col_in_payload_2_real;
  wire       [17:0]   fft_col_in_payload_2_imag;
  wire       [17:0]   fft_col_in_payload_3_real;
  wire       [17:0]   fft_col_in_payload_3_imag;
  wire       [17:0]   fft_col_in_payload_4_real;
  wire       [17:0]   fft_col_in_payload_4_imag;
  wire       [17:0]   fft_col_in_payload_5_real;
  wire       [17:0]   fft_col_in_payload_5_imag;
  wire       [17:0]   fft_col_in_payload_6_real;
  wire       [17:0]   fft_col_in_payload_6_imag;
  wire       [17:0]   fft_col_in_payload_7_real;
  wire       [17:0]   fft_col_in_payload_7_imag;
  wire       [17:0]   fft_col_in_payload_8_real;
  wire       [17:0]   fft_col_in_payload_8_imag;
  wire       [17:0]   fft_col_in_payload_9_real;
  wire       [17:0]   fft_col_in_payload_9_imag;
  wire       [17:0]   fft_col_in_payload_10_real;
  wire       [17:0]   fft_col_in_payload_10_imag;
  wire       [17:0]   fft_col_in_payload_11_real;
  wire       [17:0]   fft_col_in_payload_11_imag;
  wire       [17:0]   fft_col_in_payload_12_real;
  wire       [17:0]   fft_col_in_payload_12_imag;
  wire       [17:0]   fft_col_in_payload_13_real;
  wire       [17:0]   fft_col_in_payload_13_imag;
  wire       [17:0]   fft_col_in_payload_14_real;
  wire       [17:0]   fft_col_in_payload_14_imag;
  wire       [17:0]   fft_col_in_payload_15_real;
  wire       [17:0]   fft_col_in_payload_15_imag;
  wire       [17:0]   fft_col_in_payload_16_real;
  wire       [17:0]   fft_col_in_payload_16_imag;
  wire       [17:0]   fft_col_in_payload_17_real;
  wire       [17:0]   fft_col_in_payload_17_imag;
  wire       [17:0]   fft_col_in_payload_18_real;
  wire       [17:0]   fft_col_in_payload_18_imag;
  wire       [17:0]   fft_col_in_payload_19_real;
  wire       [17:0]   fft_col_in_payload_19_imag;
  wire       [17:0]   fft_col_in_payload_20_real;
  wire       [17:0]   fft_col_in_payload_20_imag;
  wire       [17:0]   fft_col_in_payload_21_real;
  wire       [17:0]   fft_col_in_payload_21_imag;
  wire       [17:0]   fft_col_in_payload_22_real;
  wire       [17:0]   fft_col_in_payload_22_imag;
  wire       [17:0]   fft_col_in_payload_23_real;
  wire       [17:0]   fft_col_in_payload_23_imag;
  wire       [17:0]   fft_col_in_payload_24_real;
  wire       [17:0]   fft_col_in_payload_24_imag;
  wire       [17:0]   fft_col_in_payload_25_real;
  wire       [17:0]   fft_col_in_payload_25_imag;
  wire       [17:0]   fft_col_in_payload_26_real;
  wire       [17:0]   fft_col_in_payload_26_imag;
  wire       [17:0]   fft_col_in_payload_27_real;
  wire       [17:0]   fft_col_in_payload_27_imag;
  wire       [17:0]   fft_col_in_payload_28_real;
  wire       [17:0]   fft_col_in_payload_28_imag;
  wire       [17:0]   fft_col_in_payload_29_real;
  wire       [17:0]   fft_col_in_payload_29_imag;
  wire       [17:0]   fft_col_in_payload_30_real;
  wire       [17:0]   fft_col_in_payload_30_imag;
  wire       [17:0]   fft_col_in_payload_31_real;
  wire       [17:0]   fft_col_in_payload_31_imag;
  wire       [17:0]   fft_col_in_payload_32_real;
  wire       [17:0]   fft_col_in_payload_32_imag;
  wire       [17:0]   fft_col_in_payload_33_real;
  wire       [17:0]   fft_col_in_payload_33_imag;
  wire       [17:0]   fft_col_in_payload_34_real;
  wire       [17:0]   fft_col_in_payload_34_imag;
  wire       [17:0]   fft_col_in_payload_35_real;
  wire       [17:0]   fft_col_in_payload_35_imag;
  wire       [17:0]   fft_col_in_payload_36_real;
  wire       [17:0]   fft_col_in_payload_36_imag;
  wire       [17:0]   fft_col_in_payload_37_real;
  wire       [17:0]   fft_col_in_payload_37_imag;
  wire       [17:0]   fft_col_in_payload_38_real;
  wire       [17:0]   fft_col_in_payload_38_imag;
  wire       [17:0]   fft_col_in_payload_39_real;
  wire       [17:0]   fft_col_in_payload_39_imag;
  wire       [17:0]   fft_col_in_payload_40_real;
  wire       [17:0]   fft_col_in_payload_40_imag;
  wire       [17:0]   fft_col_in_payload_41_real;
  wire       [17:0]   fft_col_in_payload_41_imag;
  wire       [17:0]   fft_col_in_payload_42_real;
  wire       [17:0]   fft_col_in_payload_42_imag;
  wire       [17:0]   fft_col_in_payload_43_real;
  wire       [17:0]   fft_col_in_payload_43_imag;
  wire       [17:0]   fft_col_in_payload_44_real;
  wire       [17:0]   fft_col_in_payload_44_imag;
  wire       [17:0]   fft_col_in_payload_45_real;
  wire       [17:0]   fft_col_in_payload_45_imag;
  wire       [17:0]   fft_col_in_payload_46_real;
  wire       [17:0]   fft_col_in_payload_46_imag;
  wire       [17:0]   fft_col_in_payload_47_real;
  wire       [17:0]   fft_col_in_payload_47_imag;
  wire       [17:0]   fft_col_in_payload_48_real;
  wire       [17:0]   fft_col_in_payload_48_imag;
  wire       [17:0]   fft_col_in_payload_49_real;
  wire       [17:0]   fft_col_in_payload_49_imag;
  wire       [17:0]   fft_col_in_payload_50_real;
  wire       [17:0]   fft_col_in_payload_50_imag;
  wire       [17:0]   fft_col_in_payload_51_real;
  wire       [17:0]   fft_col_in_payload_51_imag;
  wire       [17:0]   fft_col_in_payload_52_real;
  wire       [17:0]   fft_col_in_payload_52_imag;
  wire       [17:0]   fft_col_in_payload_53_real;
  wire       [17:0]   fft_col_in_payload_53_imag;
  wire       [17:0]   fft_col_in_payload_54_real;
  wire       [17:0]   fft_col_in_payload_54_imag;
  wire       [17:0]   fft_col_in_payload_55_real;
  wire       [17:0]   fft_col_in_payload_55_imag;
  wire       [17:0]   fft_col_in_payload_56_real;
  wire       [17:0]   fft_col_in_payload_56_imag;
  wire       [17:0]   fft_col_in_payload_57_real;
  wire       [17:0]   fft_col_in_payload_57_imag;
  wire       [17:0]   fft_col_in_payload_58_real;
  wire       [17:0]   fft_col_in_payload_58_imag;
  wire       [17:0]   fft_col_in_payload_59_real;
  wire       [17:0]   fft_col_in_payload_59_imag;
  wire       [17:0]   fft_col_in_payload_60_real;
  wire       [17:0]   fft_col_in_payload_60_imag;
  wire       [17:0]   fft_col_in_payload_61_real;
  wire       [17:0]   fft_col_in_payload_61_imag;
  wire       [17:0]   fft_col_in_payload_62_real;
  wire       [17:0]   fft_col_in_payload_62_imag;
  wire       [17:0]   fft_col_in_payload_63_real;
  wire       [17:0]   fft_col_in_payload_63_imag;
  reg                 null_cond_period_regNext;
  reg                 myFFT_3_fft_col_out_regNext_valid;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_0_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_0_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_1_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_1_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_2_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_2_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_3_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_3_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_4_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_4_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_5_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_5_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_6_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_6_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_7_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_7_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_8_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_8_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_9_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_9_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_10_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_10_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_11_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_11_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_12_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_12_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_13_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_13_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_14_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_14_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_15_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_15_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_16_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_16_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_17_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_17_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_18_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_18_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_19_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_19_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_20_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_20_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_21_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_21_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_22_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_22_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_23_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_23_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_24_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_24_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_25_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_25_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_26_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_26_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_27_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_27_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_28_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_28_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_29_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_29_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_30_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_30_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_31_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_31_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_32_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_32_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_33_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_33_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_34_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_34_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_35_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_35_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_36_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_36_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_37_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_37_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_38_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_38_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_39_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_39_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_40_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_40_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_41_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_41_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_42_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_42_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_43_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_43_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_44_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_44_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_45_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_45_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_46_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_46_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_47_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_47_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_48_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_48_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_49_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_49_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_50_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_50_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_51_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_51_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_52_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_52_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_53_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_53_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_54_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_54_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_55_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_55_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_56_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_56_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_57_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_57_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_58_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_58_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_59_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_59_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_60_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_60_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_61_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_61_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_62_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_62_imag;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_63_real;
  reg        [17:0]   myFFT_3_fft_col_out_regNext_payload_63_imag;

  assign _zz_322 = row_addr_willIncrement;
  assign _zz_323 = {5'd0, _zz_322};
  assign _zz_324 = null_cnt_willIncrement;
  assign _zz_325 = {5'd0, _zz_324};
  MyFFT myFFT_2 (
    .io_data_in_valid              (io_line_in_valid                       ), //i
    .io_data_in_payload_0_real     (io_line_in_payload_0_real[17:0]        ), //i
    .io_data_in_payload_0_imag     (io_line_in_payload_0_imag[17:0]        ), //i
    .io_data_in_payload_1_real     (io_line_in_payload_1_real[17:0]        ), //i
    .io_data_in_payload_1_imag     (io_line_in_payload_1_imag[17:0]        ), //i
    .io_data_in_payload_2_real     (io_line_in_payload_2_real[17:0]        ), //i
    .io_data_in_payload_2_imag     (io_line_in_payload_2_imag[17:0]        ), //i
    .io_data_in_payload_3_real     (io_line_in_payload_3_real[17:0]        ), //i
    .io_data_in_payload_3_imag     (io_line_in_payload_3_imag[17:0]        ), //i
    .io_data_in_payload_4_real     (io_line_in_payload_4_real[17:0]        ), //i
    .io_data_in_payload_4_imag     (io_line_in_payload_4_imag[17:0]        ), //i
    .io_data_in_payload_5_real     (io_line_in_payload_5_real[17:0]        ), //i
    .io_data_in_payload_5_imag     (io_line_in_payload_5_imag[17:0]        ), //i
    .io_data_in_payload_6_real     (io_line_in_payload_6_real[17:0]        ), //i
    .io_data_in_payload_6_imag     (io_line_in_payload_6_imag[17:0]        ), //i
    .io_data_in_payload_7_real     (io_line_in_payload_7_real[17:0]        ), //i
    .io_data_in_payload_7_imag     (io_line_in_payload_7_imag[17:0]        ), //i
    .io_data_in_payload_8_real     (io_line_in_payload_8_real[17:0]        ), //i
    .io_data_in_payload_8_imag     (io_line_in_payload_8_imag[17:0]        ), //i
    .io_data_in_payload_9_real     (io_line_in_payload_9_real[17:0]        ), //i
    .io_data_in_payload_9_imag     (io_line_in_payload_9_imag[17:0]        ), //i
    .io_data_in_payload_10_real    (io_line_in_payload_10_real[17:0]       ), //i
    .io_data_in_payload_10_imag    (io_line_in_payload_10_imag[17:0]       ), //i
    .io_data_in_payload_11_real    (io_line_in_payload_11_real[17:0]       ), //i
    .io_data_in_payload_11_imag    (io_line_in_payload_11_imag[17:0]       ), //i
    .io_data_in_payload_12_real    (io_line_in_payload_12_real[17:0]       ), //i
    .io_data_in_payload_12_imag    (io_line_in_payload_12_imag[17:0]       ), //i
    .io_data_in_payload_13_real    (io_line_in_payload_13_real[17:0]       ), //i
    .io_data_in_payload_13_imag    (io_line_in_payload_13_imag[17:0]       ), //i
    .io_data_in_payload_14_real    (io_line_in_payload_14_real[17:0]       ), //i
    .io_data_in_payload_14_imag    (io_line_in_payload_14_imag[17:0]       ), //i
    .io_data_in_payload_15_real    (io_line_in_payload_15_real[17:0]       ), //i
    .io_data_in_payload_15_imag    (io_line_in_payload_15_imag[17:0]       ), //i
    .io_data_in_payload_16_real    (io_line_in_payload_16_real[17:0]       ), //i
    .io_data_in_payload_16_imag    (io_line_in_payload_16_imag[17:0]       ), //i
    .io_data_in_payload_17_real    (io_line_in_payload_17_real[17:0]       ), //i
    .io_data_in_payload_17_imag    (io_line_in_payload_17_imag[17:0]       ), //i
    .io_data_in_payload_18_real    (io_line_in_payload_18_real[17:0]       ), //i
    .io_data_in_payload_18_imag    (io_line_in_payload_18_imag[17:0]       ), //i
    .io_data_in_payload_19_real    (io_line_in_payload_19_real[17:0]       ), //i
    .io_data_in_payload_19_imag    (io_line_in_payload_19_imag[17:0]       ), //i
    .io_data_in_payload_20_real    (io_line_in_payload_20_real[17:0]       ), //i
    .io_data_in_payload_20_imag    (io_line_in_payload_20_imag[17:0]       ), //i
    .io_data_in_payload_21_real    (io_line_in_payload_21_real[17:0]       ), //i
    .io_data_in_payload_21_imag    (io_line_in_payload_21_imag[17:0]       ), //i
    .io_data_in_payload_22_real    (io_line_in_payload_22_real[17:0]       ), //i
    .io_data_in_payload_22_imag    (io_line_in_payload_22_imag[17:0]       ), //i
    .io_data_in_payload_23_real    (io_line_in_payload_23_real[17:0]       ), //i
    .io_data_in_payload_23_imag    (io_line_in_payload_23_imag[17:0]       ), //i
    .io_data_in_payload_24_real    (io_line_in_payload_24_real[17:0]       ), //i
    .io_data_in_payload_24_imag    (io_line_in_payload_24_imag[17:0]       ), //i
    .io_data_in_payload_25_real    (io_line_in_payload_25_real[17:0]       ), //i
    .io_data_in_payload_25_imag    (io_line_in_payload_25_imag[17:0]       ), //i
    .io_data_in_payload_26_real    (io_line_in_payload_26_real[17:0]       ), //i
    .io_data_in_payload_26_imag    (io_line_in_payload_26_imag[17:0]       ), //i
    .io_data_in_payload_27_real    (io_line_in_payload_27_real[17:0]       ), //i
    .io_data_in_payload_27_imag    (io_line_in_payload_27_imag[17:0]       ), //i
    .io_data_in_payload_28_real    (io_line_in_payload_28_real[17:0]       ), //i
    .io_data_in_payload_28_imag    (io_line_in_payload_28_imag[17:0]       ), //i
    .io_data_in_payload_29_real    (io_line_in_payload_29_real[17:0]       ), //i
    .io_data_in_payload_29_imag    (io_line_in_payload_29_imag[17:0]       ), //i
    .io_data_in_payload_30_real    (io_line_in_payload_30_real[17:0]       ), //i
    .io_data_in_payload_30_imag    (io_line_in_payload_30_imag[17:0]       ), //i
    .io_data_in_payload_31_real    (io_line_in_payload_31_real[17:0]       ), //i
    .io_data_in_payload_31_imag    (io_line_in_payload_31_imag[17:0]       ), //i
    .io_data_in_payload_32_real    (io_line_in_payload_32_real[17:0]       ), //i
    .io_data_in_payload_32_imag    (io_line_in_payload_32_imag[17:0]       ), //i
    .io_data_in_payload_33_real    (io_line_in_payload_33_real[17:0]       ), //i
    .io_data_in_payload_33_imag    (io_line_in_payload_33_imag[17:0]       ), //i
    .io_data_in_payload_34_real    (io_line_in_payload_34_real[17:0]       ), //i
    .io_data_in_payload_34_imag    (io_line_in_payload_34_imag[17:0]       ), //i
    .io_data_in_payload_35_real    (io_line_in_payload_35_real[17:0]       ), //i
    .io_data_in_payload_35_imag    (io_line_in_payload_35_imag[17:0]       ), //i
    .io_data_in_payload_36_real    (io_line_in_payload_36_real[17:0]       ), //i
    .io_data_in_payload_36_imag    (io_line_in_payload_36_imag[17:0]       ), //i
    .io_data_in_payload_37_real    (io_line_in_payload_37_real[17:0]       ), //i
    .io_data_in_payload_37_imag    (io_line_in_payload_37_imag[17:0]       ), //i
    .io_data_in_payload_38_real    (io_line_in_payload_38_real[17:0]       ), //i
    .io_data_in_payload_38_imag    (io_line_in_payload_38_imag[17:0]       ), //i
    .io_data_in_payload_39_real    (io_line_in_payload_39_real[17:0]       ), //i
    .io_data_in_payload_39_imag    (io_line_in_payload_39_imag[17:0]       ), //i
    .io_data_in_payload_40_real    (io_line_in_payload_40_real[17:0]       ), //i
    .io_data_in_payload_40_imag    (io_line_in_payload_40_imag[17:0]       ), //i
    .io_data_in_payload_41_real    (io_line_in_payload_41_real[17:0]       ), //i
    .io_data_in_payload_41_imag    (io_line_in_payload_41_imag[17:0]       ), //i
    .io_data_in_payload_42_real    (io_line_in_payload_42_real[17:0]       ), //i
    .io_data_in_payload_42_imag    (io_line_in_payload_42_imag[17:0]       ), //i
    .io_data_in_payload_43_real    (io_line_in_payload_43_real[17:0]       ), //i
    .io_data_in_payload_43_imag    (io_line_in_payload_43_imag[17:0]       ), //i
    .io_data_in_payload_44_real    (io_line_in_payload_44_real[17:0]       ), //i
    .io_data_in_payload_44_imag    (io_line_in_payload_44_imag[17:0]       ), //i
    .io_data_in_payload_45_real    (io_line_in_payload_45_real[17:0]       ), //i
    .io_data_in_payload_45_imag    (io_line_in_payload_45_imag[17:0]       ), //i
    .io_data_in_payload_46_real    (io_line_in_payload_46_real[17:0]       ), //i
    .io_data_in_payload_46_imag    (io_line_in_payload_46_imag[17:0]       ), //i
    .io_data_in_payload_47_real    (io_line_in_payload_47_real[17:0]       ), //i
    .io_data_in_payload_47_imag    (io_line_in_payload_47_imag[17:0]       ), //i
    .io_data_in_payload_48_real    (io_line_in_payload_48_real[17:0]       ), //i
    .io_data_in_payload_48_imag    (io_line_in_payload_48_imag[17:0]       ), //i
    .io_data_in_payload_49_real    (io_line_in_payload_49_real[17:0]       ), //i
    .io_data_in_payload_49_imag    (io_line_in_payload_49_imag[17:0]       ), //i
    .io_data_in_payload_50_real    (io_line_in_payload_50_real[17:0]       ), //i
    .io_data_in_payload_50_imag    (io_line_in_payload_50_imag[17:0]       ), //i
    .io_data_in_payload_51_real    (io_line_in_payload_51_real[17:0]       ), //i
    .io_data_in_payload_51_imag    (io_line_in_payload_51_imag[17:0]       ), //i
    .io_data_in_payload_52_real    (io_line_in_payload_52_real[17:0]       ), //i
    .io_data_in_payload_52_imag    (io_line_in_payload_52_imag[17:0]       ), //i
    .io_data_in_payload_53_real    (io_line_in_payload_53_real[17:0]       ), //i
    .io_data_in_payload_53_imag    (io_line_in_payload_53_imag[17:0]       ), //i
    .io_data_in_payload_54_real    (io_line_in_payload_54_real[17:0]       ), //i
    .io_data_in_payload_54_imag    (io_line_in_payload_54_imag[17:0]       ), //i
    .io_data_in_payload_55_real    (io_line_in_payload_55_real[17:0]       ), //i
    .io_data_in_payload_55_imag    (io_line_in_payload_55_imag[17:0]       ), //i
    .io_data_in_payload_56_real    (io_line_in_payload_56_real[17:0]       ), //i
    .io_data_in_payload_56_imag    (io_line_in_payload_56_imag[17:0]       ), //i
    .io_data_in_payload_57_real    (io_line_in_payload_57_real[17:0]       ), //i
    .io_data_in_payload_57_imag    (io_line_in_payload_57_imag[17:0]       ), //i
    .io_data_in_payload_58_real    (io_line_in_payload_58_real[17:0]       ), //i
    .io_data_in_payload_58_imag    (io_line_in_payload_58_imag[17:0]       ), //i
    .io_data_in_payload_59_real    (io_line_in_payload_59_real[17:0]       ), //i
    .io_data_in_payload_59_imag    (io_line_in_payload_59_imag[17:0]       ), //i
    .io_data_in_payload_60_real    (io_line_in_payload_60_real[17:0]       ), //i
    .io_data_in_payload_60_imag    (io_line_in_payload_60_imag[17:0]       ), //i
    .io_data_in_payload_61_real    (io_line_in_payload_61_real[17:0]       ), //i
    .io_data_in_payload_61_imag    (io_line_in_payload_61_imag[17:0]       ), //i
    .io_data_in_payload_62_real    (io_line_in_payload_62_real[17:0]       ), //i
    .io_data_in_payload_62_imag    (io_line_in_payload_62_imag[17:0]       ), //i
    .io_data_in_payload_63_real    (io_line_in_payload_63_real[17:0]       ), //i
    .io_data_in_payload_63_imag    (io_line_in_payload_63_imag[17:0]       ), //i
    .fft_row_valid                 (myFFT_2_fft_row_valid                  ), //o
    .fft_row_payload_0_real        (myFFT_2_fft_row_payload_0_real[17:0]   ), //o
    .fft_row_payload_0_imag        (myFFT_2_fft_row_payload_0_imag[17:0]   ), //o
    .fft_row_payload_1_real        (myFFT_2_fft_row_payload_1_real[17:0]   ), //o
    .fft_row_payload_1_imag        (myFFT_2_fft_row_payload_1_imag[17:0]   ), //o
    .fft_row_payload_2_real        (myFFT_2_fft_row_payload_2_real[17:0]   ), //o
    .fft_row_payload_2_imag        (myFFT_2_fft_row_payload_2_imag[17:0]   ), //o
    .fft_row_payload_3_real        (myFFT_2_fft_row_payload_3_real[17:0]   ), //o
    .fft_row_payload_3_imag        (myFFT_2_fft_row_payload_3_imag[17:0]   ), //o
    .fft_row_payload_4_real        (myFFT_2_fft_row_payload_4_real[17:0]   ), //o
    .fft_row_payload_4_imag        (myFFT_2_fft_row_payload_4_imag[17:0]   ), //o
    .fft_row_payload_5_real        (myFFT_2_fft_row_payload_5_real[17:0]   ), //o
    .fft_row_payload_5_imag        (myFFT_2_fft_row_payload_5_imag[17:0]   ), //o
    .fft_row_payload_6_real        (myFFT_2_fft_row_payload_6_real[17:0]   ), //o
    .fft_row_payload_6_imag        (myFFT_2_fft_row_payload_6_imag[17:0]   ), //o
    .fft_row_payload_7_real        (myFFT_2_fft_row_payload_7_real[17:0]   ), //o
    .fft_row_payload_7_imag        (myFFT_2_fft_row_payload_7_imag[17:0]   ), //o
    .fft_row_payload_8_real        (myFFT_2_fft_row_payload_8_real[17:0]   ), //o
    .fft_row_payload_8_imag        (myFFT_2_fft_row_payload_8_imag[17:0]   ), //o
    .fft_row_payload_9_real        (myFFT_2_fft_row_payload_9_real[17:0]   ), //o
    .fft_row_payload_9_imag        (myFFT_2_fft_row_payload_9_imag[17:0]   ), //o
    .fft_row_payload_10_real       (myFFT_2_fft_row_payload_10_real[17:0]  ), //o
    .fft_row_payload_10_imag       (myFFT_2_fft_row_payload_10_imag[17:0]  ), //o
    .fft_row_payload_11_real       (myFFT_2_fft_row_payload_11_real[17:0]  ), //o
    .fft_row_payload_11_imag       (myFFT_2_fft_row_payload_11_imag[17:0]  ), //o
    .fft_row_payload_12_real       (myFFT_2_fft_row_payload_12_real[17:0]  ), //o
    .fft_row_payload_12_imag       (myFFT_2_fft_row_payload_12_imag[17:0]  ), //o
    .fft_row_payload_13_real       (myFFT_2_fft_row_payload_13_real[17:0]  ), //o
    .fft_row_payload_13_imag       (myFFT_2_fft_row_payload_13_imag[17:0]  ), //o
    .fft_row_payload_14_real       (myFFT_2_fft_row_payload_14_real[17:0]  ), //o
    .fft_row_payload_14_imag       (myFFT_2_fft_row_payload_14_imag[17:0]  ), //o
    .fft_row_payload_15_real       (myFFT_2_fft_row_payload_15_real[17:0]  ), //o
    .fft_row_payload_15_imag       (myFFT_2_fft_row_payload_15_imag[17:0]  ), //o
    .fft_row_payload_16_real       (myFFT_2_fft_row_payload_16_real[17:0]  ), //o
    .fft_row_payload_16_imag       (myFFT_2_fft_row_payload_16_imag[17:0]  ), //o
    .fft_row_payload_17_real       (myFFT_2_fft_row_payload_17_real[17:0]  ), //o
    .fft_row_payload_17_imag       (myFFT_2_fft_row_payload_17_imag[17:0]  ), //o
    .fft_row_payload_18_real       (myFFT_2_fft_row_payload_18_real[17:0]  ), //o
    .fft_row_payload_18_imag       (myFFT_2_fft_row_payload_18_imag[17:0]  ), //o
    .fft_row_payload_19_real       (myFFT_2_fft_row_payload_19_real[17:0]  ), //o
    .fft_row_payload_19_imag       (myFFT_2_fft_row_payload_19_imag[17:0]  ), //o
    .fft_row_payload_20_real       (myFFT_2_fft_row_payload_20_real[17:0]  ), //o
    .fft_row_payload_20_imag       (myFFT_2_fft_row_payload_20_imag[17:0]  ), //o
    .fft_row_payload_21_real       (myFFT_2_fft_row_payload_21_real[17:0]  ), //o
    .fft_row_payload_21_imag       (myFFT_2_fft_row_payload_21_imag[17:0]  ), //o
    .fft_row_payload_22_real       (myFFT_2_fft_row_payload_22_real[17:0]  ), //o
    .fft_row_payload_22_imag       (myFFT_2_fft_row_payload_22_imag[17:0]  ), //o
    .fft_row_payload_23_real       (myFFT_2_fft_row_payload_23_real[17:0]  ), //o
    .fft_row_payload_23_imag       (myFFT_2_fft_row_payload_23_imag[17:0]  ), //o
    .fft_row_payload_24_real       (myFFT_2_fft_row_payload_24_real[17:0]  ), //o
    .fft_row_payload_24_imag       (myFFT_2_fft_row_payload_24_imag[17:0]  ), //o
    .fft_row_payload_25_real       (myFFT_2_fft_row_payload_25_real[17:0]  ), //o
    .fft_row_payload_25_imag       (myFFT_2_fft_row_payload_25_imag[17:0]  ), //o
    .fft_row_payload_26_real       (myFFT_2_fft_row_payload_26_real[17:0]  ), //o
    .fft_row_payload_26_imag       (myFFT_2_fft_row_payload_26_imag[17:0]  ), //o
    .fft_row_payload_27_real       (myFFT_2_fft_row_payload_27_real[17:0]  ), //o
    .fft_row_payload_27_imag       (myFFT_2_fft_row_payload_27_imag[17:0]  ), //o
    .fft_row_payload_28_real       (myFFT_2_fft_row_payload_28_real[17:0]  ), //o
    .fft_row_payload_28_imag       (myFFT_2_fft_row_payload_28_imag[17:0]  ), //o
    .fft_row_payload_29_real       (myFFT_2_fft_row_payload_29_real[17:0]  ), //o
    .fft_row_payload_29_imag       (myFFT_2_fft_row_payload_29_imag[17:0]  ), //o
    .fft_row_payload_30_real       (myFFT_2_fft_row_payload_30_real[17:0]  ), //o
    .fft_row_payload_30_imag       (myFFT_2_fft_row_payload_30_imag[17:0]  ), //o
    .fft_row_payload_31_real       (myFFT_2_fft_row_payload_31_real[17:0]  ), //o
    .fft_row_payload_31_imag       (myFFT_2_fft_row_payload_31_imag[17:0]  ), //o
    .fft_row_payload_32_real       (myFFT_2_fft_row_payload_32_real[17:0]  ), //o
    .fft_row_payload_32_imag       (myFFT_2_fft_row_payload_32_imag[17:0]  ), //o
    .fft_row_payload_33_real       (myFFT_2_fft_row_payload_33_real[17:0]  ), //o
    .fft_row_payload_33_imag       (myFFT_2_fft_row_payload_33_imag[17:0]  ), //o
    .fft_row_payload_34_real       (myFFT_2_fft_row_payload_34_real[17:0]  ), //o
    .fft_row_payload_34_imag       (myFFT_2_fft_row_payload_34_imag[17:0]  ), //o
    .fft_row_payload_35_real       (myFFT_2_fft_row_payload_35_real[17:0]  ), //o
    .fft_row_payload_35_imag       (myFFT_2_fft_row_payload_35_imag[17:0]  ), //o
    .fft_row_payload_36_real       (myFFT_2_fft_row_payload_36_real[17:0]  ), //o
    .fft_row_payload_36_imag       (myFFT_2_fft_row_payload_36_imag[17:0]  ), //o
    .fft_row_payload_37_real       (myFFT_2_fft_row_payload_37_real[17:0]  ), //o
    .fft_row_payload_37_imag       (myFFT_2_fft_row_payload_37_imag[17:0]  ), //o
    .fft_row_payload_38_real       (myFFT_2_fft_row_payload_38_real[17:0]  ), //o
    .fft_row_payload_38_imag       (myFFT_2_fft_row_payload_38_imag[17:0]  ), //o
    .fft_row_payload_39_real       (myFFT_2_fft_row_payload_39_real[17:0]  ), //o
    .fft_row_payload_39_imag       (myFFT_2_fft_row_payload_39_imag[17:0]  ), //o
    .fft_row_payload_40_real       (myFFT_2_fft_row_payload_40_real[17:0]  ), //o
    .fft_row_payload_40_imag       (myFFT_2_fft_row_payload_40_imag[17:0]  ), //o
    .fft_row_payload_41_real       (myFFT_2_fft_row_payload_41_real[17:0]  ), //o
    .fft_row_payload_41_imag       (myFFT_2_fft_row_payload_41_imag[17:0]  ), //o
    .fft_row_payload_42_real       (myFFT_2_fft_row_payload_42_real[17:0]  ), //o
    .fft_row_payload_42_imag       (myFFT_2_fft_row_payload_42_imag[17:0]  ), //o
    .fft_row_payload_43_real       (myFFT_2_fft_row_payload_43_real[17:0]  ), //o
    .fft_row_payload_43_imag       (myFFT_2_fft_row_payload_43_imag[17:0]  ), //o
    .fft_row_payload_44_real       (myFFT_2_fft_row_payload_44_real[17:0]  ), //o
    .fft_row_payload_44_imag       (myFFT_2_fft_row_payload_44_imag[17:0]  ), //o
    .fft_row_payload_45_real       (myFFT_2_fft_row_payload_45_real[17:0]  ), //o
    .fft_row_payload_45_imag       (myFFT_2_fft_row_payload_45_imag[17:0]  ), //o
    .fft_row_payload_46_real       (myFFT_2_fft_row_payload_46_real[17:0]  ), //o
    .fft_row_payload_46_imag       (myFFT_2_fft_row_payload_46_imag[17:0]  ), //o
    .fft_row_payload_47_real       (myFFT_2_fft_row_payload_47_real[17:0]  ), //o
    .fft_row_payload_47_imag       (myFFT_2_fft_row_payload_47_imag[17:0]  ), //o
    .fft_row_payload_48_real       (myFFT_2_fft_row_payload_48_real[17:0]  ), //o
    .fft_row_payload_48_imag       (myFFT_2_fft_row_payload_48_imag[17:0]  ), //o
    .fft_row_payload_49_real       (myFFT_2_fft_row_payload_49_real[17:0]  ), //o
    .fft_row_payload_49_imag       (myFFT_2_fft_row_payload_49_imag[17:0]  ), //o
    .fft_row_payload_50_real       (myFFT_2_fft_row_payload_50_real[17:0]  ), //o
    .fft_row_payload_50_imag       (myFFT_2_fft_row_payload_50_imag[17:0]  ), //o
    .fft_row_payload_51_real       (myFFT_2_fft_row_payload_51_real[17:0]  ), //o
    .fft_row_payload_51_imag       (myFFT_2_fft_row_payload_51_imag[17:0]  ), //o
    .fft_row_payload_52_real       (myFFT_2_fft_row_payload_52_real[17:0]  ), //o
    .fft_row_payload_52_imag       (myFFT_2_fft_row_payload_52_imag[17:0]  ), //o
    .fft_row_payload_53_real       (myFFT_2_fft_row_payload_53_real[17:0]  ), //o
    .fft_row_payload_53_imag       (myFFT_2_fft_row_payload_53_imag[17:0]  ), //o
    .fft_row_payload_54_real       (myFFT_2_fft_row_payload_54_real[17:0]  ), //o
    .fft_row_payload_54_imag       (myFFT_2_fft_row_payload_54_imag[17:0]  ), //o
    .fft_row_payload_55_real       (myFFT_2_fft_row_payload_55_real[17:0]  ), //o
    .fft_row_payload_55_imag       (myFFT_2_fft_row_payload_55_imag[17:0]  ), //o
    .fft_row_payload_56_real       (myFFT_2_fft_row_payload_56_real[17:0]  ), //o
    .fft_row_payload_56_imag       (myFFT_2_fft_row_payload_56_imag[17:0]  ), //o
    .fft_row_payload_57_real       (myFFT_2_fft_row_payload_57_real[17:0]  ), //o
    .fft_row_payload_57_imag       (myFFT_2_fft_row_payload_57_imag[17:0]  ), //o
    .fft_row_payload_58_real       (myFFT_2_fft_row_payload_58_real[17:0]  ), //o
    .fft_row_payload_58_imag       (myFFT_2_fft_row_payload_58_imag[17:0]  ), //o
    .fft_row_payload_59_real       (myFFT_2_fft_row_payload_59_real[17:0]  ), //o
    .fft_row_payload_59_imag       (myFFT_2_fft_row_payload_59_imag[17:0]  ), //o
    .fft_row_payload_60_real       (myFFT_2_fft_row_payload_60_real[17:0]  ), //o
    .fft_row_payload_60_imag       (myFFT_2_fft_row_payload_60_imag[17:0]  ), //o
    .fft_row_payload_61_real       (myFFT_2_fft_row_payload_61_real[17:0]  ), //o
    .fft_row_payload_61_imag       (myFFT_2_fft_row_payload_61_imag[17:0]  ), //o
    .fft_row_payload_62_real       (myFFT_2_fft_row_payload_62_real[17:0]  ), //o
    .fft_row_payload_62_imag       (myFFT_2_fft_row_payload_62_imag[17:0]  ), //o
    .fft_row_payload_63_real       (myFFT_2_fft_row_payload_63_real[17:0]  ), //o
    .fft_row_payload_63_imag       (myFFT_2_fft_row_payload_63_imag[17:0]  ), //o
    .clk                           (clk                                    ), //i
    .reset                         (reset                                  )  //i
  );
  MyFFT_1 myFFT_3 (
    .io_data_in_valid               (fft_col_in_valid                           ), //i
    .io_data_in_payload_0_real      (fft_col_in_payload_0_real[17:0]            ), //i
    .io_data_in_payload_0_imag      (fft_col_in_payload_0_imag[17:0]            ), //i
    .io_data_in_payload_1_real      (fft_col_in_payload_1_real[17:0]            ), //i
    .io_data_in_payload_1_imag      (fft_col_in_payload_1_imag[17:0]            ), //i
    .io_data_in_payload_2_real      (fft_col_in_payload_2_real[17:0]            ), //i
    .io_data_in_payload_2_imag      (fft_col_in_payload_2_imag[17:0]            ), //i
    .io_data_in_payload_3_real      (fft_col_in_payload_3_real[17:0]            ), //i
    .io_data_in_payload_3_imag      (fft_col_in_payload_3_imag[17:0]            ), //i
    .io_data_in_payload_4_real      (fft_col_in_payload_4_real[17:0]            ), //i
    .io_data_in_payload_4_imag      (fft_col_in_payload_4_imag[17:0]            ), //i
    .io_data_in_payload_5_real      (fft_col_in_payload_5_real[17:0]            ), //i
    .io_data_in_payload_5_imag      (fft_col_in_payload_5_imag[17:0]            ), //i
    .io_data_in_payload_6_real      (fft_col_in_payload_6_real[17:0]            ), //i
    .io_data_in_payload_6_imag      (fft_col_in_payload_6_imag[17:0]            ), //i
    .io_data_in_payload_7_real      (fft_col_in_payload_7_real[17:0]            ), //i
    .io_data_in_payload_7_imag      (fft_col_in_payload_7_imag[17:0]            ), //i
    .io_data_in_payload_8_real      (fft_col_in_payload_8_real[17:0]            ), //i
    .io_data_in_payload_8_imag      (fft_col_in_payload_8_imag[17:0]            ), //i
    .io_data_in_payload_9_real      (fft_col_in_payload_9_real[17:0]            ), //i
    .io_data_in_payload_9_imag      (fft_col_in_payload_9_imag[17:0]            ), //i
    .io_data_in_payload_10_real     (fft_col_in_payload_10_real[17:0]           ), //i
    .io_data_in_payload_10_imag     (fft_col_in_payload_10_imag[17:0]           ), //i
    .io_data_in_payload_11_real     (fft_col_in_payload_11_real[17:0]           ), //i
    .io_data_in_payload_11_imag     (fft_col_in_payload_11_imag[17:0]           ), //i
    .io_data_in_payload_12_real     (fft_col_in_payload_12_real[17:0]           ), //i
    .io_data_in_payload_12_imag     (fft_col_in_payload_12_imag[17:0]           ), //i
    .io_data_in_payload_13_real     (fft_col_in_payload_13_real[17:0]           ), //i
    .io_data_in_payload_13_imag     (fft_col_in_payload_13_imag[17:0]           ), //i
    .io_data_in_payload_14_real     (fft_col_in_payload_14_real[17:0]           ), //i
    .io_data_in_payload_14_imag     (fft_col_in_payload_14_imag[17:0]           ), //i
    .io_data_in_payload_15_real     (fft_col_in_payload_15_real[17:0]           ), //i
    .io_data_in_payload_15_imag     (fft_col_in_payload_15_imag[17:0]           ), //i
    .io_data_in_payload_16_real     (fft_col_in_payload_16_real[17:0]           ), //i
    .io_data_in_payload_16_imag     (fft_col_in_payload_16_imag[17:0]           ), //i
    .io_data_in_payload_17_real     (fft_col_in_payload_17_real[17:0]           ), //i
    .io_data_in_payload_17_imag     (fft_col_in_payload_17_imag[17:0]           ), //i
    .io_data_in_payload_18_real     (fft_col_in_payload_18_real[17:0]           ), //i
    .io_data_in_payload_18_imag     (fft_col_in_payload_18_imag[17:0]           ), //i
    .io_data_in_payload_19_real     (fft_col_in_payload_19_real[17:0]           ), //i
    .io_data_in_payload_19_imag     (fft_col_in_payload_19_imag[17:0]           ), //i
    .io_data_in_payload_20_real     (fft_col_in_payload_20_real[17:0]           ), //i
    .io_data_in_payload_20_imag     (fft_col_in_payload_20_imag[17:0]           ), //i
    .io_data_in_payload_21_real     (fft_col_in_payload_21_real[17:0]           ), //i
    .io_data_in_payload_21_imag     (fft_col_in_payload_21_imag[17:0]           ), //i
    .io_data_in_payload_22_real     (fft_col_in_payload_22_real[17:0]           ), //i
    .io_data_in_payload_22_imag     (fft_col_in_payload_22_imag[17:0]           ), //i
    .io_data_in_payload_23_real     (fft_col_in_payload_23_real[17:0]           ), //i
    .io_data_in_payload_23_imag     (fft_col_in_payload_23_imag[17:0]           ), //i
    .io_data_in_payload_24_real     (fft_col_in_payload_24_real[17:0]           ), //i
    .io_data_in_payload_24_imag     (fft_col_in_payload_24_imag[17:0]           ), //i
    .io_data_in_payload_25_real     (fft_col_in_payload_25_real[17:0]           ), //i
    .io_data_in_payload_25_imag     (fft_col_in_payload_25_imag[17:0]           ), //i
    .io_data_in_payload_26_real     (fft_col_in_payload_26_real[17:0]           ), //i
    .io_data_in_payload_26_imag     (fft_col_in_payload_26_imag[17:0]           ), //i
    .io_data_in_payload_27_real     (fft_col_in_payload_27_real[17:0]           ), //i
    .io_data_in_payload_27_imag     (fft_col_in_payload_27_imag[17:0]           ), //i
    .io_data_in_payload_28_real     (fft_col_in_payload_28_real[17:0]           ), //i
    .io_data_in_payload_28_imag     (fft_col_in_payload_28_imag[17:0]           ), //i
    .io_data_in_payload_29_real     (fft_col_in_payload_29_real[17:0]           ), //i
    .io_data_in_payload_29_imag     (fft_col_in_payload_29_imag[17:0]           ), //i
    .io_data_in_payload_30_real     (fft_col_in_payload_30_real[17:0]           ), //i
    .io_data_in_payload_30_imag     (fft_col_in_payload_30_imag[17:0]           ), //i
    .io_data_in_payload_31_real     (fft_col_in_payload_31_real[17:0]           ), //i
    .io_data_in_payload_31_imag     (fft_col_in_payload_31_imag[17:0]           ), //i
    .io_data_in_payload_32_real     (fft_col_in_payload_32_real[17:0]           ), //i
    .io_data_in_payload_32_imag     (fft_col_in_payload_32_imag[17:0]           ), //i
    .io_data_in_payload_33_real     (fft_col_in_payload_33_real[17:0]           ), //i
    .io_data_in_payload_33_imag     (fft_col_in_payload_33_imag[17:0]           ), //i
    .io_data_in_payload_34_real     (fft_col_in_payload_34_real[17:0]           ), //i
    .io_data_in_payload_34_imag     (fft_col_in_payload_34_imag[17:0]           ), //i
    .io_data_in_payload_35_real     (fft_col_in_payload_35_real[17:0]           ), //i
    .io_data_in_payload_35_imag     (fft_col_in_payload_35_imag[17:0]           ), //i
    .io_data_in_payload_36_real     (fft_col_in_payload_36_real[17:0]           ), //i
    .io_data_in_payload_36_imag     (fft_col_in_payload_36_imag[17:0]           ), //i
    .io_data_in_payload_37_real     (fft_col_in_payload_37_real[17:0]           ), //i
    .io_data_in_payload_37_imag     (fft_col_in_payload_37_imag[17:0]           ), //i
    .io_data_in_payload_38_real     (fft_col_in_payload_38_real[17:0]           ), //i
    .io_data_in_payload_38_imag     (fft_col_in_payload_38_imag[17:0]           ), //i
    .io_data_in_payload_39_real     (fft_col_in_payload_39_real[17:0]           ), //i
    .io_data_in_payload_39_imag     (fft_col_in_payload_39_imag[17:0]           ), //i
    .io_data_in_payload_40_real     (fft_col_in_payload_40_real[17:0]           ), //i
    .io_data_in_payload_40_imag     (fft_col_in_payload_40_imag[17:0]           ), //i
    .io_data_in_payload_41_real     (fft_col_in_payload_41_real[17:0]           ), //i
    .io_data_in_payload_41_imag     (fft_col_in_payload_41_imag[17:0]           ), //i
    .io_data_in_payload_42_real     (fft_col_in_payload_42_real[17:0]           ), //i
    .io_data_in_payload_42_imag     (fft_col_in_payload_42_imag[17:0]           ), //i
    .io_data_in_payload_43_real     (fft_col_in_payload_43_real[17:0]           ), //i
    .io_data_in_payload_43_imag     (fft_col_in_payload_43_imag[17:0]           ), //i
    .io_data_in_payload_44_real     (fft_col_in_payload_44_real[17:0]           ), //i
    .io_data_in_payload_44_imag     (fft_col_in_payload_44_imag[17:0]           ), //i
    .io_data_in_payload_45_real     (fft_col_in_payload_45_real[17:0]           ), //i
    .io_data_in_payload_45_imag     (fft_col_in_payload_45_imag[17:0]           ), //i
    .io_data_in_payload_46_real     (fft_col_in_payload_46_real[17:0]           ), //i
    .io_data_in_payload_46_imag     (fft_col_in_payload_46_imag[17:0]           ), //i
    .io_data_in_payload_47_real     (fft_col_in_payload_47_real[17:0]           ), //i
    .io_data_in_payload_47_imag     (fft_col_in_payload_47_imag[17:0]           ), //i
    .io_data_in_payload_48_real     (fft_col_in_payload_48_real[17:0]           ), //i
    .io_data_in_payload_48_imag     (fft_col_in_payload_48_imag[17:0]           ), //i
    .io_data_in_payload_49_real     (fft_col_in_payload_49_real[17:0]           ), //i
    .io_data_in_payload_49_imag     (fft_col_in_payload_49_imag[17:0]           ), //i
    .io_data_in_payload_50_real     (fft_col_in_payload_50_real[17:0]           ), //i
    .io_data_in_payload_50_imag     (fft_col_in_payload_50_imag[17:0]           ), //i
    .io_data_in_payload_51_real     (fft_col_in_payload_51_real[17:0]           ), //i
    .io_data_in_payload_51_imag     (fft_col_in_payload_51_imag[17:0]           ), //i
    .io_data_in_payload_52_real     (fft_col_in_payload_52_real[17:0]           ), //i
    .io_data_in_payload_52_imag     (fft_col_in_payload_52_imag[17:0]           ), //i
    .io_data_in_payload_53_real     (fft_col_in_payload_53_real[17:0]           ), //i
    .io_data_in_payload_53_imag     (fft_col_in_payload_53_imag[17:0]           ), //i
    .io_data_in_payload_54_real     (fft_col_in_payload_54_real[17:0]           ), //i
    .io_data_in_payload_54_imag     (fft_col_in_payload_54_imag[17:0]           ), //i
    .io_data_in_payload_55_real     (fft_col_in_payload_55_real[17:0]           ), //i
    .io_data_in_payload_55_imag     (fft_col_in_payload_55_imag[17:0]           ), //i
    .io_data_in_payload_56_real     (fft_col_in_payload_56_real[17:0]           ), //i
    .io_data_in_payload_56_imag     (fft_col_in_payload_56_imag[17:0]           ), //i
    .io_data_in_payload_57_real     (fft_col_in_payload_57_real[17:0]           ), //i
    .io_data_in_payload_57_imag     (fft_col_in_payload_57_imag[17:0]           ), //i
    .io_data_in_payload_58_real     (fft_col_in_payload_58_real[17:0]           ), //i
    .io_data_in_payload_58_imag     (fft_col_in_payload_58_imag[17:0]           ), //i
    .io_data_in_payload_59_real     (fft_col_in_payload_59_real[17:0]           ), //i
    .io_data_in_payload_59_imag     (fft_col_in_payload_59_imag[17:0]           ), //i
    .io_data_in_payload_60_real     (fft_col_in_payload_60_real[17:0]           ), //i
    .io_data_in_payload_60_imag     (fft_col_in_payload_60_imag[17:0]           ), //i
    .io_data_in_payload_61_real     (fft_col_in_payload_61_real[17:0]           ), //i
    .io_data_in_payload_61_imag     (fft_col_in_payload_61_imag[17:0]           ), //i
    .io_data_in_payload_62_real     (fft_col_in_payload_62_real[17:0]           ), //i
    .io_data_in_payload_62_imag     (fft_col_in_payload_62_imag[17:0]           ), //i
    .io_data_in_payload_63_real     (fft_col_in_payload_63_real[17:0]           ), //i
    .io_data_in_payload_63_imag     (fft_col_in_payload_63_imag[17:0]           ), //i
    .fft_col_out_valid              (myFFT_3_fft_col_out_valid                  ), //o
    .fft_col_out_payload_0_real     (myFFT_3_fft_col_out_payload_0_real[17:0]   ), //o
    .fft_col_out_payload_0_imag     (myFFT_3_fft_col_out_payload_0_imag[17:0]   ), //o
    .fft_col_out_payload_1_real     (myFFT_3_fft_col_out_payload_1_real[17:0]   ), //o
    .fft_col_out_payload_1_imag     (myFFT_3_fft_col_out_payload_1_imag[17:0]   ), //o
    .fft_col_out_payload_2_real     (myFFT_3_fft_col_out_payload_2_real[17:0]   ), //o
    .fft_col_out_payload_2_imag     (myFFT_3_fft_col_out_payload_2_imag[17:0]   ), //o
    .fft_col_out_payload_3_real     (myFFT_3_fft_col_out_payload_3_real[17:0]   ), //o
    .fft_col_out_payload_3_imag     (myFFT_3_fft_col_out_payload_3_imag[17:0]   ), //o
    .fft_col_out_payload_4_real     (myFFT_3_fft_col_out_payload_4_real[17:0]   ), //o
    .fft_col_out_payload_4_imag     (myFFT_3_fft_col_out_payload_4_imag[17:0]   ), //o
    .fft_col_out_payload_5_real     (myFFT_3_fft_col_out_payload_5_real[17:0]   ), //o
    .fft_col_out_payload_5_imag     (myFFT_3_fft_col_out_payload_5_imag[17:0]   ), //o
    .fft_col_out_payload_6_real     (myFFT_3_fft_col_out_payload_6_real[17:0]   ), //o
    .fft_col_out_payload_6_imag     (myFFT_3_fft_col_out_payload_6_imag[17:0]   ), //o
    .fft_col_out_payload_7_real     (myFFT_3_fft_col_out_payload_7_real[17:0]   ), //o
    .fft_col_out_payload_7_imag     (myFFT_3_fft_col_out_payload_7_imag[17:0]   ), //o
    .fft_col_out_payload_8_real     (myFFT_3_fft_col_out_payload_8_real[17:0]   ), //o
    .fft_col_out_payload_8_imag     (myFFT_3_fft_col_out_payload_8_imag[17:0]   ), //o
    .fft_col_out_payload_9_real     (myFFT_3_fft_col_out_payload_9_real[17:0]   ), //o
    .fft_col_out_payload_9_imag     (myFFT_3_fft_col_out_payload_9_imag[17:0]   ), //o
    .fft_col_out_payload_10_real    (myFFT_3_fft_col_out_payload_10_real[17:0]  ), //o
    .fft_col_out_payload_10_imag    (myFFT_3_fft_col_out_payload_10_imag[17:0]  ), //o
    .fft_col_out_payload_11_real    (myFFT_3_fft_col_out_payload_11_real[17:0]  ), //o
    .fft_col_out_payload_11_imag    (myFFT_3_fft_col_out_payload_11_imag[17:0]  ), //o
    .fft_col_out_payload_12_real    (myFFT_3_fft_col_out_payload_12_real[17:0]  ), //o
    .fft_col_out_payload_12_imag    (myFFT_3_fft_col_out_payload_12_imag[17:0]  ), //o
    .fft_col_out_payload_13_real    (myFFT_3_fft_col_out_payload_13_real[17:0]  ), //o
    .fft_col_out_payload_13_imag    (myFFT_3_fft_col_out_payload_13_imag[17:0]  ), //o
    .fft_col_out_payload_14_real    (myFFT_3_fft_col_out_payload_14_real[17:0]  ), //o
    .fft_col_out_payload_14_imag    (myFFT_3_fft_col_out_payload_14_imag[17:0]  ), //o
    .fft_col_out_payload_15_real    (myFFT_3_fft_col_out_payload_15_real[17:0]  ), //o
    .fft_col_out_payload_15_imag    (myFFT_3_fft_col_out_payload_15_imag[17:0]  ), //o
    .fft_col_out_payload_16_real    (myFFT_3_fft_col_out_payload_16_real[17:0]  ), //o
    .fft_col_out_payload_16_imag    (myFFT_3_fft_col_out_payload_16_imag[17:0]  ), //o
    .fft_col_out_payload_17_real    (myFFT_3_fft_col_out_payload_17_real[17:0]  ), //o
    .fft_col_out_payload_17_imag    (myFFT_3_fft_col_out_payload_17_imag[17:0]  ), //o
    .fft_col_out_payload_18_real    (myFFT_3_fft_col_out_payload_18_real[17:0]  ), //o
    .fft_col_out_payload_18_imag    (myFFT_3_fft_col_out_payload_18_imag[17:0]  ), //o
    .fft_col_out_payload_19_real    (myFFT_3_fft_col_out_payload_19_real[17:0]  ), //o
    .fft_col_out_payload_19_imag    (myFFT_3_fft_col_out_payload_19_imag[17:0]  ), //o
    .fft_col_out_payload_20_real    (myFFT_3_fft_col_out_payload_20_real[17:0]  ), //o
    .fft_col_out_payload_20_imag    (myFFT_3_fft_col_out_payload_20_imag[17:0]  ), //o
    .fft_col_out_payload_21_real    (myFFT_3_fft_col_out_payload_21_real[17:0]  ), //o
    .fft_col_out_payload_21_imag    (myFFT_3_fft_col_out_payload_21_imag[17:0]  ), //o
    .fft_col_out_payload_22_real    (myFFT_3_fft_col_out_payload_22_real[17:0]  ), //o
    .fft_col_out_payload_22_imag    (myFFT_3_fft_col_out_payload_22_imag[17:0]  ), //o
    .fft_col_out_payload_23_real    (myFFT_3_fft_col_out_payload_23_real[17:0]  ), //o
    .fft_col_out_payload_23_imag    (myFFT_3_fft_col_out_payload_23_imag[17:0]  ), //o
    .fft_col_out_payload_24_real    (myFFT_3_fft_col_out_payload_24_real[17:0]  ), //o
    .fft_col_out_payload_24_imag    (myFFT_3_fft_col_out_payload_24_imag[17:0]  ), //o
    .fft_col_out_payload_25_real    (myFFT_3_fft_col_out_payload_25_real[17:0]  ), //o
    .fft_col_out_payload_25_imag    (myFFT_3_fft_col_out_payload_25_imag[17:0]  ), //o
    .fft_col_out_payload_26_real    (myFFT_3_fft_col_out_payload_26_real[17:0]  ), //o
    .fft_col_out_payload_26_imag    (myFFT_3_fft_col_out_payload_26_imag[17:0]  ), //o
    .fft_col_out_payload_27_real    (myFFT_3_fft_col_out_payload_27_real[17:0]  ), //o
    .fft_col_out_payload_27_imag    (myFFT_3_fft_col_out_payload_27_imag[17:0]  ), //o
    .fft_col_out_payload_28_real    (myFFT_3_fft_col_out_payload_28_real[17:0]  ), //o
    .fft_col_out_payload_28_imag    (myFFT_3_fft_col_out_payload_28_imag[17:0]  ), //o
    .fft_col_out_payload_29_real    (myFFT_3_fft_col_out_payload_29_real[17:0]  ), //o
    .fft_col_out_payload_29_imag    (myFFT_3_fft_col_out_payload_29_imag[17:0]  ), //o
    .fft_col_out_payload_30_real    (myFFT_3_fft_col_out_payload_30_real[17:0]  ), //o
    .fft_col_out_payload_30_imag    (myFFT_3_fft_col_out_payload_30_imag[17:0]  ), //o
    .fft_col_out_payload_31_real    (myFFT_3_fft_col_out_payload_31_real[17:0]  ), //o
    .fft_col_out_payload_31_imag    (myFFT_3_fft_col_out_payload_31_imag[17:0]  ), //o
    .fft_col_out_payload_32_real    (myFFT_3_fft_col_out_payload_32_real[17:0]  ), //o
    .fft_col_out_payload_32_imag    (myFFT_3_fft_col_out_payload_32_imag[17:0]  ), //o
    .fft_col_out_payload_33_real    (myFFT_3_fft_col_out_payload_33_real[17:0]  ), //o
    .fft_col_out_payload_33_imag    (myFFT_3_fft_col_out_payload_33_imag[17:0]  ), //o
    .fft_col_out_payload_34_real    (myFFT_3_fft_col_out_payload_34_real[17:0]  ), //o
    .fft_col_out_payload_34_imag    (myFFT_3_fft_col_out_payload_34_imag[17:0]  ), //o
    .fft_col_out_payload_35_real    (myFFT_3_fft_col_out_payload_35_real[17:0]  ), //o
    .fft_col_out_payload_35_imag    (myFFT_3_fft_col_out_payload_35_imag[17:0]  ), //o
    .fft_col_out_payload_36_real    (myFFT_3_fft_col_out_payload_36_real[17:0]  ), //o
    .fft_col_out_payload_36_imag    (myFFT_3_fft_col_out_payload_36_imag[17:0]  ), //o
    .fft_col_out_payload_37_real    (myFFT_3_fft_col_out_payload_37_real[17:0]  ), //o
    .fft_col_out_payload_37_imag    (myFFT_3_fft_col_out_payload_37_imag[17:0]  ), //o
    .fft_col_out_payload_38_real    (myFFT_3_fft_col_out_payload_38_real[17:0]  ), //o
    .fft_col_out_payload_38_imag    (myFFT_3_fft_col_out_payload_38_imag[17:0]  ), //o
    .fft_col_out_payload_39_real    (myFFT_3_fft_col_out_payload_39_real[17:0]  ), //o
    .fft_col_out_payload_39_imag    (myFFT_3_fft_col_out_payload_39_imag[17:0]  ), //o
    .fft_col_out_payload_40_real    (myFFT_3_fft_col_out_payload_40_real[17:0]  ), //o
    .fft_col_out_payload_40_imag    (myFFT_3_fft_col_out_payload_40_imag[17:0]  ), //o
    .fft_col_out_payload_41_real    (myFFT_3_fft_col_out_payload_41_real[17:0]  ), //o
    .fft_col_out_payload_41_imag    (myFFT_3_fft_col_out_payload_41_imag[17:0]  ), //o
    .fft_col_out_payload_42_real    (myFFT_3_fft_col_out_payload_42_real[17:0]  ), //o
    .fft_col_out_payload_42_imag    (myFFT_3_fft_col_out_payload_42_imag[17:0]  ), //o
    .fft_col_out_payload_43_real    (myFFT_3_fft_col_out_payload_43_real[17:0]  ), //o
    .fft_col_out_payload_43_imag    (myFFT_3_fft_col_out_payload_43_imag[17:0]  ), //o
    .fft_col_out_payload_44_real    (myFFT_3_fft_col_out_payload_44_real[17:0]  ), //o
    .fft_col_out_payload_44_imag    (myFFT_3_fft_col_out_payload_44_imag[17:0]  ), //o
    .fft_col_out_payload_45_real    (myFFT_3_fft_col_out_payload_45_real[17:0]  ), //o
    .fft_col_out_payload_45_imag    (myFFT_3_fft_col_out_payload_45_imag[17:0]  ), //o
    .fft_col_out_payload_46_real    (myFFT_3_fft_col_out_payload_46_real[17:0]  ), //o
    .fft_col_out_payload_46_imag    (myFFT_3_fft_col_out_payload_46_imag[17:0]  ), //o
    .fft_col_out_payload_47_real    (myFFT_3_fft_col_out_payload_47_real[17:0]  ), //o
    .fft_col_out_payload_47_imag    (myFFT_3_fft_col_out_payload_47_imag[17:0]  ), //o
    .fft_col_out_payload_48_real    (myFFT_3_fft_col_out_payload_48_real[17:0]  ), //o
    .fft_col_out_payload_48_imag    (myFFT_3_fft_col_out_payload_48_imag[17:0]  ), //o
    .fft_col_out_payload_49_real    (myFFT_3_fft_col_out_payload_49_real[17:0]  ), //o
    .fft_col_out_payload_49_imag    (myFFT_3_fft_col_out_payload_49_imag[17:0]  ), //o
    .fft_col_out_payload_50_real    (myFFT_3_fft_col_out_payload_50_real[17:0]  ), //o
    .fft_col_out_payload_50_imag    (myFFT_3_fft_col_out_payload_50_imag[17:0]  ), //o
    .fft_col_out_payload_51_real    (myFFT_3_fft_col_out_payload_51_real[17:0]  ), //o
    .fft_col_out_payload_51_imag    (myFFT_3_fft_col_out_payload_51_imag[17:0]  ), //o
    .fft_col_out_payload_52_real    (myFFT_3_fft_col_out_payload_52_real[17:0]  ), //o
    .fft_col_out_payload_52_imag    (myFFT_3_fft_col_out_payload_52_imag[17:0]  ), //o
    .fft_col_out_payload_53_real    (myFFT_3_fft_col_out_payload_53_real[17:0]  ), //o
    .fft_col_out_payload_53_imag    (myFFT_3_fft_col_out_payload_53_imag[17:0]  ), //o
    .fft_col_out_payload_54_real    (myFFT_3_fft_col_out_payload_54_real[17:0]  ), //o
    .fft_col_out_payload_54_imag    (myFFT_3_fft_col_out_payload_54_imag[17:0]  ), //o
    .fft_col_out_payload_55_real    (myFFT_3_fft_col_out_payload_55_real[17:0]  ), //o
    .fft_col_out_payload_55_imag    (myFFT_3_fft_col_out_payload_55_imag[17:0]  ), //o
    .fft_col_out_payload_56_real    (myFFT_3_fft_col_out_payload_56_real[17:0]  ), //o
    .fft_col_out_payload_56_imag    (myFFT_3_fft_col_out_payload_56_imag[17:0]  ), //o
    .fft_col_out_payload_57_real    (myFFT_3_fft_col_out_payload_57_real[17:0]  ), //o
    .fft_col_out_payload_57_imag    (myFFT_3_fft_col_out_payload_57_imag[17:0]  ), //o
    .fft_col_out_payload_58_real    (myFFT_3_fft_col_out_payload_58_real[17:0]  ), //o
    .fft_col_out_payload_58_imag    (myFFT_3_fft_col_out_payload_58_imag[17:0]  ), //o
    .fft_col_out_payload_59_real    (myFFT_3_fft_col_out_payload_59_real[17:0]  ), //o
    .fft_col_out_payload_59_imag    (myFFT_3_fft_col_out_payload_59_imag[17:0]  ), //o
    .fft_col_out_payload_60_real    (myFFT_3_fft_col_out_payload_60_real[17:0]  ), //o
    .fft_col_out_payload_60_imag    (myFFT_3_fft_col_out_payload_60_imag[17:0]  ), //o
    .fft_col_out_payload_61_real    (myFFT_3_fft_col_out_payload_61_real[17:0]  ), //o
    .fft_col_out_payload_61_imag    (myFFT_3_fft_col_out_payload_61_imag[17:0]  ), //o
    .fft_col_out_payload_62_real    (myFFT_3_fft_col_out_payload_62_real[17:0]  ), //o
    .fft_col_out_payload_62_imag    (myFFT_3_fft_col_out_payload_62_imag[17:0]  ), //o
    .fft_col_out_payload_63_real    (myFFT_3_fft_col_out_payload_63_real[17:0]  ), //o
    .fft_col_out_payload_63_imag    (myFFT_3_fft_col_out_payload_63_imag[17:0]  ), //o
    .clk                            (clk                                        ), //i
    .reset                          (reset                                      )  //i
  );
  always @(*) begin
    case(col_addr)
      6'b000000 : begin
        _zz_194 = img_reg_array_0_0_real;
        _zz_195 = img_reg_array_0_0_imag;
        _zz_196 = img_reg_array_1_0_real;
        _zz_197 = img_reg_array_1_0_imag;
        _zz_198 = img_reg_array_2_0_real;
        _zz_199 = img_reg_array_2_0_imag;
        _zz_200 = img_reg_array_3_0_real;
        _zz_201 = img_reg_array_3_0_imag;
        _zz_202 = img_reg_array_4_0_real;
        _zz_203 = img_reg_array_4_0_imag;
        _zz_204 = img_reg_array_5_0_real;
        _zz_205 = img_reg_array_5_0_imag;
        _zz_206 = img_reg_array_6_0_real;
        _zz_207 = img_reg_array_6_0_imag;
        _zz_208 = img_reg_array_7_0_real;
        _zz_209 = img_reg_array_7_0_imag;
        _zz_210 = img_reg_array_8_0_real;
        _zz_211 = img_reg_array_8_0_imag;
        _zz_212 = img_reg_array_9_0_real;
        _zz_213 = img_reg_array_9_0_imag;
        _zz_214 = img_reg_array_10_0_real;
        _zz_215 = img_reg_array_10_0_imag;
        _zz_216 = img_reg_array_11_0_real;
        _zz_217 = img_reg_array_11_0_imag;
        _zz_218 = img_reg_array_12_0_real;
        _zz_219 = img_reg_array_12_0_imag;
        _zz_220 = img_reg_array_13_0_real;
        _zz_221 = img_reg_array_13_0_imag;
        _zz_222 = img_reg_array_14_0_real;
        _zz_223 = img_reg_array_14_0_imag;
        _zz_224 = img_reg_array_15_0_real;
        _zz_225 = img_reg_array_15_0_imag;
        _zz_226 = img_reg_array_16_0_real;
        _zz_227 = img_reg_array_16_0_imag;
        _zz_228 = img_reg_array_17_0_real;
        _zz_229 = img_reg_array_17_0_imag;
        _zz_230 = img_reg_array_18_0_real;
        _zz_231 = img_reg_array_18_0_imag;
        _zz_232 = img_reg_array_19_0_real;
        _zz_233 = img_reg_array_19_0_imag;
        _zz_234 = img_reg_array_20_0_real;
        _zz_235 = img_reg_array_20_0_imag;
        _zz_236 = img_reg_array_21_0_real;
        _zz_237 = img_reg_array_21_0_imag;
        _zz_238 = img_reg_array_22_0_real;
        _zz_239 = img_reg_array_22_0_imag;
        _zz_240 = img_reg_array_23_0_real;
        _zz_241 = img_reg_array_23_0_imag;
        _zz_242 = img_reg_array_24_0_real;
        _zz_243 = img_reg_array_24_0_imag;
        _zz_244 = img_reg_array_25_0_real;
        _zz_245 = img_reg_array_25_0_imag;
        _zz_246 = img_reg_array_26_0_real;
        _zz_247 = img_reg_array_26_0_imag;
        _zz_248 = img_reg_array_27_0_real;
        _zz_249 = img_reg_array_27_0_imag;
        _zz_250 = img_reg_array_28_0_real;
        _zz_251 = img_reg_array_28_0_imag;
        _zz_252 = img_reg_array_29_0_real;
        _zz_253 = img_reg_array_29_0_imag;
        _zz_254 = img_reg_array_30_0_real;
        _zz_255 = img_reg_array_30_0_imag;
        _zz_256 = img_reg_array_31_0_real;
        _zz_257 = img_reg_array_31_0_imag;
        _zz_258 = img_reg_array_32_0_real;
        _zz_259 = img_reg_array_32_0_imag;
        _zz_260 = img_reg_array_33_0_real;
        _zz_261 = img_reg_array_33_0_imag;
        _zz_262 = img_reg_array_34_0_real;
        _zz_263 = img_reg_array_34_0_imag;
        _zz_264 = img_reg_array_35_0_real;
        _zz_265 = img_reg_array_35_0_imag;
        _zz_266 = img_reg_array_36_0_real;
        _zz_267 = img_reg_array_36_0_imag;
        _zz_268 = img_reg_array_37_0_real;
        _zz_269 = img_reg_array_37_0_imag;
        _zz_270 = img_reg_array_38_0_real;
        _zz_271 = img_reg_array_38_0_imag;
        _zz_272 = img_reg_array_39_0_real;
        _zz_273 = img_reg_array_39_0_imag;
        _zz_274 = img_reg_array_40_0_real;
        _zz_275 = img_reg_array_40_0_imag;
        _zz_276 = img_reg_array_41_0_real;
        _zz_277 = img_reg_array_41_0_imag;
        _zz_278 = img_reg_array_42_0_real;
        _zz_279 = img_reg_array_42_0_imag;
        _zz_280 = img_reg_array_43_0_real;
        _zz_281 = img_reg_array_43_0_imag;
        _zz_282 = img_reg_array_44_0_real;
        _zz_283 = img_reg_array_44_0_imag;
        _zz_284 = img_reg_array_45_0_real;
        _zz_285 = img_reg_array_45_0_imag;
        _zz_286 = img_reg_array_46_0_real;
        _zz_287 = img_reg_array_46_0_imag;
        _zz_288 = img_reg_array_47_0_real;
        _zz_289 = img_reg_array_47_0_imag;
        _zz_290 = img_reg_array_48_0_real;
        _zz_291 = img_reg_array_48_0_imag;
        _zz_292 = img_reg_array_49_0_real;
        _zz_293 = img_reg_array_49_0_imag;
        _zz_294 = img_reg_array_50_0_real;
        _zz_295 = img_reg_array_50_0_imag;
        _zz_296 = img_reg_array_51_0_real;
        _zz_297 = img_reg_array_51_0_imag;
        _zz_298 = img_reg_array_52_0_real;
        _zz_299 = img_reg_array_52_0_imag;
        _zz_300 = img_reg_array_53_0_real;
        _zz_301 = img_reg_array_53_0_imag;
        _zz_302 = img_reg_array_54_0_real;
        _zz_303 = img_reg_array_54_0_imag;
        _zz_304 = img_reg_array_55_0_real;
        _zz_305 = img_reg_array_55_0_imag;
        _zz_306 = img_reg_array_56_0_real;
        _zz_307 = img_reg_array_56_0_imag;
        _zz_308 = img_reg_array_57_0_real;
        _zz_309 = img_reg_array_57_0_imag;
        _zz_310 = img_reg_array_58_0_real;
        _zz_311 = img_reg_array_58_0_imag;
        _zz_312 = img_reg_array_59_0_real;
        _zz_313 = img_reg_array_59_0_imag;
        _zz_314 = img_reg_array_60_0_real;
        _zz_315 = img_reg_array_60_0_imag;
        _zz_316 = img_reg_array_61_0_real;
        _zz_317 = img_reg_array_61_0_imag;
        _zz_318 = img_reg_array_62_0_real;
        _zz_319 = img_reg_array_62_0_imag;
        _zz_320 = img_reg_array_63_0_real;
        _zz_321 = img_reg_array_63_0_imag;
      end
      6'b000001 : begin
        _zz_194 = img_reg_array_0_1_real;
        _zz_195 = img_reg_array_0_1_imag;
        _zz_196 = img_reg_array_1_1_real;
        _zz_197 = img_reg_array_1_1_imag;
        _zz_198 = img_reg_array_2_1_real;
        _zz_199 = img_reg_array_2_1_imag;
        _zz_200 = img_reg_array_3_1_real;
        _zz_201 = img_reg_array_3_1_imag;
        _zz_202 = img_reg_array_4_1_real;
        _zz_203 = img_reg_array_4_1_imag;
        _zz_204 = img_reg_array_5_1_real;
        _zz_205 = img_reg_array_5_1_imag;
        _zz_206 = img_reg_array_6_1_real;
        _zz_207 = img_reg_array_6_1_imag;
        _zz_208 = img_reg_array_7_1_real;
        _zz_209 = img_reg_array_7_1_imag;
        _zz_210 = img_reg_array_8_1_real;
        _zz_211 = img_reg_array_8_1_imag;
        _zz_212 = img_reg_array_9_1_real;
        _zz_213 = img_reg_array_9_1_imag;
        _zz_214 = img_reg_array_10_1_real;
        _zz_215 = img_reg_array_10_1_imag;
        _zz_216 = img_reg_array_11_1_real;
        _zz_217 = img_reg_array_11_1_imag;
        _zz_218 = img_reg_array_12_1_real;
        _zz_219 = img_reg_array_12_1_imag;
        _zz_220 = img_reg_array_13_1_real;
        _zz_221 = img_reg_array_13_1_imag;
        _zz_222 = img_reg_array_14_1_real;
        _zz_223 = img_reg_array_14_1_imag;
        _zz_224 = img_reg_array_15_1_real;
        _zz_225 = img_reg_array_15_1_imag;
        _zz_226 = img_reg_array_16_1_real;
        _zz_227 = img_reg_array_16_1_imag;
        _zz_228 = img_reg_array_17_1_real;
        _zz_229 = img_reg_array_17_1_imag;
        _zz_230 = img_reg_array_18_1_real;
        _zz_231 = img_reg_array_18_1_imag;
        _zz_232 = img_reg_array_19_1_real;
        _zz_233 = img_reg_array_19_1_imag;
        _zz_234 = img_reg_array_20_1_real;
        _zz_235 = img_reg_array_20_1_imag;
        _zz_236 = img_reg_array_21_1_real;
        _zz_237 = img_reg_array_21_1_imag;
        _zz_238 = img_reg_array_22_1_real;
        _zz_239 = img_reg_array_22_1_imag;
        _zz_240 = img_reg_array_23_1_real;
        _zz_241 = img_reg_array_23_1_imag;
        _zz_242 = img_reg_array_24_1_real;
        _zz_243 = img_reg_array_24_1_imag;
        _zz_244 = img_reg_array_25_1_real;
        _zz_245 = img_reg_array_25_1_imag;
        _zz_246 = img_reg_array_26_1_real;
        _zz_247 = img_reg_array_26_1_imag;
        _zz_248 = img_reg_array_27_1_real;
        _zz_249 = img_reg_array_27_1_imag;
        _zz_250 = img_reg_array_28_1_real;
        _zz_251 = img_reg_array_28_1_imag;
        _zz_252 = img_reg_array_29_1_real;
        _zz_253 = img_reg_array_29_1_imag;
        _zz_254 = img_reg_array_30_1_real;
        _zz_255 = img_reg_array_30_1_imag;
        _zz_256 = img_reg_array_31_1_real;
        _zz_257 = img_reg_array_31_1_imag;
        _zz_258 = img_reg_array_32_1_real;
        _zz_259 = img_reg_array_32_1_imag;
        _zz_260 = img_reg_array_33_1_real;
        _zz_261 = img_reg_array_33_1_imag;
        _zz_262 = img_reg_array_34_1_real;
        _zz_263 = img_reg_array_34_1_imag;
        _zz_264 = img_reg_array_35_1_real;
        _zz_265 = img_reg_array_35_1_imag;
        _zz_266 = img_reg_array_36_1_real;
        _zz_267 = img_reg_array_36_1_imag;
        _zz_268 = img_reg_array_37_1_real;
        _zz_269 = img_reg_array_37_1_imag;
        _zz_270 = img_reg_array_38_1_real;
        _zz_271 = img_reg_array_38_1_imag;
        _zz_272 = img_reg_array_39_1_real;
        _zz_273 = img_reg_array_39_1_imag;
        _zz_274 = img_reg_array_40_1_real;
        _zz_275 = img_reg_array_40_1_imag;
        _zz_276 = img_reg_array_41_1_real;
        _zz_277 = img_reg_array_41_1_imag;
        _zz_278 = img_reg_array_42_1_real;
        _zz_279 = img_reg_array_42_1_imag;
        _zz_280 = img_reg_array_43_1_real;
        _zz_281 = img_reg_array_43_1_imag;
        _zz_282 = img_reg_array_44_1_real;
        _zz_283 = img_reg_array_44_1_imag;
        _zz_284 = img_reg_array_45_1_real;
        _zz_285 = img_reg_array_45_1_imag;
        _zz_286 = img_reg_array_46_1_real;
        _zz_287 = img_reg_array_46_1_imag;
        _zz_288 = img_reg_array_47_1_real;
        _zz_289 = img_reg_array_47_1_imag;
        _zz_290 = img_reg_array_48_1_real;
        _zz_291 = img_reg_array_48_1_imag;
        _zz_292 = img_reg_array_49_1_real;
        _zz_293 = img_reg_array_49_1_imag;
        _zz_294 = img_reg_array_50_1_real;
        _zz_295 = img_reg_array_50_1_imag;
        _zz_296 = img_reg_array_51_1_real;
        _zz_297 = img_reg_array_51_1_imag;
        _zz_298 = img_reg_array_52_1_real;
        _zz_299 = img_reg_array_52_1_imag;
        _zz_300 = img_reg_array_53_1_real;
        _zz_301 = img_reg_array_53_1_imag;
        _zz_302 = img_reg_array_54_1_real;
        _zz_303 = img_reg_array_54_1_imag;
        _zz_304 = img_reg_array_55_1_real;
        _zz_305 = img_reg_array_55_1_imag;
        _zz_306 = img_reg_array_56_1_real;
        _zz_307 = img_reg_array_56_1_imag;
        _zz_308 = img_reg_array_57_1_real;
        _zz_309 = img_reg_array_57_1_imag;
        _zz_310 = img_reg_array_58_1_real;
        _zz_311 = img_reg_array_58_1_imag;
        _zz_312 = img_reg_array_59_1_real;
        _zz_313 = img_reg_array_59_1_imag;
        _zz_314 = img_reg_array_60_1_real;
        _zz_315 = img_reg_array_60_1_imag;
        _zz_316 = img_reg_array_61_1_real;
        _zz_317 = img_reg_array_61_1_imag;
        _zz_318 = img_reg_array_62_1_real;
        _zz_319 = img_reg_array_62_1_imag;
        _zz_320 = img_reg_array_63_1_real;
        _zz_321 = img_reg_array_63_1_imag;
      end
      6'b000010 : begin
        _zz_194 = img_reg_array_0_2_real;
        _zz_195 = img_reg_array_0_2_imag;
        _zz_196 = img_reg_array_1_2_real;
        _zz_197 = img_reg_array_1_2_imag;
        _zz_198 = img_reg_array_2_2_real;
        _zz_199 = img_reg_array_2_2_imag;
        _zz_200 = img_reg_array_3_2_real;
        _zz_201 = img_reg_array_3_2_imag;
        _zz_202 = img_reg_array_4_2_real;
        _zz_203 = img_reg_array_4_2_imag;
        _zz_204 = img_reg_array_5_2_real;
        _zz_205 = img_reg_array_5_2_imag;
        _zz_206 = img_reg_array_6_2_real;
        _zz_207 = img_reg_array_6_2_imag;
        _zz_208 = img_reg_array_7_2_real;
        _zz_209 = img_reg_array_7_2_imag;
        _zz_210 = img_reg_array_8_2_real;
        _zz_211 = img_reg_array_8_2_imag;
        _zz_212 = img_reg_array_9_2_real;
        _zz_213 = img_reg_array_9_2_imag;
        _zz_214 = img_reg_array_10_2_real;
        _zz_215 = img_reg_array_10_2_imag;
        _zz_216 = img_reg_array_11_2_real;
        _zz_217 = img_reg_array_11_2_imag;
        _zz_218 = img_reg_array_12_2_real;
        _zz_219 = img_reg_array_12_2_imag;
        _zz_220 = img_reg_array_13_2_real;
        _zz_221 = img_reg_array_13_2_imag;
        _zz_222 = img_reg_array_14_2_real;
        _zz_223 = img_reg_array_14_2_imag;
        _zz_224 = img_reg_array_15_2_real;
        _zz_225 = img_reg_array_15_2_imag;
        _zz_226 = img_reg_array_16_2_real;
        _zz_227 = img_reg_array_16_2_imag;
        _zz_228 = img_reg_array_17_2_real;
        _zz_229 = img_reg_array_17_2_imag;
        _zz_230 = img_reg_array_18_2_real;
        _zz_231 = img_reg_array_18_2_imag;
        _zz_232 = img_reg_array_19_2_real;
        _zz_233 = img_reg_array_19_2_imag;
        _zz_234 = img_reg_array_20_2_real;
        _zz_235 = img_reg_array_20_2_imag;
        _zz_236 = img_reg_array_21_2_real;
        _zz_237 = img_reg_array_21_2_imag;
        _zz_238 = img_reg_array_22_2_real;
        _zz_239 = img_reg_array_22_2_imag;
        _zz_240 = img_reg_array_23_2_real;
        _zz_241 = img_reg_array_23_2_imag;
        _zz_242 = img_reg_array_24_2_real;
        _zz_243 = img_reg_array_24_2_imag;
        _zz_244 = img_reg_array_25_2_real;
        _zz_245 = img_reg_array_25_2_imag;
        _zz_246 = img_reg_array_26_2_real;
        _zz_247 = img_reg_array_26_2_imag;
        _zz_248 = img_reg_array_27_2_real;
        _zz_249 = img_reg_array_27_2_imag;
        _zz_250 = img_reg_array_28_2_real;
        _zz_251 = img_reg_array_28_2_imag;
        _zz_252 = img_reg_array_29_2_real;
        _zz_253 = img_reg_array_29_2_imag;
        _zz_254 = img_reg_array_30_2_real;
        _zz_255 = img_reg_array_30_2_imag;
        _zz_256 = img_reg_array_31_2_real;
        _zz_257 = img_reg_array_31_2_imag;
        _zz_258 = img_reg_array_32_2_real;
        _zz_259 = img_reg_array_32_2_imag;
        _zz_260 = img_reg_array_33_2_real;
        _zz_261 = img_reg_array_33_2_imag;
        _zz_262 = img_reg_array_34_2_real;
        _zz_263 = img_reg_array_34_2_imag;
        _zz_264 = img_reg_array_35_2_real;
        _zz_265 = img_reg_array_35_2_imag;
        _zz_266 = img_reg_array_36_2_real;
        _zz_267 = img_reg_array_36_2_imag;
        _zz_268 = img_reg_array_37_2_real;
        _zz_269 = img_reg_array_37_2_imag;
        _zz_270 = img_reg_array_38_2_real;
        _zz_271 = img_reg_array_38_2_imag;
        _zz_272 = img_reg_array_39_2_real;
        _zz_273 = img_reg_array_39_2_imag;
        _zz_274 = img_reg_array_40_2_real;
        _zz_275 = img_reg_array_40_2_imag;
        _zz_276 = img_reg_array_41_2_real;
        _zz_277 = img_reg_array_41_2_imag;
        _zz_278 = img_reg_array_42_2_real;
        _zz_279 = img_reg_array_42_2_imag;
        _zz_280 = img_reg_array_43_2_real;
        _zz_281 = img_reg_array_43_2_imag;
        _zz_282 = img_reg_array_44_2_real;
        _zz_283 = img_reg_array_44_2_imag;
        _zz_284 = img_reg_array_45_2_real;
        _zz_285 = img_reg_array_45_2_imag;
        _zz_286 = img_reg_array_46_2_real;
        _zz_287 = img_reg_array_46_2_imag;
        _zz_288 = img_reg_array_47_2_real;
        _zz_289 = img_reg_array_47_2_imag;
        _zz_290 = img_reg_array_48_2_real;
        _zz_291 = img_reg_array_48_2_imag;
        _zz_292 = img_reg_array_49_2_real;
        _zz_293 = img_reg_array_49_2_imag;
        _zz_294 = img_reg_array_50_2_real;
        _zz_295 = img_reg_array_50_2_imag;
        _zz_296 = img_reg_array_51_2_real;
        _zz_297 = img_reg_array_51_2_imag;
        _zz_298 = img_reg_array_52_2_real;
        _zz_299 = img_reg_array_52_2_imag;
        _zz_300 = img_reg_array_53_2_real;
        _zz_301 = img_reg_array_53_2_imag;
        _zz_302 = img_reg_array_54_2_real;
        _zz_303 = img_reg_array_54_2_imag;
        _zz_304 = img_reg_array_55_2_real;
        _zz_305 = img_reg_array_55_2_imag;
        _zz_306 = img_reg_array_56_2_real;
        _zz_307 = img_reg_array_56_2_imag;
        _zz_308 = img_reg_array_57_2_real;
        _zz_309 = img_reg_array_57_2_imag;
        _zz_310 = img_reg_array_58_2_real;
        _zz_311 = img_reg_array_58_2_imag;
        _zz_312 = img_reg_array_59_2_real;
        _zz_313 = img_reg_array_59_2_imag;
        _zz_314 = img_reg_array_60_2_real;
        _zz_315 = img_reg_array_60_2_imag;
        _zz_316 = img_reg_array_61_2_real;
        _zz_317 = img_reg_array_61_2_imag;
        _zz_318 = img_reg_array_62_2_real;
        _zz_319 = img_reg_array_62_2_imag;
        _zz_320 = img_reg_array_63_2_real;
        _zz_321 = img_reg_array_63_2_imag;
      end
      6'b000011 : begin
        _zz_194 = img_reg_array_0_3_real;
        _zz_195 = img_reg_array_0_3_imag;
        _zz_196 = img_reg_array_1_3_real;
        _zz_197 = img_reg_array_1_3_imag;
        _zz_198 = img_reg_array_2_3_real;
        _zz_199 = img_reg_array_2_3_imag;
        _zz_200 = img_reg_array_3_3_real;
        _zz_201 = img_reg_array_3_3_imag;
        _zz_202 = img_reg_array_4_3_real;
        _zz_203 = img_reg_array_4_3_imag;
        _zz_204 = img_reg_array_5_3_real;
        _zz_205 = img_reg_array_5_3_imag;
        _zz_206 = img_reg_array_6_3_real;
        _zz_207 = img_reg_array_6_3_imag;
        _zz_208 = img_reg_array_7_3_real;
        _zz_209 = img_reg_array_7_3_imag;
        _zz_210 = img_reg_array_8_3_real;
        _zz_211 = img_reg_array_8_3_imag;
        _zz_212 = img_reg_array_9_3_real;
        _zz_213 = img_reg_array_9_3_imag;
        _zz_214 = img_reg_array_10_3_real;
        _zz_215 = img_reg_array_10_3_imag;
        _zz_216 = img_reg_array_11_3_real;
        _zz_217 = img_reg_array_11_3_imag;
        _zz_218 = img_reg_array_12_3_real;
        _zz_219 = img_reg_array_12_3_imag;
        _zz_220 = img_reg_array_13_3_real;
        _zz_221 = img_reg_array_13_3_imag;
        _zz_222 = img_reg_array_14_3_real;
        _zz_223 = img_reg_array_14_3_imag;
        _zz_224 = img_reg_array_15_3_real;
        _zz_225 = img_reg_array_15_3_imag;
        _zz_226 = img_reg_array_16_3_real;
        _zz_227 = img_reg_array_16_3_imag;
        _zz_228 = img_reg_array_17_3_real;
        _zz_229 = img_reg_array_17_3_imag;
        _zz_230 = img_reg_array_18_3_real;
        _zz_231 = img_reg_array_18_3_imag;
        _zz_232 = img_reg_array_19_3_real;
        _zz_233 = img_reg_array_19_3_imag;
        _zz_234 = img_reg_array_20_3_real;
        _zz_235 = img_reg_array_20_3_imag;
        _zz_236 = img_reg_array_21_3_real;
        _zz_237 = img_reg_array_21_3_imag;
        _zz_238 = img_reg_array_22_3_real;
        _zz_239 = img_reg_array_22_3_imag;
        _zz_240 = img_reg_array_23_3_real;
        _zz_241 = img_reg_array_23_3_imag;
        _zz_242 = img_reg_array_24_3_real;
        _zz_243 = img_reg_array_24_3_imag;
        _zz_244 = img_reg_array_25_3_real;
        _zz_245 = img_reg_array_25_3_imag;
        _zz_246 = img_reg_array_26_3_real;
        _zz_247 = img_reg_array_26_3_imag;
        _zz_248 = img_reg_array_27_3_real;
        _zz_249 = img_reg_array_27_3_imag;
        _zz_250 = img_reg_array_28_3_real;
        _zz_251 = img_reg_array_28_3_imag;
        _zz_252 = img_reg_array_29_3_real;
        _zz_253 = img_reg_array_29_3_imag;
        _zz_254 = img_reg_array_30_3_real;
        _zz_255 = img_reg_array_30_3_imag;
        _zz_256 = img_reg_array_31_3_real;
        _zz_257 = img_reg_array_31_3_imag;
        _zz_258 = img_reg_array_32_3_real;
        _zz_259 = img_reg_array_32_3_imag;
        _zz_260 = img_reg_array_33_3_real;
        _zz_261 = img_reg_array_33_3_imag;
        _zz_262 = img_reg_array_34_3_real;
        _zz_263 = img_reg_array_34_3_imag;
        _zz_264 = img_reg_array_35_3_real;
        _zz_265 = img_reg_array_35_3_imag;
        _zz_266 = img_reg_array_36_3_real;
        _zz_267 = img_reg_array_36_3_imag;
        _zz_268 = img_reg_array_37_3_real;
        _zz_269 = img_reg_array_37_3_imag;
        _zz_270 = img_reg_array_38_3_real;
        _zz_271 = img_reg_array_38_3_imag;
        _zz_272 = img_reg_array_39_3_real;
        _zz_273 = img_reg_array_39_3_imag;
        _zz_274 = img_reg_array_40_3_real;
        _zz_275 = img_reg_array_40_3_imag;
        _zz_276 = img_reg_array_41_3_real;
        _zz_277 = img_reg_array_41_3_imag;
        _zz_278 = img_reg_array_42_3_real;
        _zz_279 = img_reg_array_42_3_imag;
        _zz_280 = img_reg_array_43_3_real;
        _zz_281 = img_reg_array_43_3_imag;
        _zz_282 = img_reg_array_44_3_real;
        _zz_283 = img_reg_array_44_3_imag;
        _zz_284 = img_reg_array_45_3_real;
        _zz_285 = img_reg_array_45_3_imag;
        _zz_286 = img_reg_array_46_3_real;
        _zz_287 = img_reg_array_46_3_imag;
        _zz_288 = img_reg_array_47_3_real;
        _zz_289 = img_reg_array_47_3_imag;
        _zz_290 = img_reg_array_48_3_real;
        _zz_291 = img_reg_array_48_3_imag;
        _zz_292 = img_reg_array_49_3_real;
        _zz_293 = img_reg_array_49_3_imag;
        _zz_294 = img_reg_array_50_3_real;
        _zz_295 = img_reg_array_50_3_imag;
        _zz_296 = img_reg_array_51_3_real;
        _zz_297 = img_reg_array_51_3_imag;
        _zz_298 = img_reg_array_52_3_real;
        _zz_299 = img_reg_array_52_3_imag;
        _zz_300 = img_reg_array_53_3_real;
        _zz_301 = img_reg_array_53_3_imag;
        _zz_302 = img_reg_array_54_3_real;
        _zz_303 = img_reg_array_54_3_imag;
        _zz_304 = img_reg_array_55_3_real;
        _zz_305 = img_reg_array_55_3_imag;
        _zz_306 = img_reg_array_56_3_real;
        _zz_307 = img_reg_array_56_3_imag;
        _zz_308 = img_reg_array_57_3_real;
        _zz_309 = img_reg_array_57_3_imag;
        _zz_310 = img_reg_array_58_3_real;
        _zz_311 = img_reg_array_58_3_imag;
        _zz_312 = img_reg_array_59_3_real;
        _zz_313 = img_reg_array_59_3_imag;
        _zz_314 = img_reg_array_60_3_real;
        _zz_315 = img_reg_array_60_3_imag;
        _zz_316 = img_reg_array_61_3_real;
        _zz_317 = img_reg_array_61_3_imag;
        _zz_318 = img_reg_array_62_3_real;
        _zz_319 = img_reg_array_62_3_imag;
        _zz_320 = img_reg_array_63_3_real;
        _zz_321 = img_reg_array_63_3_imag;
      end
      6'b000100 : begin
        _zz_194 = img_reg_array_0_4_real;
        _zz_195 = img_reg_array_0_4_imag;
        _zz_196 = img_reg_array_1_4_real;
        _zz_197 = img_reg_array_1_4_imag;
        _zz_198 = img_reg_array_2_4_real;
        _zz_199 = img_reg_array_2_4_imag;
        _zz_200 = img_reg_array_3_4_real;
        _zz_201 = img_reg_array_3_4_imag;
        _zz_202 = img_reg_array_4_4_real;
        _zz_203 = img_reg_array_4_4_imag;
        _zz_204 = img_reg_array_5_4_real;
        _zz_205 = img_reg_array_5_4_imag;
        _zz_206 = img_reg_array_6_4_real;
        _zz_207 = img_reg_array_6_4_imag;
        _zz_208 = img_reg_array_7_4_real;
        _zz_209 = img_reg_array_7_4_imag;
        _zz_210 = img_reg_array_8_4_real;
        _zz_211 = img_reg_array_8_4_imag;
        _zz_212 = img_reg_array_9_4_real;
        _zz_213 = img_reg_array_9_4_imag;
        _zz_214 = img_reg_array_10_4_real;
        _zz_215 = img_reg_array_10_4_imag;
        _zz_216 = img_reg_array_11_4_real;
        _zz_217 = img_reg_array_11_4_imag;
        _zz_218 = img_reg_array_12_4_real;
        _zz_219 = img_reg_array_12_4_imag;
        _zz_220 = img_reg_array_13_4_real;
        _zz_221 = img_reg_array_13_4_imag;
        _zz_222 = img_reg_array_14_4_real;
        _zz_223 = img_reg_array_14_4_imag;
        _zz_224 = img_reg_array_15_4_real;
        _zz_225 = img_reg_array_15_4_imag;
        _zz_226 = img_reg_array_16_4_real;
        _zz_227 = img_reg_array_16_4_imag;
        _zz_228 = img_reg_array_17_4_real;
        _zz_229 = img_reg_array_17_4_imag;
        _zz_230 = img_reg_array_18_4_real;
        _zz_231 = img_reg_array_18_4_imag;
        _zz_232 = img_reg_array_19_4_real;
        _zz_233 = img_reg_array_19_4_imag;
        _zz_234 = img_reg_array_20_4_real;
        _zz_235 = img_reg_array_20_4_imag;
        _zz_236 = img_reg_array_21_4_real;
        _zz_237 = img_reg_array_21_4_imag;
        _zz_238 = img_reg_array_22_4_real;
        _zz_239 = img_reg_array_22_4_imag;
        _zz_240 = img_reg_array_23_4_real;
        _zz_241 = img_reg_array_23_4_imag;
        _zz_242 = img_reg_array_24_4_real;
        _zz_243 = img_reg_array_24_4_imag;
        _zz_244 = img_reg_array_25_4_real;
        _zz_245 = img_reg_array_25_4_imag;
        _zz_246 = img_reg_array_26_4_real;
        _zz_247 = img_reg_array_26_4_imag;
        _zz_248 = img_reg_array_27_4_real;
        _zz_249 = img_reg_array_27_4_imag;
        _zz_250 = img_reg_array_28_4_real;
        _zz_251 = img_reg_array_28_4_imag;
        _zz_252 = img_reg_array_29_4_real;
        _zz_253 = img_reg_array_29_4_imag;
        _zz_254 = img_reg_array_30_4_real;
        _zz_255 = img_reg_array_30_4_imag;
        _zz_256 = img_reg_array_31_4_real;
        _zz_257 = img_reg_array_31_4_imag;
        _zz_258 = img_reg_array_32_4_real;
        _zz_259 = img_reg_array_32_4_imag;
        _zz_260 = img_reg_array_33_4_real;
        _zz_261 = img_reg_array_33_4_imag;
        _zz_262 = img_reg_array_34_4_real;
        _zz_263 = img_reg_array_34_4_imag;
        _zz_264 = img_reg_array_35_4_real;
        _zz_265 = img_reg_array_35_4_imag;
        _zz_266 = img_reg_array_36_4_real;
        _zz_267 = img_reg_array_36_4_imag;
        _zz_268 = img_reg_array_37_4_real;
        _zz_269 = img_reg_array_37_4_imag;
        _zz_270 = img_reg_array_38_4_real;
        _zz_271 = img_reg_array_38_4_imag;
        _zz_272 = img_reg_array_39_4_real;
        _zz_273 = img_reg_array_39_4_imag;
        _zz_274 = img_reg_array_40_4_real;
        _zz_275 = img_reg_array_40_4_imag;
        _zz_276 = img_reg_array_41_4_real;
        _zz_277 = img_reg_array_41_4_imag;
        _zz_278 = img_reg_array_42_4_real;
        _zz_279 = img_reg_array_42_4_imag;
        _zz_280 = img_reg_array_43_4_real;
        _zz_281 = img_reg_array_43_4_imag;
        _zz_282 = img_reg_array_44_4_real;
        _zz_283 = img_reg_array_44_4_imag;
        _zz_284 = img_reg_array_45_4_real;
        _zz_285 = img_reg_array_45_4_imag;
        _zz_286 = img_reg_array_46_4_real;
        _zz_287 = img_reg_array_46_4_imag;
        _zz_288 = img_reg_array_47_4_real;
        _zz_289 = img_reg_array_47_4_imag;
        _zz_290 = img_reg_array_48_4_real;
        _zz_291 = img_reg_array_48_4_imag;
        _zz_292 = img_reg_array_49_4_real;
        _zz_293 = img_reg_array_49_4_imag;
        _zz_294 = img_reg_array_50_4_real;
        _zz_295 = img_reg_array_50_4_imag;
        _zz_296 = img_reg_array_51_4_real;
        _zz_297 = img_reg_array_51_4_imag;
        _zz_298 = img_reg_array_52_4_real;
        _zz_299 = img_reg_array_52_4_imag;
        _zz_300 = img_reg_array_53_4_real;
        _zz_301 = img_reg_array_53_4_imag;
        _zz_302 = img_reg_array_54_4_real;
        _zz_303 = img_reg_array_54_4_imag;
        _zz_304 = img_reg_array_55_4_real;
        _zz_305 = img_reg_array_55_4_imag;
        _zz_306 = img_reg_array_56_4_real;
        _zz_307 = img_reg_array_56_4_imag;
        _zz_308 = img_reg_array_57_4_real;
        _zz_309 = img_reg_array_57_4_imag;
        _zz_310 = img_reg_array_58_4_real;
        _zz_311 = img_reg_array_58_4_imag;
        _zz_312 = img_reg_array_59_4_real;
        _zz_313 = img_reg_array_59_4_imag;
        _zz_314 = img_reg_array_60_4_real;
        _zz_315 = img_reg_array_60_4_imag;
        _zz_316 = img_reg_array_61_4_real;
        _zz_317 = img_reg_array_61_4_imag;
        _zz_318 = img_reg_array_62_4_real;
        _zz_319 = img_reg_array_62_4_imag;
        _zz_320 = img_reg_array_63_4_real;
        _zz_321 = img_reg_array_63_4_imag;
      end
      6'b000101 : begin
        _zz_194 = img_reg_array_0_5_real;
        _zz_195 = img_reg_array_0_5_imag;
        _zz_196 = img_reg_array_1_5_real;
        _zz_197 = img_reg_array_1_5_imag;
        _zz_198 = img_reg_array_2_5_real;
        _zz_199 = img_reg_array_2_5_imag;
        _zz_200 = img_reg_array_3_5_real;
        _zz_201 = img_reg_array_3_5_imag;
        _zz_202 = img_reg_array_4_5_real;
        _zz_203 = img_reg_array_4_5_imag;
        _zz_204 = img_reg_array_5_5_real;
        _zz_205 = img_reg_array_5_5_imag;
        _zz_206 = img_reg_array_6_5_real;
        _zz_207 = img_reg_array_6_5_imag;
        _zz_208 = img_reg_array_7_5_real;
        _zz_209 = img_reg_array_7_5_imag;
        _zz_210 = img_reg_array_8_5_real;
        _zz_211 = img_reg_array_8_5_imag;
        _zz_212 = img_reg_array_9_5_real;
        _zz_213 = img_reg_array_9_5_imag;
        _zz_214 = img_reg_array_10_5_real;
        _zz_215 = img_reg_array_10_5_imag;
        _zz_216 = img_reg_array_11_5_real;
        _zz_217 = img_reg_array_11_5_imag;
        _zz_218 = img_reg_array_12_5_real;
        _zz_219 = img_reg_array_12_5_imag;
        _zz_220 = img_reg_array_13_5_real;
        _zz_221 = img_reg_array_13_5_imag;
        _zz_222 = img_reg_array_14_5_real;
        _zz_223 = img_reg_array_14_5_imag;
        _zz_224 = img_reg_array_15_5_real;
        _zz_225 = img_reg_array_15_5_imag;
        _zz_226 = img_reg_array_16_5_real;
        _zz_227 = img_reg_array_16_5_imag;
        _zz_228 = img_reg_array_17_5_real;
        _zz_229 = img_reg_array_17_5_imag;
        _zz_230 = img_reg_array_18_5_real;
        _zz_231 = img_reg_array_18_5_imag;
        _zz_232 = img_reg_array_19_5_real;
        _zz_233 = img_reg_array_19_5_imag;
        _zz_234 = img_reg_array_20_5_real;
        _zz_235 = img_reg_array_20_5_imag;
        _zz_236 = img_reg_array_21_5_real;
        _zz_237 = img_reg_array_21_5_imag;
        _zz_238 = img_reg_array_22_5_real;
        _zz_239 = img_reg_array_22_5_imag;
        _zz_240 = img_reg_array_23_5_real;
        _zz_241 = img_reg_array_23_5_imag;
        _zz_242 = img_reg_array_24_5_real;
        _zz_243 = img_reg_array_24_5_imag;
        _zz_244 = img_reg_array_25_5_real;
        _zz_245 = img_reg_array_25_5_imag;
        _zz_246 = img_reg_array_26_5_real;
        _zz_247 = img_reg_array_26_5_imag;
        _zz_248 = img_reg_array_27_5_real;
        _zz_249 = img_reg_array_27_5_imag;
        _zz_250 = img_reg_array_28_5_real;
        _zz_251 = img_reg_array_28_5_imag;
        _zz_252 = img_reg_array_29_5_real;
        _zz_253 = img_reg_array_29_5_imag;
        _zz_254 = img_reg_array_30_5_real;
        _zz_255 = img_reg_array_30_5_imag;
        _zz_256 = img_reg_array_31_5_real;
        _zz_257 = img_reg_array_31_5_imag;
        _zz_258 = img_reg_array_32_5_real;
        _zz_259 = img_reg_array_32_5_imag;
        _zz_260 = img_reg_array_33_5_real;
        _zz_261 = img_reg_array_33_5_imag;
        _zz_262 = img_reg_array_34_5_real;
        _zz_263 = img_reg_array_34_5_imag;
        _zz_264 = img_reg_array_35_5_real;
        _zz_265 = img_reg_array_35_5_imag;
        _zz_266 = img_reg_array_36_5_real;
        _zz_267 = img_reg_array_36_5_imag;
        _zz_268 = img_reg_array_37_5_real;
        _zz_269 = img_reg_array_37_5_imag;
        _zz_270 = img_reg_array_38_5_real;
        _zz_271 = img_reg_array_38_5_imag;
        _zz_272 = img_reg_array_39_5_real;
        _zz_273 = img_reg_array_39_5_imag;
        _zz_274 = img_reg_array_40_5_real;
        _zz_275 = img_reg_array_40_5_imag;
        _zz_276 = img_reg_array_41_5_real;
        _zz_277 = img_reg_array_41_5_imag;
        _zz_278 = img_reg_array_42_5_real;
        _zz_279 = img_reg_array_42_5_imag;
        _zz_280 = img_reg_array_43_5_real;
        _zz_281 = img_reg_array_43_5_imag;
        _zz_282 = img_reg_array_44_5_real;
        _zz_283 = img_reg_array_44_5_imag;
        _zz_284 = img_reg_array_45_5_real;
        _zz_285 = img_reg_array_45_5_imag;
        _zz_286 = img_reg_array_46_5_real;
        _zz_287 = img_reg_array_46_5_imag;
        _zz_288 = img_reg_array_47_5_real;
        _zz_289 = img_reg_array_47_5_imag;
        _zz_290 = img_reg_array_48_5_real;
        _zz_291 = img_reg_array_48_5_imag;
        _zz_292 = img_reg_array_49_5_real;
        _zz_293 = img_reg_array_49_5_imag;
        _zz_294 = img_reg_array_50_5_real;
        _zz_295 = img_reg_array_50_5_imag;
        _zz_296 = img_reg_array_51_5_real;
        _zz_297 = img_reg_array_51_5_imag;
        _zz_298 = img_reg_array_52_5_real;
        _zz_299 = img_reg_array_52_5_imag;
        _zz_300 = img_reg_array_53_5_real;
        _zz_301 = img_reg_array_53_5_imag;
        _zz_302 = img_reg_array_54_5_real;
        _zz_303 = img_reg_array_54_5_imag;
        _zz_304 = img_reg_array_55_5_real;
        _zz_305 = img_reg_array_55_5_imag;
        _zz_306 = img_reg_array_56_5_real;
        _zz_307 = img_reg_array_56_5_imag;
        _zz_308 = img_reg_array_57_5_real;
        _zz_309 = img_reg_array_57_5_imag;
        _zz_310 = img_reg_array_58_5_real;
        _zz_311 = img_reg_array_58_5_imag;
        _zz_312 = img_reg_array_59_5_real;
        _zz_313 = img_reg_array_59_5_imag;
        _zz_314 = img_reg_array_60_5_real;
        _zz_315 = img_reg_array_60_5_imag;
        _zz_316 = img_reg_array_61_5_real;
        _zz_317 = img_reg_array_61_5_imag;
        _zz_318 = img_reg_array_62_5_real;
        _zz_319 = img_reg_array_62_5_imag;
        _zz_320 = img_reg_array_63_5_real;
        _zz_321 = img_reg_array_63_5_imag;
      end
      6'b000110 : begin
        _zz_194 = img_reg_array_0_6_real;
        _zz_195 = img_reg_array_0_6_imag;
        _zz_196 = img_reg_array_1_6_real;
        _zz_197 = img_reg_array_1_6_imag;
        _zz_198 = img_reg_array_2_6_real;
        _zz_199 = img_reg_array_2_6_imag;
        _zz_200 = img_reg_array_3_6_real;
        _zz_201 = img_reg_array_3_6_imag;
        _zz_202 = img_reg_array_4_6_real;
        _zz_203 = img_reg_array_4_6_imag;
        _zz_204 = img_reg_array_5_6_real;
        _zz_205 = img_reg_array_5_6_imag;
        _zz_206 = img_reg_array_6_6_real;
        _zz_207 = img_reg_array_6_6_imag;
        _zz_208 = img_reg_array_7_6_real;
        _zz_209 = img_reg_array_7_6_imag;
        _zz_210 = img_reg_array_8_6_real;
        _zz_211 = img_reg_array_8_6_imag;
        _zz_212 = img_reg_array_9_6_real;
        _zz_213 = img_reg_array_9_6_imag;
        _zz_214 = img_reg_array_10_6_real;
        _zz_215 = img_reg_array_10_6_imag;
        _zz_216 = img_reg_array_11_6_real;
        _zz_217 = img_reg_array_11_6_imag;
        _zz_218 = img_reg_array_12_6_real;
        _zz_219 = img_reg_array_12_6_imag;
        _zz_220 = img_reg_array_13_6_real;
        _zz_221 = img_reg_array_13_6_imag;
        _zz_222 = img_reg_array_14_6_real;
        _zz_223 = img_reg_array_14_6_imag;
        _zz_224 = img_reg_array_15_6_real;
        _zz_225 = img_reg_array_15_6_imag;
        _zz_226 = img_reg_array_16_6_real;
        _zz_227 = img_reg_array_16_6_imag;
        _zz_228 = img_reg_array_17_6_real;
        _zz_229 = img_reg_array_17_6_imag;
        _zz_230 = img_reg_array_18_6_real;
        _zz_231 = img_reg_array_18_6_imag;
        _zz_232 = img_reg_array_19_6_real;
        _zz_233 = img_reg_array_19_6_imag;
        _zz_234 = img_reg_array_20_6_real;
        _zz_235 = img_reg_array_20_6_imag;
        _zz_236 = img_reg_array_21_6_real;
        _zz_237 = img_reg_array_21_6_imag;
        _zz_238 = img_reg_array_22_6_real;
        _zz_239 = img_reg_array_22_6_imag;
        _zz_240 = img_reg_array_23_6_real;
        _zz_241 = img_reg_array_23_6_imag;
        _zz_242 = img_reg_array_24_6_real;
        _zz_243 = img_reg_array_24_6_imag;
        _zz_244 = img_reg_array_25_6_real;
        _zz_245 = img_reg_array_25_6_imag;
        _zz_246 = img_reg_array_26_6_real;
        _zz_247 = img_reg_array_26_6_imag;
        _zz_248 = img_reg_array_27_6_real;
        _zz_249 = img_reg_array_27_6_imag;
        _zz_250 = img_reg_array_28_6_real;
        _zz_251 = img_reg_array_28_6_imag;
        _zz_252 = img_reg_array_29_6_real;
        _zz_253 = img_reg_array_29_6_imag;
        _zz_254 = img_reg_array_30_6_real;
        _zz_255 = img_reg_array_30_6_imag;
        _zz_256 = img_reg_array_31_6_real;
        _zz_257 = img_reg_array_31_6_imag;
        _zz_258 = img_reg_array_32_6_real;
        _zz_259 = img_reg_array_32_6_imag;
        _zz_260 = img_reg_array_33_6_real;
        _zz_261 = img_reg_array_33_6_imag;
        _zz_262 = img_reg_array_34_6_real;
        _zz_263 = img_reg_array_34_6_imag;
        _zz_264 = img_reg_array_35_6_real;
        _zz_265 = img_reg_array_35_6_imag;
        _zz_266 = img_reg_array_36_6_real;
        _zz_267 = img_reg_array_36_6_imag;
        _zz_268 = img_reg_array_37_6_real;
        _zz_269 = img_reg_array_37_6_imag;
        _zz_270 = img_reg_array_38_6_real;
        _zz_271 = img_reg_array_38_6_imag;
        _zz_272 = img_reg_array_39_6_real;
        _zz_273 = img_reg_array_39_6_imag;
        _zz_274 = img_reg_array_40_6_real;
        _zz_275 = img_reg_array_40_6_imag;
        _zz_276 = img_reg_array_41_6_real;
        _zz_277 = img_reg_array_41_6_imag;
        _zz_278 = img_reg_array_42_6_real;
        _zz_279 = img_reg_array_42_6_imag;
        _zz_280 = img_reg_array_43_6_real;
        _zz_281 = img_reg_array_43_6_imag;
        _zz_282 = img_reg_array_44_6_real;
        _zz_283 = img_reg_array_44_6_imag;
        _zz_284 = img_reg_array_45_6_real;
        _zz_285 = img_reg_array_45_6_imag;
        _zz_286 = img_reg_array_46_6_real;
        _zz_287 = img_reg_array_46_6_imag;
        _zz_288 = img_reg_array_47_6_real;
        _zz_289 = img_reg_array_47_6_imag;
        _zz_290 = img_reg_array_48_6_real;
        _zz_291 = img_reg_array_48_6_imag;
        _zz_292 = img_reg_array_49_6_real;
        _zz_293 = img_reg_array_49_6_imag;
        _zz_294 = img_reg_array_50_6_real;
        _zz_295 = img_reg_array_50_6_imag;
        _zz_296 = img_reg_array_51_6_real;
        _zz_297 = img_reg_array_51_6_imag;
        _zz_298 = img_reg_array_52_6_real;
        _zz_299 = img_reg_array_52_6_imag;
        _zz_300 = img_reg_array_53_6_real;
        _zz_301 = img_reg_array_53_6_imag;
        _zz_302 = img_reg_array_54_6_real;
        _zz_303 = img_reg_array_54_6_imag;
        _zz_304 = img_reg_array_55_6_real;
        _zz_305 = img_reg_array_55_6_imag;
        _zz_306 = img_reg_array_56_6_real;
        _zz_307 = img_reg_array_56_6_imag;
        _zz_308 = img_reg_array_57_6_real;
        _zz_309 = img_reg_array_57_6_imag;
        _zz_310 = img_reg_array_58_6_real;
        _zz_311 = img_reg_array_58_6_imag;
        _zz_312 = img_reg_array_59_6_real;
        _zz_313 = img_reg_array_59_6_imag;
        _zz_314 = img_reg_array_60_6_real;
        _zz_315 = img_reg_array_60_6_imag;
        _zz_316 = img_reg_array_61_6_real;
        _zz_317 = img_reg_array_61_6_imag;
        _zz_318 = img_reg_array_62_6_real;
        _zz_319 = img_reg_array_62_6_imag;
        _zz_320 = img_reg_array_63_6_real;
        _zz_321 = img_reg_array_63_6_imag;
      end
      6'b000111 : begin
        _zz_194 = img_reg_array_0_7_real;
        _zz_195 = img_reg_array_0_7_imag;
        _zz_196 = img_reg_array_1_7_real;
        _zz_197 = img_reg_array_1_7_imag;
        _zz_198 = img_reg_array_2_7_real;
        _zz_199 = img_reg_array_2_7_imag;
        _zz_200 = img_reg_array_3_7_real;
        _zz_201 = img_reg_array_3_7_imag;
        _zz_202 = img_reg_array_4_7_real;
        _zz_203 = img_reg_array_4_7_imag;
        _zz_204 = img_reg_array_5_7_real;
        _zz_205 = img_reg_array_5_7_imag;
        _zz_206 = img_reg_array_6_7_real;
        _zz_207 = img_reg_array_6_7_imag;
        _zz_208 = img_reg_array_7_7_real;
        _zz_209 = img_reg_array_7_7_imag;
        _zz_210 = img_reg_array_8_7_real;
        _zz_211 = img_reg_array_8_7_imag;
        _zz_212 = img_reg_array_9_7_real;
        _zz_213 = img_reg_array_9_7_imag;
        _zz_214 = img_reg_array_10_7_real;
        _zz_215 = img_reg_array_10_7_imag;
        _zz_216 = img_reg_array_11_7_real;
        _zz_217 = img_reg_array_11_7_imag;
        _zz_218 = img_reg_array_12_7_real;
        _zz_219 = img_reg_array_12_7_imag;
        _zz_220 = img_reg_array_13_7_real;
        _zz_221 = img_reg_array_13_7_imag;
        _zz_222 = img_reg_array_14_7_real;
        _zz_223 = img_reg_array_14_7_imag;
        _zz_224 = img_reg_array_15_7_real;
        _zz_225 = img_reg_array_15_7_imag;
        _zz_226 = img_reg_array_16_7_real;
        _zz_227 = img_reg_array_16_7_imag;
        _zz_228 = img_reg_array_17_7_real;
        _zz_229 = img_reg_array_17_7_imag;
        _zz_230 = img_reg_array_18_7_real;
        _zz_231 = img_reg_array_18_7_imag;
        _zz_232 = img_reg_array_19_7_real;
        _zz_233 = img_reg_array_19_7_imag;
        _zz_234 = img_reg_array_20_7_real;
        _zz_235 = img_reg_array_20_7_imag;
        _zz_236 = img_reg_array_21_7_real;
        _zz_237 = img_reg_array_21_7_imag;
        _zz_238 = img_reg_array_22_7_real;
        _zz_239 = img_reg_array_22_7_imag;
        _zz_240 = img_reg_array_23_7_real;
        _zz_241 = img_reg_array_23_7_imag;
        _zz_242 = img_reg_array_24_7_real;
        _zz_243 = img_reg_array_24_7_imag;
        _zz_244 = img_reg_array_25_7_real;
        _zz_245 = img_reg_array_25_7_imag;
        _zz_246 = img_reg_array_26_7_real;
        _zz_247 = img_reg_array_26_7_imag;
        _zz_248 = img_reg_array_27_7_real;
        _zz_249 = img_reg_array_27_7_imag;
        _zz_250 = img_reg_array_28_7_real;
        _zz_251 = img_reg_array_28_7_imag;
        _zz_252 = img_reg_array_29_7_real;
        _zz_253 = img_reg_array_29_7_imag;
        _zz_254 = img_reg_array_30_7_real;
        _zz_255 = img_reg_array_30_7_imag;
        _zz_256 = img_reg_array_31_7_real;
        _zz_257 = img_reg_array_31_7_imag;
        _zz_258 = img_reg_array_32_7_real;
        _zz_259 = img_reg_array_32_7_imag;
        _zz_260 = img_reg_array_33_7_real;
        _zz_261 = img_reg_array_33_7_imag;
        _zz_262 = img_reg_array_34_7_real;
        _zz_263 = img_reg_array_34_7_imag;
        _zz_264 = img_reg_array_35_7_real;
        _zz_265 = img_reg_array_35_7_imag;
        _zz_266 = img_reg_array_36_7_real;
        _zz_267 = img_reg_array_36_7_imag;
        _zz_268 = img_reg_array_37_7_real;
        _zz_269 = img_reg_array_37_7_imag;
        _zz_270 = img_reg_array_38_7_real;
        _zz_271 = img_reg_array_38_7_imag;
        _zz_272 = img_reg_array_39_7_real;
        _zz_273 = img_reg_array_39_7_imag;
        _zz_274 = img_reg_array_40_7_real;
        _zz_275 = img_reg_array_40_7_imag;
        _zz_276 = img_reg_array_41_7_real;
        _zz_277 = img_reg_array_41_7_imag;
        _zz_278 = img_reg_array_42_7_real;
        _zz_279 = img_reg_array_42_7_imag;
        _zz_280 = img_reg_array_43_7_real;
        _zz_281 = img_reg_array_43_7_imag;
        _zz_282 = img_reg_array_44_7_real;
        _zz_283 = img_reg_array_44_7_imag;
        _zz_284 = img_reg_array_45_7_real;
        _zz_285 = img_reg_array_45_7_imag;
        _zz_286 = img_reg_array_46_7_real;
        _zz_287 = img_reg_array_46_7_imag;
        _zz_288 = img_reg_array_47_7_real;
        _zz_289 = img_reg_array_47_7_imag;
        _zz_290 = img_reg_array_48_7_real;
        _zz_291 = img_reg_array_48_7_imag;
        _zz_292 = img_reg_array_49_7_real;
        _zz_293 = img_reg_array_49_7_imag;
        _zz_294 = img_reg_array_50_7_real;
        _zz_295 = img_reg_array_50_7_imag;
        _zz_296 = img_reg_array_51_7_real;
        _zz_297 = img_reg_array_51_7_imag;
        _zz_298 = img_reg_array_52_7_real;
        _zz_299 = img_reg_array_52_7_imag;
        _zz_300 = img_reg_array_53_7_real;
        _zz_301 = img_reg_array_53_7_imag;
        _zz_302 = img_reg_array_54_7_real;
        _zz_303 = img_reg_array_54_7_imag;
        _zz_304 = img_reg_array_55_7_real;
        _zz_305 = img_reg_array_55_7_imag;
        _zz_306 = img_reg_array_56_7_real;
        _zz_307 = img_reg_array_56_7_imag;
        _zz_308 = img_reg_array_57_7_real;
        _zz_309 = img_reg_array_57_7_imag;
        _zz_310 = img_reg_array_58_7_real;
        _zz_311 = img_reg_array_58_7_imag;
        _zz_312 = img_reg_array_59_7_real;
        _zz_313 = img_reg_array_59_7_imag;
        _zz_314 = img_reg_array_60_7_real;
        _zz_315 = img_reg_array_60_7_imag;
        _zz_316 = img_reg_array_61_7_real;
        _zz_317 = img_reg_array_61_7_imag;
        _zz_318 = img_reg_array_62_7_real;
        _zz_319 = img_reg_array_62_7_imag;
        _zz_320 = img_reg_array_63_7_real;
        _zz_321 = img_reg_array_63_7_imag;
      end
      6'b001000 : begin
        _zz_194 = img_reg_array_0_8_real;
        _zz_195 = img_reg_array_0_8_imag;
        _zz_196 = img_reg_array_1_8_real;
        _zz_197 = img_reg_array_1_8_imag;
        _zz_198 = img_reg_array_2_8_real;
        _zz_199 = img_reg_array_2_8_imag;
        _zz_200 = img_reg_array_3_8_real;
        _zz_201 = img_reg_array_3_8_imag;
        _zz_202 = img_reg_array_4_8_real;
        _zz_203 = img_reg_array_4_8_imag;
        _zz_204 = img_reg_array_5_8_real;
        _zz_205 = img_reg_array_5_8_imag;
        _zz_206 = img_reg_array_6_8_real;
        _zz_207 = img_reg_array_6_8_imag;
        _zz_208 = img_reg_array_7_8_real;
        _zz_209 = img_reg_array_7_8_imag;
        _zz_210 = img_reg_array_8_8_real;
        _zz_211 = img_reg_array_8_8_imag;
        _zz_212 = img_reg_array_9_8_real;
        _zz_213 = img_reg_array_9_8_imag;
        _zz_214 = img_reg_array_10_8_real;
        _zz_215 = img_reg_array_10_8_imag;
        _zz_216 = img_reg_array_11_8_real;
        _zz_217 = img_reg_array_11_8_imag;
        _zz_218 = img_reg_array_12_8_real;
        _zz_219 = img_reg_array_12_8_imag;
        _zz_220 = img_reg_array_13_8_real;
        _zz_221 = img_reg_array_13_8_imag;
        _zz_222 = img_reg_array_14_8_real;
        _zz_223 = img_reg_array_14_8_imag;
        _zz_224 = img_reg_array_15_8_real;
        _zz_225 = img_reg_array_15_8_imag;
        _zz_226 = img_reg_array_16_8_real;
        _zz_227 = img_reg_array_16_8_imag;
        _zz_228 = img_reg_array_17_8_real;
        _zz_229 = img_reg_array_17_8_imag;
        _zz_230 = img_reg_array_18_8_real;
        _zz_231 = img_reg_array_18_8_imag;
        _zz_232 = img_reg_array_19_8_real;
        _zz_233 = img_reg_array_19_8_imag;
        _zz_234 = img_reg_array_20_8_real;
        _zz_235 = img_reg_array_20_8_imag;
        _zz_236 = img_reg_array_21_8_real;
        _zz_237 = img_reg_array_21_8_imag;
        _zz_238 = img_reg_array_22_8_real;
        _zz_239 = img_reg_array_22_8_imag;
        _zz_240 = img_reg_array_23_8_real;
        _zz_241 = img_reg_array_23_8_imag;
        _zz_242 = img_reg_array_24_8_real;
        _zz_243 = img_reg_array_24_8_imag;
        _zz_244 = img_reg_array_25_8_real;
        _zz_245 = img_reg_array_25_8_imag;
        _zz_246 = img_reg_array_26_8_real;
        _zz_247 = img_reg_array_26_8_imag;
        _zz_248 = img_reg_array_27_8_real;
        _zz_249 = img_reg_array_27_8_imag;
        _zz_250 = img_reg_array_28_8_real;
        _zz_251 = img_reg_array_28_8_imag;
        _zz_252 = img_reg_array_29_8_real;
        _zz_253 = img_reg_array_29_8_imag;
        _zz_254 = img_reg_array_30_8_real;
        _zz_255 = img_reg_array_30_8_imag;
        _zz_256 = img_reg_array_31_8_real;
        _zz_257 = img_reg_array_31_8_imag;
        _zz_258 = img_reg_array_32_8_real;
        _zz_259 = img_reg_array_32_8_imag;
        _zz_260 = img_reg_array_33_8_real;
        _zz_261 = img_reg_array_33_8_imag;
        _zz_262 = img_reg_array_34_8_real;
        _zz_263 = img_reg_array_34_8_imag;
        _zz_264 = img_reg_array_35_8_real;
        _zz_265 = img_reg_array_35_8_imag;
        _zz_266 = img_reg_array_36_8_real;
        _zz_267 = img_reg_array_36_8_imag;
        _zz_268 = img_reg_array_37_8_real;
        _zz_269 = img_reg_array_37_8_imag;
        _zz_270 = img_reg_array_38_8_real;
        _zz_271 = img_reg_array_38_8_imag;
        _zz_272 = img_reg_array_39_8_real;
        _zz_273 = img_reg_array_39_8_imag;
        _zz_274 = img_reg_array_40_8_real;
        _zz_275 = img_reg_array_40_8_imag;
        _zz_276 = img_reg_array_41_8_real;
        _zz_277 = img_reg_array_41_8_imag;
        _zz_278 = img_reg_array_42_8_real;
        _zz_279 = img_reg_array_42_8_imag;
        _zz_280 = img_reg_array_43_8_real;
        _zz_281 = img_reg_array_43_8_imag;
        _zz_282 = img_reg_array_44_8_real;
        _zz_283 = img_reg_array_44_8_imag;
        _zz_284 = img_reg_array_45_8_real;
        _zz_285 = img_reg_array_45_8_imag;
        _zz_286 = img_reg_array_46_8_real;
        _zz_287 = img_reg_array_46_8_imag;
        _zz_288 = img_reg_array_47_8_real;
        _zz_289 = img_reg_array_47_8_imag;
        _zz_290 = img_reg_array_48_8_real;
        _zz_291 = img_reg_array_48_8_imag;
        _zz_292 = img_reg_array_49_8_real;
        _zz_293 = img_reg_array_49_8_imag;
        _zz_294 = img_reg_array_50_8_real;
        _zz_295 = img_reg_array_50_8_imag;
        _zz_296 = img_reg_array_51_8_real;
        _zz_297 = img_reg_array_51_8_imag;
        _zz_298 = img_reg_array_52_8_real;
        _zz_299 = img_reg_array_52_8_imag;
        _zz_300 = img_reg_array_53_8_real;
        _zz_301 = img_reg_array_53_8_imag;
        _zz_302 = img_reg_array_54_8_real;
        _zz_303 = img_reg_array_54_8_imag;
        _zz_304 = img_reg_array_55_8_real;
        _zz_305 = img_reg_array_55_8_imag;
        _zz_306 = img_reg_array_56_8_real;
        _zz_307 = img_reg_array_56_8_imag;
        _zz_308 = img_reg_array_57_8_real;
        _zz_309 = img_reg_array_57_8_imag;
        _zz_310 = img_reg_array_58_8_real;
        _zz_311 = img_reg_array_58_8_imag;
        _zz_312 = img_reg_array_59_8_real;
        _zz_313 = img_reg_array_59_8_imag;
        _zz_314 = img_reg_array_60_8_real;
        _zz_315 = img_reg_array_60_8_imag;
        _zz_316 = img_reg_array_61_8_real;
        _zz_317 = img_reg_array_61_8_imag;
        _zz_318 = img_reg_array_62_8_real;
        _zz_319 = img_reg_array_62_8_imag;
        _zz_320 = img_reg_array_63_8_real;
        _zz_321 = img_reg_array_63_8_imag;
      end
      6'b001001 : begin
        _zz_194 = img_reg_array_0_9_real;
        _zz_195 = img_reg_array_0_9_imag;
        _zz_196 = img_reg_array_1_9_real;
        _zz_197 = img_reg_array_1_9_imag;
        _zz_198 = img_reg_array_2_9_real;
        _zz_199 = img_reg_array_2_9_imag;
        _zz_200 = img_reg_array_3_9_real;
        _zz_201 = img_reg_array_3_9_imag;
        _zz_202 = img_reg_array_4_9_real;
        _zz_203 = img_reg_array_4_9_imag;
        _zz_204 = img_reg_array_5_9_real;
        _zz_205 = img_reg_array_5_9_imag;
        _zz_206 = img_reg_array_6_9_real;
        _zz_207 = img_reg_array_6_9_imag;
        _zz_208 = img_reg_array_7_9_real;
        _zz_209 = img_reg_array_7_9_imag;
        _zz_210 = img_reg_array_8_9_real;
        _zz_211 = img_reg_array_8_9_imag;
        _zz_212 = img_reg_array_9_9_real;
        _zz_213 = img_reg_array_9_9_imag;
        _zz_214 = img_reg_array_10_9_real;
        _zz_215 = img_reg_array_10_9_imag;
        _zz_216 = img_reg_array_11_9_real;
        _zz_217 = img_reg_array_11_9_imag;
        _zz_218 = img_reg_array_12_9_real;
        _zz_219 = img_reg_array_12_9_imag;
        _zz_220 = img_reg_array_13_9_real;
        _zz_221 = img_reg_array_13_9_imag;
        _zz_222 = img_reg_array_14_9_real;
        _zz_223 = img_reg_array_14_9_imag;
        _zz_224 = img_reg_array_15_9_real;
        _zz_225 = img_reg_array_15_9_imag;
        _zz_226 = img_reg_array_16_9_real;
        _zz_227 = img_reg_array_16_9_imag;
        _zz_228 = img_reg_array_17_9_real;
        _zz_229 = img_reg_array_17_9_imag;
        _zz_230 = img_reg_array_18_9_real;
        _zz_231 = img_reg_array_18_9_imag;
        _zz_232 = img_reg_array_19_9_real;
        _zz_233 = img_reg_array_19_9_imag;
        _zz_234 = img_reg_array_20_9_real;
        _zz_235 = img_reg_array_20_9_imag;
        _zz_236 = img_reg_array_21_9_real;
        _zz_237 = img_reg_array_21_9_imag;
        _zz_238 = img_reg_array_22_9_real;
        _zz_239 = img_reg_array_22_9_imag;
        _zz_240 = img_reg_array_23_9_real;
        _zz_241 = img_reg_array_23_9_imag;
        _zz_242 = img_reg_array_24_9_real;
        _zz_243 = img_reg_array_24_9_imag;
        _zz_244 = img_reg_array_25_9_real;
        _zz_245 = img_reg_array_25_9_imag;
        _zz_246 = img_reg_array_26_9_real;
        _zz_247 = img_reg_array_26_9_imag;
        _zz_248 = img_reg_array_27_9_real;
        _zz_249 = img_reg_array_27_9_imag;
        _zz_250 = img_reg_array_28_9_real;
        _zz_251 = img_reg_array_28_9_imag;
        _zz_252 = img_reg_array_29_9_real;
        _zz_253 = img_reg_array_29_9_imag;
        _zz_254 = img_reg_array_30_9_real;
        _zz_255 = img_reg_array_30_9_imag;
        _zz_256 = img_reg_array_31_9_real;
        _zz_257 = img_reg_array_31_9_imag;
        _zz_258 = img_reg_array_32_9_real;
        _zz_259 = img_reg_array_32_9_imag;
        _zz_260 = img_reg_array_33_9_real;
        _zz_261 = img_reg_array_33_9_imag;
        _zz_262 = img_reg_array_34_9_real;
        _zz_263 = img_reg_array_34_9_imag;
        _zz_264 = img_reg_array_35_9_real;
        _zz_265 = img_reg_array_35_9_imag;
        _zz_266 = img_reg_array_36_9_real;
        _zz_267 = img_reg_array_36_9_imag;
        _zz_268 = img_reg_array_37_9_real;
        _zz_269 = img_reg_array_37_9_imag;
        _zz_270 = img_reg_array_38_9_real;
        _zz_271 = img_reg_array_38_9_imag;
        _zz_272 = img_reg_array_39_9_real;
        _zz_273 = img_reg_array_39_9_imag;
        _zz_274 = img_reg_array_40_9_real;
        _zz_275 = img_reg_array_40_9_imag;
        _zz_276 = img_reg_array_41_9_real;
        _zz_277 = img_reg_array_41_9_imag;
        _zz_278 = img_reg_array_42_9_real;
        _zz_279 = img_reg_array_42_9_imag;
        _zz_280 = img_reg_array_43_9_real;
        _zz_281 = img_reg_array_43_9_imag;
        _zz_282 = img_reg_array_44_9_real;
        _zz_283 = img_reg_array_44_9_imag;
        _zz_284 = img_reg_array_45_9_real;
        _zz_285 = img_reg_array_45_9_imag;
        _zz_286 = img_reg_array_46_9_real;
        _zz_287 = img_reg_array_46_9_imag;
        _zz_288 = img_reg_array_47_9_real;
        _zz_289 = img_reg_array_47_9_imag;
        _zz_290 = img_reg_array_48_9_real;
        _zz_291 = img_reg_array_48_9_imag;
        _zz_292 = img_reg_array_49_9_real;
        _zz_293 = img_reg_array_49_9_imag;
        _zz_294 = img_reg_array_50_9_real;
        _zz_295 = img_reg_array_50_9_imag;
        _zz_296 = img_reg_array_51_9_real;
        _zz_297 = img_reg_array_51_9_imag;
        _zz_298 = img_reg_array_52_9_real;
        _zz_299 = img_reg_array_52_9_imag;
        _zz_300 = img_reg_array_53_9_real;
        _zz_301 = img_reg_array_53_9_imag;
        _zz_302 = img_reg_array_54_9_real;
        _zz_303 = img_reg_array_54_9_imag;
        _zz_304 = img_reg_array_55_9_real;
        _zz_305 = img_reg_array_55_9_imag;
        _zz_306 = img_reg_array_56_9_real;
        _zz_307 = img_reg_array_56_9_imag;
        _zz_308 = img_reg_array_57_9_real;
        _zz_309 = img_reg_array_57_9_imag;
        _zz_310 = img_reg_array_58_9_real;
        _zz_311 = img_reg_array_58_9_imag;
        _zz_312 = img_reg_array_59_9_real;
        _zz_313 = img_reg_array_59_9_imag;
        _zz_314 = img_reg_array_60_9_real;
        _zz_315 = img_reg_array_60_9_imag;
        _zz_316 = img_reg_array_61_9_real;
        _zz_317 = img_reg_array_61_9_imag;
        _zz_318 = img_reg_array_62_9_real;
        _zz_319 = img_reg_array_62_9_imag;
        _zz_320 = img_reg_array_63_9_real;
        _zz_321 = img_reg_array_63_9_imag;
      end
      6'b001010 : begin
        _zz_194 = img_reg_array_0_10_real;
        _zz_195 = img_reg_array_0_10_imag;
        _zz_196 = img_reg_array_1_10_real;
        _zz_197 = img_reg_array_1_10_imag;
        _zz_198 = img_reg_array_2_10_real;
        _zz_199 = img_reg_array_2_10_imag;
        _zz_200 = img_reg_array_3_10_real;
        _zz_201 = img_reg_array_3_10_imag;
        _zz_202 = img_reg_array_4_10_real;
        _zz_203 = img_reg_array_4_10_imag;
        _zz_204 = img_reg_array_5_10_real;
        _zz_205 = img_reg_array_5_10_imag;
        _zz_206 = img_reg_array_6_10_real;
        _zz_207 = img_reg_array_6_10_imag;
        _zz_208 = img_reg_array_7_10_real;
        _zz_209 = img_reg_array_7_10_imag;
        _zz_210 = img_reg_array_8_10_real;
        _zz_211 = img_reg_array_8_10_imag;
        _zz_212 = img_reg_array_9_10_real;
        _zz_213 = img_reg_array_9_10_imag;
        _zz_214 = img_reg_array_10_10_real;
        _zz_215 = img_reg_array_10_10_imag;
        _zz_216 = img_reg_array_11_10_real;
        _zz_217 = img_reg_array_11_10_imag;
        _zz_218 = img_reg_array_12_10_real;
        _zz_219 = img_reg_array_12_10_imag;
        _zz_220 = img_reg_array_13_10_real;
        _zz_221 = img_reg_array_13_10_imag;
        _zz_222 = img_reg_array_14_10_real;
        _zz_223 = img_reg_array_14_10_imag;
        _zz_224 = img_reg_array_15_10_real;
        _zz_225 = img_reg_array_15_10_imag;
        _zz_226 = img_reg_array_16_10_real;
        _zz_227 = img_reg_array_16_10_imag;
        _zz_228 = img_reg_array_17_10_real;
        _zz_229 = img_reg_array_17_10_imag;
        _zz_230 = img_reg_array_18_10_real;
        _zz_231 = img_reg_array_18_10_imag;
        _zz_232 = img_reg_array_19_10_real;
        _zz_233 = img_reg_array_19_10_imag;
        _zz_234 = img_reg_array_20_10_real;
        _zz_235 = img_reg_array_20_10_imag;
        _zz_236 = img_reg_array_21_10_real;
        _zz_237 = img_reg_array_21_10_imag;
        _zz_238 = img_reg_array_22_10_real;
        _zz_239 = img_reg_array_22_10_imag;
        _zz_240 = img_reg_array_23_10_real;
        _zz_241 = img_reg_array_23_10_imag;
        _zz_242 = img_reg_array_24_10_real;
        _zz_243 = img_reg_array_24_10_imag;
        _zz_244 = img_reg_array_25_10_real;
        _zz_245 = img_reg_array_25_10_imag;
        _zz_246 = img_reg_array_26_10_real;
        _zz_247 = img_reg_array_26_10_imag;
        _zz_248 = img_reg_array_27_10_real;
        _zz_249 = img_reg_array_27_10_imag;
        _zz_250 = img_reg_array_28_10_real;
        _zz_251 = img_reg_array_28_10_imag;
        _zz_252 = img_reg_array_29_10_real;
        _zz_253 = img_reg_array_29_10_imag;
        _zz_254 = img_reg_array_30_10_real;
        _zz_255 = img_reg_array_30_10_imag;
        _zz_256 = img_reg_array_31_10_real;
        _zz_257 = img_reg_array_31_10_imag;
        _zz_258 = img_reg_array_32_10_real;
        _zz_259 = img_reg_array_32_10_imag;
        _zz_260 = img_reg_array_33_10_real;
        _zz_261 = img_reg_array_33_10_imag;
        _zz_262 = img_reg_array_34_10_real;
        _zz_263 = img_reg_array_34_10_imag;
        _zz_264 = img_reg_array_35_10_real;
        _zz_265 = img_reg_array_35_10_imag;
        _zz_266 = img_reg_array_36_10_real;
        _zz_267 = img_reg_array_36_10_imag;
        _zz_268 = img_reg_array_37_10_real;
        _zz_269 = img_reg_array_37_10_imag;
        _zz_270 = img_reg_array_38_10_real;
        _zz_271 = img_reg_array_38_10_imag;
        _zz_272 = img_reg_array_39_10_real;
        _zz_273 = img_reg_array_39_10_imag;
        _zz_274 = img_reg_array_40_10_real;
        _zz_275 = img_reg_array_40_10_imag;
        _zz_276 = img_reg_array_41_10_real;
        _zz_277 = img_reg_array_41_10_imag;
        _zz_278 = img_reg_array_42_10_real;
        _zz_279 = img_reg_array_42_10_imag;
        _zz_280 = img_reg_array_43_10_real;
        _zz_281 = img_reg_array_43_10_imag;
        _zz_282 = img_reg_array_44_10_real;
        _zz_283 = img_reg_array_44_10_imag;
        _zz_284 = img_reg_array_45_10_real;
        _zz_285 = img_reg_array_45_10_imag;
        _zz_286 = img_reg_array_46_10_real;
        _zz_287 = img_reg_array_46_10_imag;
        _zz_288 = img_reg_array_47_10_real;
        _zz_289 = img_reg_array_47_10_imag;
        _zz_290 = img_reg_array_48_10_real;
        _zz_291 = img_reg_array_48_10_imag;
        _zz_292 = img_reg_array_49_10_real;
        _zz_293 = img_reg_array_49_10_imag;
        _zz_294 = img_reg_array_50_10_real;
        _zz_295 = img_reg_array_50_10_imag;
        _zz_296 = img_reg_array_51_10_real;
        _zz_297 = img_reg_array_51_10_imag;
        _zz_298 = img_reg_array_52_10_real;
        _zz_299 = img_reg_array_52_10_imag;
        _zz_300 = img_reg_array_53_10_real;
        _zz_301 = img_reg_array_53_10_imag;
        _zz_302 = img_reg_array_54_10_real;
        _zz_303 = img_reg_array_54_10_imag;
        _zz_304 = img_reg_array_55_10_real;
        _zz_305 = img_reg_array_55_10_imag;
        _zz_306 = img_reg_array_56_10_real;
        _zz_307 = img_reg_array_56_10_imag;
        _zz_308 = img_reg_array_57_10_real;
        _zz_309 = img_reg_array_57_10_imag;
        _zz_310 = img_reg_array_58_10_real;
        _zz_311 = img_reg_array_58_10_imag;
        _zz_312 = img_reg_array_59_10_real;
        _zz_313 = img_reg_array_59_10_imag;
        _zz_314 = img_reg_array_60_10_real;
        _zz_315 = img_reg_array_60_10_imag;
        _zz_316 = img_reg_array_61_10_real;
        _zz_317 = img_reg_array_61_10_imag;
        _zz_318 = img_reg_array_62_10_real;
        _zz_319 = img_reg_array_62_10_imag;
        _zz_320 = img_reg_array_63_10_real;
        _zz_321 = img_reg_array_63_10_imag;
      end
      6'b001011 : begin
        _zz_194 = img_reg_array_0_11_real;
        _zz_195 = img_reg_array_0_11_imag;
        _zz_196 = img_reg_array_1_11_real;
        _zz_197 = img_reg_array_1_11_imag;
        _zz_198 = img_reg_array_2_11_real;
        _zz_199 = img_reg_array_2_11_imag;
        _zz_200 = img_reg_array_3_11_real;
        _zz_201 = img_reg_array_3_11_imag;
        _zz_202 = img_reg_array_4_11_real;
        _zz_203 = img_reg_array_4_11_imag;
        _zz_204 = img_reg_array_5_11_real;
        _zz_205 = img_reg_array_5_11_imag;
        _zz_206 = img_reg_array_6_11_real;
        _zz_207 = img_reg_array_6_11_imag;
        _zz_208 = img_reg_array_7_11_real;
        _zz_209 = img_reg_array_7_11_imag;
        _zz_210 = img_reg_array_8_11_real;
        _zz_211 = img_reg_array_8_11_imag;
        _zz_212 = img_reg_array_9_11_real;
        _zz_213 = img_reg_array_9_11_imag;
        _zz_214 = img_reg_array_10_11_real;
        _zz_215 = img_reg_array_10_11_imag;
        _zz_216 = img_reg_array_11_11_real;
        _zz_217 = img_reg_array_11_11_imag;
        _zz_218 = img_reg_array_12_11_real;
        _zz_219 = img_reg_array_12_11_imag;
        _zz_220 = img_reg_array_13_11_real;
        _zz_221 = img_reg_array_13_11_imag;
        _zz_222 = img_reg_array_14_11_real;
        _zz_223 = img_reg_array_14_11_imag;
        _zz_224 = img_reg_array_15_11_real;
        _zz_225 = img_reg_array_15_11_imag;
        _zz_226 = img_reg_array_16_11_real;
        _zz_227 = img_reg_array_16_11_imag;
        _zz_228 = img_reg_array_17_11_real;
        _zz_229 = img_reg_array_17_11_imag;
        _zz_230 = img_reg_array_18_11_real;
        _zz_231 = img_reg_array_18_11_imag;
        _zz_232 = img_reg_array_19_11_real;
        _zz_233 = img_reg_array_19_11_imag;
        _zz_234 = img_reg_array_20_11_real;
        _zz_235 = img_reg_array_20_11_imag;
        _zz_236 = img_reg_array_21_11_real;
        _zz_237 = img_reg_array_21_11_imag;
        _zz_238 = img_reg_array_22_11_real;
        _zz_239 = img_reg_array_22_11_imag;
        _zz_240 = img_reg_array_23_11_real;
        _zz_241 = img_reg_array_23_11_imag;
        _zz_242 = img_reg_array_24_11_real;
        _zz_243 = img_reg_array_24_11_imag;
        _zz_244 = img_reg_array_25_11_real;
        _zz_245 = img_reg_array_25_11_imag;
        _zz_246 = img_reg_array_26_11_real;
        _zz_247 = img_reg_array_26_11_imag;
        _zz_248 = img_reg_array_27_11_real;
        _zz_249 = img_reg_array_27_11_imag;
        _zz_250 = img_reg_array_28_11_real;
        _zz_251 = img_reg_array_28_11_imag;
        _zz_252 = img_reg_array_29_11_real;
        _zz_253 = img_reg_array_29_11_imag;
        _zz_254 = img_reg_array_30_11_real;
        _zz_255 = img_reg_array_30_11_imag;
        _zz_256 = img_reg_array_31_11_real;
        _zz_257 = img_reg_array_31_11_imag;
        _zz_258 = img_reg_array_32_11_real;
        _zz_259 = img_reg_array_32_11_imag;
        _zz_260 = img_reg_array_33_11_real;
        _zz_261 = img_reg_array_33_11_imag;
        _zz_262 = img_reg_array_34_11_real;
        _zz_263 = img_reg_array_34_11_imag;
        _zz_264 = img_reg_array_35_11_real;
        _zz_265 = img_reg_array_35_11_imag;
        _zz_266 = img_reg_array_36_11_real;
        _zz_267 = img_reg_array_36_11_imag;
        _zz_268 = img_reg_array_37_11_real;
        _zz_269 = img_reg_array_37_11_imag;
        _zz_270 = img_reg_array_38_11_real;
        _zz_271 = img_reg_array_38_11_imag;
        _zz_272 = img_reg_array_39_11_real;
        _zz_273 = img_reg_array_39_11_imag;
        _zz_274 = img_reg_array_40_11_real;
        _zz_275 = img_reg_array_40_11_imag;
        _zz_276 = img_reg_array_41_11_real;
        _zz_277 = img_reg_array_41_11_imag;
        _zz_278 = img_reg_array_42_11_real;
        _zz_279 = img_reg_array_42_11_imag;
        _zz_280 = img_reg_array_43_11_real;
        _zz_281 = img_reg_array_43_11_imag;
        _zz_282 = img_reg_array_44_11_real;
        _zz_283 = img_reg_array_44_11_imag;
        _zz_284 = img_reg_array_45_11_real;
        _zz_285 = img_reg_array_45_11_imag;
        _zz_286 = img_reg_array_46_11_real;
        _zz_287 = img_reg_array_46_11_imag;
        _zz_288 = img_reg_array_47_11_real;
        _zz_289 = img_reg_array_47_11_imag;
        _zz_290 = img_reg_array_48_11_real;
        _zz_291 = img_reg_array_48_11_imag;
        _zz_292 = img_reg_array_49_11_real;
        _zz_293 = img_reg_array_49_11_imag;
        _zz_294 = img_reg_array_50_11_real;
        _zz_295 = img_reg_array_50_11_imag;
        _zz_296 = img_reg_array_51_11_real;
        _zz_297 = img_reg_array_51_11_imag;
        _zz_298 = img_reg_array_52_11_real;
        _zz_299 = img_reg_array_52_11_imag;
        _zz_300 = img_reg_array_53_11_real;
        _zz_301 = img_reg_array_53_11_imag;
        _zz_302 = img_reg_array_54_11_real;
        _zz_303 = img_reg_array_54_11_imag;
        _zz_304 = img_reg_array_55_11_real;
        _zz_305 = img_reg_array_55_11_imag;
        _zz_306 = img_reg_array_56_11_real;
        _zz_307 = img_reg_array_56_11_imag;
        _zz_308 = img_reg_array_57_11_real;
        _zz_309 = img_reg_array_57_11_imag;
        _zz_310 = img_reg_array_58_11_real;
        _zz_311 = img_reg_array_58_11_imag;
        _zz_312 = img_reg_array_59_11_real;
        _zz_313 = img_reg_array_59_11_imag;
        _zz_314 = img_reg_array_60_11_real;
        _zz_315 = img_reg_array_60_11_imag;
        _zz_316 = img_reg_array_61_11_real;
        _zz_317 = img_reg_array_61_11_imag;
        _zz_318 = img_reg_array_62_11_real;
        _zz_319 = img_reg_array_62_11_imag;
        _zz_320 = img_reg_array_63_11_real;
        _zz_321 = img_reg_array_63_11_imag;
      end
      6'b001100 : begin
        _zz_194 = img_reg_array_0_12_real;
        _zz_195 = img_reg_array_0_12_imag;
        _zz_196 = img_reg_array_1_12_real;
        _zz_197 = img_reg_array_1_12_imag;
        _zz_198 = img_reg_array_2_12_real;
        _zz_199 = img_reg_array_2_12_imag;
        _zz_200 = img_reg_array_3_12_real;
        _zz_201 = img_reg_array_3_12_imag;
        _zz_202 = img_reg_array_4_12_real;
        _zz_203 = img_reg_array_4_12_imag;
        _zz_204 = img_reg_array_5_12_real;
        _zz_205 = img_reg_array_5_12_imag;
        _zz_206 = img_reg_array_6_12_real;
        _zz_207 = img_reg_array_6_12_imag;
        _zz_208 = img_reg_array_7_12_real;
        _zz_209 = img_reg_array_7_12_imag;
        _zz_210 = img_reg_array_8_12_real;
        _zz_211 = img_reg_array_8_12_imag;
        _zz_212 = img_reg_array_9_12_real;
        _zz_213 = img_reg_array_9_12_imag;
        _zz_214 = img_reg_array_10_12_real;
        _zz_215 = img_reg_array_10_12_imag;
        _zz_216 = img_reg_array_11_12_real;
        _zz_217 = img_reg_array_11_12_imag;
        _zz_218 = img_reg_array_12_12_real;
        _zz_219 = img_reg_array_12_12_imag;
        _zz_220 = img_reg_array_13_12_real;
        _zz_221 = img_reg_array_13_12_imag;
        _zz_222 = img_reg_array_14_12_real;
        _zz_223 = img_reg_array_14_12_imag;
        _zz_224 = img_reg_array_15_12_real;
        _zz_225 = img_reg_array_15_12_imag;
        _zz_226 = img_reg_array_16_12_real;
        _zz_227 = img_reg_array_16_12_imag;
        _zz_228 = img_reg_array_17_12_real;
        _zz_229 = img_reg_array_17_12_imag;
        _zz_230 = img_reg_array_18_12_real;
        _zz_231 = img_reg_array_18_12_imag;
        _zz_232 = img_reg_array_19_12_real;
        _zz_233 = img_reg_array_19_12_imag;
        _zz_234 = img_reg_array_20_12_real;
        _zz_235 = img_reg_array_20_12_imag;
        _zz_236 = img_reg_array_21_12_real;
        _zz_237 = img_reg_array_21_12_imag;
        _zz_238 = img_reg_array_22_12_real;
        _zz_239 = img_reg_array_22_12_imag;
        _zz_240 = img_reg_array_23_12_real;
        _zz_241 = img_reg_array_23_12_imag;
        _zz_242 = img_reg_array_24_12_real;
        _zz_243 = img_reg_array_24_12_imag;
        _zz_244 = img_reg_array_25_12_real;
        _zz_245 = img_reg_array_25_12_imag;
        _zz_246 = img_reg_array_26_12_real;
        _zz_247 = img_reg_array_26_12_imag;
        _zz_248 = img_reg_array_27_12_real;
        _zz_249 = img_reg_array_27_12_imag;
        _zz_250 = img_reg_array_28_12_real;
        _zz_251 = img_reg_array_28_12_imag;
        _zz_252 = img_reg_array_29_12_real;
        _zz_253 = img_reg_array_29_12_imag;
        _zz_254 = img_reg_array_30_12_real;
        _zz_255 = img_reg_array_30_12_imag;
        _zz_256 = img_reg_array_31_12_real;
        _zz_257 = img_reg_array_31_12_imag;
        _zz_258 = img_reg_array_32_12_real;
        _zz_259 = img_reg_array_32_12_imag;
        _zz_260 = img_reg_array_33_12_real;
        _zz_261 = img_reg_array_33_12_imag;
        _zz_262 = img_reg_array_34_12_real;
        _zz_263 = img_reg_array_34_12_imag;
        _zz_264 = img_reg_array_35_12_real;
        _zz_265 = img_reg_array_35_12_imag;
        _zz_266 = img_reg_array_36_12_real;
        _zz_267 = img_reg_array_36_12_imag;
        _zz_268 = img_reg_array_37_12_real;
        _zz_269 = img_reg_array_37_12_imag;
        _zz_270 = img_reg_array_38_12_real;
        _zz_271 = img_reg_array_38_12_imag;
        _zz_272 = img_reg_array_39_12_real;
        _zz_273 = img_reg_array_39_12_imag;
        _zz_274 = img_reg_array_40_12_real;
        _zz_275 = img_reg_array_40_12_imag;
        _zz_276 = img_reg_array_41_12_real;
        _zz_277 = img_reg_array_41_12_imag;
        _zz_278 = img_reg_array_42_12_real;
        _zz_279 = img_reg_array_42_12_imag;
        _zz_280 = img_reg_array_43_12_real;
        _zz_281 = img_reg_array_43_12_imag;
        _zz_282 = img_reg_array_44_12_real;
        _zz_283 = img_reg_array_44_12_imag;
        _zz_284 = img_reg_array_45_12_real;
        _zz_285 = img_reg_array_45_12_imag;
        _zz_286 = img_reg_array_46_12_real;
        _zz_287 = img_reg_array_46_12_imag;
        _zz_288 = img_reg_array_47_12_real;
        _zz_289 = img_reg_array_47_12_imag;
        _zz_290 = img_reg_array_48_12_real;
        _zz_291 = img_reg_array_48_12_imag;
        _zz_292 = img_reg_array_49_12_real;
        _zz_293 = img_reg_array_49_12_imag;
        _zz_294 = img_reg_array_50_12_real;
        _zz_295 = img_reg_array_50_12_imag;
        _zz_296 = img_reg_array_51_12_real;
        _zz_297 = img_reg_array_51_12_imag;
        _zz_298 = img_reg_array_52_12_real;
        _zz_299 = img_reg_array_52_12_imag;
        _zz_300 = img_reg_array_53_12_real;
        _zz_301 = img_reg_array_53_12_imag;
        _zz_302 = img_reg_array_54_12_real;
        _zz_303 = img_reg_array_54_12_imag;
        _zz_304 = img_reg_array_55_12_real;
        _zz_305 = img_reg_array_55_12_imag;
        _zz_306 = img_reg_array_56_12_real;
        _zz_307 = img_reg_array_56_12_imag;
        _zz_308 = img_reg_array_57_12_real;
        _zz_309 = img_reg_array_57_12_imag;
        _zz_310 = img_reg_array_58_12_real;
        _zz_311 = img_reg_array_58_12_imag;
        _zz_312 = img_reg_array_59_12_real;
        _zz_313 = img_reg_array_59_12_imag;
        _zz_314 = img_reg_array_60_12_real;
        _zz_315 = img_reg_array_60_12_imag;
        _zz_316 = img_reg_array_61_12_real;
        _zz_317 = img_reg_array_61_12_imag;
        _zz_318 = img_reg_array_62_12_real;
        _zz_319 = img_reg_array_62_12_imag;
        _zz_320 = img_reg_array_63_12_real;
        _zz_321 = img_reg_array_63_12_imag;
      end
      6'b001101 : begin
        _zz_194 = img_reg_array_0_13_real;
        _zz_195 = img_reg_array_0_13_imag;
        _zz_196 = img_reg_array_1_13_real;
        _zz_197 = img_reg_array_1_13_imag;
        _zz_198 = img_reg_array_2_13_real;
        _zz_199 = img_reg_array_2_13_imag;
        _zz_200 = img_reg_array_3_13_real;
        _zz_201 = img_reg_array_3_13_imag;
        _zz_202 = img_reg_array_4_13_real;
        _zz_203 = img_reg_array_4_13_imag;
        _zz_204 = img_reg_array_5_13_real;
        _zz_205 = img_reg_array_5_13_imag;
        _zz_206 = img_reg_array_6_13_real;
        _zz_207 = img_reg_array_6_13_imag;
        _zz_208 = img_reg_array_7_13_real;
        _zz_209 = img_reg_array_7_13_imag;
        _zz_210 = img_reg_array_8_13_real;
        _zz_211 = img_reg_array_8_13_imag;
        _zz_212 = img_reg_array_9_13_real;
        _zz_213 = img_reg_array_9_13_imag;
        _zz_214 = img_reg_array_10_13_real;
        _zz_215 = img_reg_array_10_13_imag;
        _zz_216 = img_reg_array_11_13_real;
        _zz_217 = img_reg_array_11_13_imag;
        _zz_218 = img_reg_array_12_13_real;
        _zz_219 = img_reg_array_12_13_imag;
        _zz_220 = img_reg_array_13_13_real;
        _zz_221 = img_reg_array_13_13_imag;
        _zz_222 = img_reg_array_14_13_real;
        _zz_223 = img_reg_array_14_13_imag;
        _zz_224 = img_reg_array_15_13_real;
        _zz_225 = img_reg_array_15_13_imag;
        _zz_226 = img_reg_array_16_13_real;
        _zz_227 = img_reg_array_16_13_imag;
        _zz_228 = img_reg_array_17_13_real;
        _zz_229 = img_reg_array_17_13_imag;
        _zz_230 = img_reg_array_18_13_real;
        _zz_231 = img_reg_array_18_13_imag;
        _zz_232 = img_reg_array_19_13_real;
        _zz_233 = img_reg_array_19_13_imag;
        _zz_234 = img_reg_array_20_13_real;
        _zz_235 = img_reg_array_20_13_imag;
        _zz_236 = img_reg_array_21_13_real;
        _zz_237 = img_reg_array_21_13_imag;
        _zz_238 = img_reg_array_22_13_real;
        _zz_239 = img_reg_array_22_13_imag;
        _zz_240 = img_reg_array_23_13_real;
        _zz_241 = img_reg_array_23_13_imag;
        _zz_242 = img_reg_array_24_13_real;
        _zz_243 = img_reg_array_24_13_imag;
        _zz_244 = img_reg_array_25_13_real;
        _zz_245 = img_reg_array_25_13_imag;
        _zz_246 = img_reg_array_26_13_real;
        _zz_247 = img_reg_array_26_13_imag;
        _zz_248 = img_reg_array_27_13_real;
        _zz_249 = img_reg_array_27_13_imag;
        _zz_250 = img_reg_array_28_13_real;
        _zz_251 = img_reg_array_28_13_imag;
        _zz_252 = img_reg_array_29_13_real;
        _zz_253 = img_reg_array_29_13_imag;
        _zz_254 = img_reg_array_30_13_real;
        _zz_255 = img_reg_array_30_13_imag;
        _zz_256 = img_reg_array_31_13_real;
        _zz_257 = img_reg_array_31_13_imag;
        _zz_258 = img_reg_array_32_13_real;
        _zz_259 = img_reg_array_32_13_imag;
        _zz_260 = img_reg_array_33_13_real;
        _zz_261 = img_reg_array_33_13_imag;
        _zz_262 = img_reg_array_34_13_real;
        _zz_263 = img_reg_array_34_13_imag;
        _zz_264 = img_reg_array_35_13_real;
        _zz_265 = img_reg_array_35_13_imag;
        _zz_266 = img_reg_array_36_13_real;
        _zz_267 = img_reg_array_36_13_imag;
        _zz_268 = img_reg_array_37_13_real;
        _zz_269 = img_reg_array_37_13_imag;
        _zz_270 = img_reg_array_38_13_real;
        _zz_271 = img_reg_array_38_13_imag;
        _zz_272 = img_reg_array_39_13_real;
        _zz_273 = img_reg_array_39_13_imag;
        _zz_274 = img_reg_array_40_13_real;
        _zz_275 = img_reg_array_40_13_imag;
        _zz_276 = img_reg_array_41_13_real;
        _zz_277 = img_reg_array_41_13_imag;
        _zz_278 = img_reg_array_42_13_real;
        _zz_279 = img_reg_array_42_13_imag;
        _zz_280 = img_reg_array_43_13_real;
        _zz_281 = img_reg_array_43_13_imag;
        _zz_282 = img_reg_array_44_13_real;
        _zz_283 = img_reg_array_44_13_imag;
        _zz_284 = img_reg_array_45_13_real;
        _zz_285 = img_reg_array_45_13_imag;
        _zz_286 = img_reg_array_46_13_real;
        _zz_287 = img_reg_array_46_13_imag;
        _zz_288 = img_reg_array_47_13_real;
        _zz_289 = img_reg_array_47_13_imag;
        _zz_290 = img_reg_array_48_13_real;
        _zz_291 = img_reg_array_48_13_imag;
        _zz_292 = img_reg_array_49_13_real;
        _zz_293 = img_reg_array_49_13_imag;
        _zz_294 = img_reg_array_50_13_real;
        _zz_295 = img_reg_array_50_13_imag;
        _zz_296 = img_reg_array_51_13_real;
        _zz_297 = img_reg_array_51_13_imag;
        _zz_298 = img_reg_array_52_13_real;
        _zz_299 = img_reg_array_52_13_imag;
        _zz_300 = img_reg_array_53_13_real;
        _zz_301 = img_reg_array_53_13_imag;
        _zz_302 = img_reg_array_54_13_real;
        _zz_303 = img_reg_array_54_13_imag;
        _zz_304 = img_reg_array_55_13_real;
        _zz_305 = img_reg_array_55_13_imag;
        _zz_306 = img_reg_array_56_13_real;
        _zz_307 = img_reg_array_56_13_imag;
        _zz_308 = img_reg_array_57_13_real;
        _zz_309 = img_reg_array_57_13_imag;
        _zz_310 = img_reg_array_58_13_real;
        _zz_311 = img_reg_array_58_13_imag;
        _zz_312 = img_reg_array_59_13_real;
        _zz_313 = img_reg_array_59_13_imag;
        _zz_314 = img_reg_array_60_13_real;
        _zz_315 = img_reg_array_60_13_imag;
        _zz_316 = img_reg_array_61_13_real;
        _zz_317 = img_reg_array_61_13_imag;
        _zz_318 = img_reg_array_62_13_real;
        _zz_319 = img_reg_array_62_13_imag;
        _zz_320 = img_reg_array_63_13_real;
        _zz_321 = img_reg_array_63_13_imag;
      end
      6'b001110 : begin
        _zz_194 = img_reg_array_0_14_real;
        _zz_195 = img_reg_array_0_14_imag;
        _zz_196 = img_reg_array_1_14_real;
        _zz_197 = img_reg_array_1_14_imag;
        _zz_198 = img_reg_array_2_14_real;
        _zz_199 = img_reg_array_2_14_imag;
        _zz_200 = img_reg_array_3_14_real;
        _zz_201 = img_reg_array_3_14_imag;
        _zz_202 = img_reg_array_4_14_real;
        _zz_203 = img_reg_array_4_14_imag;
        _zz_204 = img_reg_array_5_14_real;
        _zz_205 = img_reg_array_5_14_imag;
        _zz_206 = img_reg_array_6_14_real;
        _zz_207 = img_reg_array_6_14_imag;
        _zz_208 = img_reg_array_7_14_real;
        _zz_209 = img_reg_array_7_14_imag;
        _zz_210 = img_reg_array_8_14_real;
        _zz_211 = img_reg_array_8_14_imag;
        _zz_212 = img_reg_array_9_14_real;
        _zz_213 = img_reg_array_9_14_imag;
        _zz_214 = img_reg_array_10_14_real;
        _zz_215 = img_reg_array_10_14_imag;
        _zz_216 = img_reg_array_11_14_real;
        _zz_217 = img_reg_array_11_14_imag;
        _zz_218 = img_reg_array_12_14_real;
        _zz_219 = img_reg_array_12_14_imag;
        _zz_220 = img_reg_array_13_14_real;
        _zz_221 = img_reg_array_13_14_imag;
        _zz_222 = img_reg_array_14_14_real;
        _zz_223 = img_reg_array_14_14_imag;
        _zz_224 = img_reg_array_15_14_real;
        _zz_225 = img_reg_array_15_14_imag;
        _zz_226 = img_reg_array_16_14_real;
        _zz_227 = img_reg_array_16_14_imag;
        _zz_228 = img_reg_array_17_14_real;
        _zz_229 = img_reg_array_17_14_imag;
        _zz_230 = img_reg_array_18_14_real;
        _zz_231 = img_reg_array_18_14_imag;
        _zz_232 = img_reg_array_19_14_real;
        _zz_233 = img_reg_array_19_14_imag;
        _zz_234 = img_reg_array_20_14_real;
        _zz_235 = img_reg_array_20_14_imag;
        _zz_236 = img_reg_array_21_14_real;
        _zz_237 = img_reg_array_21_14_imag;
        _zz_238 = img_reg_array_22_14_real;
        _zz_239 = img_reg_array_22_14_imag;
        _zz_240 = img_reg_array_23_14_real;
        _zz_241 = img_reg_array_23_14_imag;
        _zz_242 = img_reg_array_24_14_real;
        _zz_243 = img_reg_array_24_14_imag;
        _zz_244 = img_reg_array_25_14_real;
        _zz_245 = img_reg_array_25_14_imag;
        _zz_246 = img_reg_array_26_14_real;
        _zz_247 = img_reg_array_26_14_imag;
        _zz_248 = img_reg_array_27_14_real;
        _zz_249 = img_reg_array_27_14_imag;
        _zz_250 = img_reg_array_28_14_real;
        _zz_251 = img_reg_array_28_14_imag;
        _zz_252 = img_reg_array_29_14_real;
        _zz_253 = img_reg_array_29_14_imag;
        _zz_254 = img_reg_array_30_14_real;
        _zz_255 = img_reg_array_30_14_imag;
        _zz_256 = img_reg_array_31_14_real;
        _zz_257 = img_reg_array_31_14_imag;
        _zz_258 = img_reg_array_32_14_real;
        _zz_259 = img_reg_array_32_14_imag;
        _zz_260 = img_reg_array_33_14_real;
        _zz_261 = img_reg_array_33_14_imag;
        _zz_262 = img_reg_array_34_14_real;
        _zz_263 = img_reg_array_34_14_imag;
        _zz_264 = img_reg_array_35_14_real;
        _zz_265 = img_reg_array_35_14_imag;
        _zz_266 = img_reg_array_36_14_real;
        _zz_267 = img_reg_array_36_14_imag;
        _zz_268 = img_reg_array_37_14_real;
        _zz_269 = img_reg_array_37_14_imag;
        _zz_270 = img_reg_array_38_14_real;
        _zz_271 = img_reg_array_38_14_imag;
        _zz_272 = img_reg_array_39_14_real;
        _zz_273 = img_reg_array_39_14_imag;
        _zz_274 = img_reg_array_40_14_real;
        _zz_275 = img_reg_array_40_14_imag;
        _zz_276 = img_reg_array_41_14_real;
        _zz_277 = img_reg_array_41_14_imag;
        _zz_278 = img_reg_array_42_14_real;
        _zz_279 = img_reg_array_42_14_imag;
        _zz_280 = img_reg_array_43_14_real;
        _zz_281 = img_reg_array_43_14_imag;
        _zz_282 = img_reg_array_44_14_real;
        _zz_283 = img_reg_array_44_14_imag;
        _zz_284 = img_reg_array_45_14_real;
        _zz_285 = img_reg_array_45_14_imag;
        _zz_286 = img_reg_array_46_14_real;
        _zz_287 = img_reg_array_46_14_imag;
        _zz_288 = img_reg_array_47_14_real;
        _zz_289 = img_reg_array_47_14_imag;
        _zz_290 = img_reg_array_48_14_real;
        _zz_291 = img_reg_array_48_14_imag;
        _zz_292 = img_reg_array_49_14_real;
        _zz_293 = img_reg_array_49_14_imag;
        _zz_294 = img_reg_array_50_14_real;
        _zz_295 = img_reg_array_50_14_imag;
        _zz_296 = img_reg_array_51_14_real;
        _zz_297 = img_reg_array_51_14_imag;
        _zz_298 = img_reg_array_52_14_real;
        _zz_299 = img_reg_array_52_14_imag;
        _zz_300 = img_reg_array_53_14_real;
        _zz_301 = img_reg_array_53_14_imag;
        _zz_302 = img_reg_array_54_14_real;
        _zz_303 = img_reg_array_54_14_imag;
        _zz_304 = img_reg_array_55_14_real;
        _zz_305 = img_reg_array_55_14_imag;
        _zz_306 = img_reg_array_56_14_real;
        _zz_307 = img_reg_array_56_14_imag;
        _zz_308 = img_reg_array_57_14_real;
        _zz_309 = img_reg_array_57_14_imag;
        _zz_310 = img_reg_array_58_14_real;
        _zz_311 = img_reg_array_58_14_imag;
        _zz_312 = img_reg_array_59_14_real;
        _zz_313 = img_reg_array_59_14_imag;
        _zz_314 = img_reg_array_60_14_real;
        _zz_315 = img_reg_array_60_14_imag;
        _zz_316 = img_reg_array_61_14_real;
        _zz_317 = img_reg_array_61_14_imag;
        _zz_318 = img_reg_array_62_14_real;
        _zz_319 = img_reg_array_62_14_imag;
        _zz_320 = img_reg_array_63_14_real;
        _zz_321 = img_reg_array_63_14_imag;
      end
      6'b001111 : begin
        _zz_194 = img_reg_array_0_15_real;
        _zz_195 = img_reg_array_0_15_imag;
        _zz_196 = img_reg_array_1_15_real;
        _zz_197 = img_reg_array_1_15_imag;
        _zz_198 = img_reg_array_2_15_real;
        _zz_199 = img_reg_array_2_15_imag;
        _zz_200 = img_reg_array_3_15_real;
        _zz_201 = img_reg_array_3_15_imag;
        _zz_202 = img_reg_array_4_15_real;
        _zz_203 = img_reg_array_4_15_imag;
        _zz_204 = img_reg_array_5_15_real;
        _zz_205 = img_reg_array_5_15_imag;
        _zz_206 = img_reg_array_6_15_real;
        _zz_207 = img_reg_array_6_15_imag;
        _zz_208 = img_reg_array_7_15_real;
        _zz_209 = img_reg_array_7_15_imag;
        _zz_210 = img_reg_array_8_15_real;
        _zz_211 = img_reg_array_8_15_imag;
        _zz_212 = img_reg_array_9_15_real;
        _zz_213 = img_reg_array_9_15_imag;
        _zz_214 = img_reg_array_10_15_real;
        _zz_215 = img_reg_array_10_15_imag;
        _zz_216 = img_reg_array_11_15_real;
        _zz_217 = img_reg_array_11_15_imag;
        _zz_218 = img_reg_array_12_15_real;
        _zz_219 = img_reg_array_12_15_imag;
        _zz_220 = img_reg_array_13_15_real;
        _zz_221 = img_reg_array_13_15_imag;
        _zz_222 = img_reg_array_14_15_real;
        _zz_223 = img_reg_array_14_15_imag;
        _zz_224 = img_reg_array_15_15_real;
        _zz_225 = img_reg_array_15_15_imag;
        _zz_226 = img_reg_array_16_15_real;
        _zz_227 = img_reg_array_16_15_imag;
        _zz_228 = img_reg_array_17_15_real;
        _zz_229 = img_reg_array_17_15_imag;
        _zz_230 = img_reg_array_18_15_real;
        _zz_231 = img_reg_array_18_15_imag;
        _zz_232 = img_reg_array_19_15_real;
        _zz_233 = img_reg_array_19_15_imag;
        _zz_234 = img_reg_array_20_15_real;
        _zz_235 = img_reg_array_20_15_imag;
        _zz_236 = img_reg_array_21_15_real;
        _zz_237 = img_reg_array_21_15_imag;
        _zz_238 = img_reg_array_22_15_real;
        _zz_239 = img_reg_array_22_15_imag;
        _zz_240 = img_reg_array_23_15_real;
        _zz_241 = img_reg_array_23_15_imag;
        _zz_242 = img_reg_array_24_15_real;
        _zz_243 = img_reg_array_24_15_imag;
        _zz_244 = img_reg_array_25_15_real;
        _zz_245 = img_reg_array_25_15_imag;
        _zz_246 = img_reg_array_26_15_real;
        _zz_247 = img_reg_array_26_15_imag;
        _zz_248 = img_reg_array_27_15_real;
        _zz_249 = img_reg_array_27_15_imag;
        _zz_250 = img_reg_array_28_15_real;
        _zz_251 = img_reg_array_28_15_imag;
        _zz_252 = img_reg_array_29_15_real;
        _zz_253 = img_reg_array_29_15_imag;
        _zz_254 = img_reg_array_30_15_real;
        _zz_255 = img_reg_array_30_15_imag;
        _zz_256 = img_reg_array_31_15_real;
        _zz_257 = img_reg_array_31_15_imag;
        _zz_258 = img_reg_array_32_15_real;
        _zz_259 = img_reg_array_32_15_imag;
        _zz_260 = img_reg_array_33_15_real;
        _zz_261 = img_reg_array_33_15_imag;
        _zz_262 = img_reg_array_34_15_real;
        _zz_263 = img_reg_array_34_15_imag;
        _zz_264 = img_reg_array_35_15_real;
        _zz_265 = img_reg_array_35_15_imag;
        _zz_266 = img_reg_array_36_15_real;
        _zz_267 = img_reg_array_36_15_imag;
        _zz_268 = img_reg_array_37_15_real;
        _zz_269 = img_reg_array_37_15_imag;
        _zz_270 = img_reg_array_38_15_real;
        _zz_271 = img_reg_array_38_15_imag;
        _zz_272 = img_reg_array_39_15_real;
        _zz_273 = img_reg_array_39_15_imag;
        _zz_274 = img_reg_array_40_15_real;
        _zz_275 = img_reg_array_40_15_imag;
        _zz_276 = img_reg_array_41_15_real;
        _zz_277 = img_reg_array_41_15_imag;
        _zz_278 = img_reg_array_42_15_real;
        _zz_279 = img_reg_array_42_15_imag;
        _zz_280 = img_reg_array_43_15_real;
        _zz_281 = img_reg_array_43_15_imag;
        _zz_282 = img_reg_array_44_15_real;
        _zz_283 = img_reg_array_44_15_imag;
        _zz_284 = img_reg_array_45_15_real;
        _zz_285 = img_reg_array_45_15_imag;
        _zz_286 = img_reg_array_46_15_real;
        _zz_287 = img_reg_array_46_15_imag;
        _zz_288 = img_reg_array_47_15_real;
        _zz_289 = img_reg_array_47_15_imag;
        _zz_290 = img_reg_array_48_15_real;
        _zz_291 = img_reg_array_48_15_imag;
        _zz_292 = img_reg_array_49_15_real;
        _zz_293 = img_reg_array_49_15_imag;
        _zz_294 = img_reg_array_50_15_real;
        _zz_295 = img_reg_array_50_15_imag;
        _zz_296 = img_reg_array_51_15_real;
        _zz_297 = img_reg_array_51_15_imag;
        _zz_298 = img_reg_array_52_15_real;
        _zz_299 = img_reg_array_52_15_imag;
        _zz_300 = img_reg_array_53_15_real;
        _zz_301 = img_reg_array_53_15_imag;
        _zz_302 = img_reg_array_54_15_real;
        _zz_303 = img_reg_array_54_15_imag;
        _zz_304 = img_reg_array_55_15_real;
        _zz_305 = img_reg_array_55_15_imag;
        _zz_306 = img_reg_array_56_15_real;
        _zz_307 = img_reg_array_56_15_imag;
        _zz_308 = img_reg_array_57_15_real;
        _zz_309 = img_reg_array_57_15_imag;
        _zz_310 = img_reg_array_58_15_real;
        _zz_311 = img_reg_array_58_15_imag;
        _zz_312 = img_reg_array_59_15_real;
        _zz_313 = img_reg_array_59_15_imag;
        _zz_314 = img_reg_array_60_15_real;
        _zz_315 = img_reg_array_60_15_imag;
        _zz_316 = img_reg_array_61_15_real;
        _zz_317 = img_reg_array_61_15_imag;
        _zz_318 = img_reg_array_62_15_real;
        _zz_319 = img_reg_array_62_15_imag;
        _zz_320 = img_reg_array_63_15_real;
        _zz_321 = img_reg_array_63_15_imag;
      end
      6'b010000 : begin
        _zz_194 = img_reg_array_0_16_real;
        _zz_195 = img_reg_array_0_16_imag;
        _zz_196 = img_reg_array_1_16_real;
        _zz_197 = img_reg_array_1_16_imag;
        _zz_198 = img_reg_array_2_16_real;
        _zz_199 = img_reg_array_2_16_imag;
        _zz_200 = img_reg_array_3_16_real;
        _zz_201 = img_reg_array_3_16_imag;
        _zz_202 = img_reg_array_4_16_real;
        _zz_203 = img_reg_array_4_16_imag;
        _zz_204 = img_reg_array_5_16_real;
        _zz_205 = img_reg_array_5_16_imag;
        _zz_206 = img_reg_array_6_16_real;
        _zz_207 = img_reg_array_6_16_imag;
        _zz_208 = img_reg_array_7_16_real;
        _zz_209 = img_reg_array_7_16_imag;
        _zz_210 = img_reg_array_8_16_real;
        _zz_211 = img_reg_array_8_16_imag;
        _zz_212 = img_reg_array_9_16_real;
        _zz_213 = img_reg_array_9_16_imag;
        _zz_214 = img_reg_array_10_16_real;
        _zz_215 = img_reg_array_10_16_imag;
        _zz_216 = img_reg_array_11_16_real;
        _zz_217 = img_reg_array_11_16_imag;
        _zz_218 = img_reg_array_12_16_real;
        _zz_219 = img_reg_array_12_16_imag;
        _zz_220 = img_reg_array_13_16_real;
        _zz_221 = img_reg_array_13_16_imag;
        _zz_222 = img_reg_array_14_16_real;
        _zz_223 = img_reg_array_14_16_imag;
        _zz_224 = img_reg_array_15_16_real;
        _zz_225 = img_reg_array_15_16_imag;
        _zz_226 = img_reg_array_16_16_real;
        _zz_227 = img_reg_array_16_16_imag;
        _zz_228 = img_reg_array_17_16_real;
        _zz_229 = img_reg_array_17_16_imag;
        _zz_230 = img_reg_array_18_16_real;
        _zz_231 = img_reg_array_18_16_imag;
        _zz_232 = img_reg_array_19_16_real;
        _zz_233 = img_reg_array_19_16_imag;
        _zz_234 = img_reg_array_20_16_real;
        _zz_235 = img_reg_array_20_16_imag;
        _zz_236 = img_reg_array_21_16_real;
        _zz_237 = img_reg_array_21_16_imag;
        _zz_238 = img_reg_array_22_16_real;
        _zz_239 = img_reg_array_22_16_imag;
        _zz_240 = img_reg_array_23_16_real;
        _zz_241 = img_reg_array_23_16_imag;
        _zz_242 = img_reg_array_24_16_real;
        _zz_243 = img_reg_array_24_16_imag;
        _zz_244 = img_reg_array_25_16_real;
        _zz_245 = img_reg_array_25_16_imag;
        _zz_246 = img_reg_array_26_16_real;
        _zz_247 = img_reg_array_26_16_imag;
        _zz_248 = img_reg_array_27_16_real;
        _zz_249 = img_reg_array_27_16_imag;
        _zz_250 = img_reg_array_28_16_real;
        _zz_251 = img_reg_array_28_16_imag;
        _zz_252 = img_reg_array_29_16_real;
        _zz_253 = img_reg_array_29_16_imag;
        _zz_254 = img_reg_array_30_16_real;
        _zz_255 = img_reg_array_30_16_imag;
        _zz_256 = img_reg_array_31_16_real;
        _zz_257 = img_reg_array_31_16_imag;
        _zz_258 = img_reg_array_32_16_real;
        _zz_259 = img_reg_array_32_16_imag;
        _zz_260 = img_reg_array_33_16_real;
        _zz_261 = img_reg_array_33_16_imag;
        _zz_262 = img_reg_array_34_16_real;
        _zz_263 = img_reg_array_34_16_imag;
        _zz_264 = img_reg_array_35_16_real;
        _zz_265 = img_reg_array_35_16_imag;
        _zz_266 = img_reg_array_36_16_real;
        _zz_267 = img_reg_array_36_16_imag;
        _zz_268 = img_reg_array_37_16_real;
        _zz_269 = img_reg_array_37_16_imag;
        _zz_270 = img_reg_array_38_16_real;
        _zz_271 = img_reg_array_38_16_imag;
        _zz_272 = img_reg_array_39_16_real;
        _zz_273 = img_reg_array_39_16_imag;
        _zz_274 = img_reg_array_40_16_real;
        _zz_275 = img_reg_array_40_16_imag;
        _zz_276 = img_reg_array_41_16_real;
        _zz_277 = img_reg_array_41_16_imag;
        _zz_278 = img_reg_array_42_16_real;
        _zz_279 = img_reg_array_42_16_imag;
        _zz_280 = img_reg_array_43_16_real;
        _zz_281 = img_reg_array_43_16_imag;
        _zz_282 = img_reg_array_44_16_real;
        _zz_283 = img_reg_array_44_16_imag;
        _zz_284 = img_reg_array_45_16_real;
        _zz_285 = img_reg_array_45_16_imag;
        _zz_286 = img_reg_array_46_16_real;
        _zz_287 = img_reg_array_46_16_imag;
        _zz_288 = img_reg_array_47_16_real;
        _zz_289 = img_reg_array_47_16_imag;
        _zz_290 = img_reg_array_48_16_real;
        _zz_291 = img_reg_array_48_16_imag;
        _zz_292 = img_reg_array_49_16_real;
        _zz_293 = img_reg_array_49_16_imag;
        _zz_294 = img_reg_array_50_16_real;
        _zz_295 = img_reg_array_50_16_imag;
        _zz_296 = img_reg_array_51_16_real;
        _zz_297 = img_reg_array_51_16_imag;
        _zz_298 = img_reg_array_52_16_real;
        _zz_299 = img_reg_array_52_16_imag;
        _zz_300 = img_reg_array_53_16_real;
        _zz_301 = img_reg_array_53_16_imag;
        _zz_302 = img_reg_array_54_16_real;
        _zz_303 = img_reg_array_54_16_imag;
        _zz_304 = img_reg_array_55_16_real;
        _zz_305 = img_reg_array_55_16_imag;
        _zz_306 = img_reg_array_56_16_real;
        _zz_307 = img_reg_array_56_16_imag;
        _zz_308 = img_reg_array_57_16_real;
        _zz_309 = img_reg_array_57_16_imag;
        _zz_310 = img_reg_array_58_16_real;
        _zz_311 = img_reg_array_58_16_imag;
        _zz_312 = img_reg_array_59_16_real;
        _zz_313 = img_reg_array_59_16_imag;
        _zz_314 = img_reg_array_60_16_real;
        _zz_315 = img_reg_array_60_16_imag;
        _zz_316 = img_reg_array_61_16_real;
        _zz_317 = img_reg_array_61_16_imag;
        _zz_318 = img_reg_array_62_16_real;
        _zz_319 = img_reg_array_62_16_imag;
        _zz_320 = img_reg_array_63_16_real;
        _zz_321 = img_reg_array_63_16_imag;
      end
      6'b010001 : begin
        _zz_194 = img_reg_array_0_17_real;
        _zz_195 = img_reg_array_0_17_imag;
        _zz_196 = img_reg_array_1_17_real;
        _zz_197 = img_reg_array_1_17_imag;
        _zz_198 = img_reg_array_2_17_real;
        _zz_199 = img_reg_array_2_17_imag;
        _zz_200 = img_reg_array_3_17_real;
        _zz_201 = img_reg_array_3_17_imag;
        _zz_202 = img_reg_array_4_17_real;
        _zz_203 = img_reg_array_4_17_imag;
        _zz_204 = img_reg_array_5_17_real;
        _zz_205 = img_reg_array_5_17_imag;
        _zz_206 = img_reg_array_6_17_real;
        _zz_207 = img_reg_array_6_17_imag;
        _zz_208 = img_reg_array_7_17_real;
        _zz_209 = img_reg_array_7_17_imag;
        _zz_210 = img_reg_array_8_17_real;
        _zz_211 = img_reg_array_8_17_imag;
        _zz_212 = img_reg_array_9_17_real;
        _zz_213 = img_reg_array_9_17_imag;
        _zz_214 = img_reg_array_10_17_real;
        _zz_215 = img_reg_array_10_17_imag;
        _zz_216 = img_reg_array_11_17_real;
        _zz_217 = img_reg_array_11_17_imag;
        _zz_218 = img_reg_array_12_17_real;
        _zz_219 = img_reg_array_12_17_imag;
        _zz_220 = img_reg_array_13_17_real;
        _zz_221 = img_reg_array_13_17_imag;
        _zz_222 = img_reg_array_14_17_real;
        _zz_223 = img_reg_array_14_17_imag;
        _zz_224 = img_reg_array_15_17_real;
        _zz_225 = img_reg_array_15_17_imag;
        _zz_226 = img_reg_array_16_17_real;
        _zz_227 = img_reg_array_16_17_imag;
        _zz_228 = img_reg_array_17_17_real;
        _zz_229 = img_reg_array_17_17_imag;
        _zz_230 = img_reg_array_18_17_real;
        _zz_231 = img_reg_array_18_17_imag;
        _zz_232 = img_reg_array_19_17_real;
        _zz_233 = img_reg_array_19_17_imag;
        _zz_234 = img_reg_array_20_17_real;
        _zz_235 = img_reg_array_20_17_imag;
        _zz_236 = img_reg_array_21_17_real;
        _zz_237 = img_reg_array_21_17_imag;
        _zz_238 = img_reg_array_22_17_real;
        _zz_239 = img_reg_array_22_17_imag;
        _zz_240 = img_reg_array_23_17_real;
        _zz_241 = img_reg_array_23_17_imag;
        _zz_242 = img_reg_array_24_17_real;
        _zz_243 = img_reg_array_24_17_imag;
        _zz_244 = img_reg_array_25_17_real;
        _zz_245 = img_reg_array_25_17_imag;
        _zz_246 = img_reg_array_26_17_real;
        _zz_247 = img_reg_array_26_17_imag;
        _zz_248 = img_reg_array_27_17_real;
        _zz_249 = img_reg_array_27_17_imag;
        _zz_250 = img_reg_array_28_17_real;
        _zz_251 = img_reg_array_28_17_imag;
        _zz_252 = img_reg_array_29_17_real;
        _zz_253 = img_reg_array_29_17_imag;
        _zz_254 = img_reg_array_30_17_real;
        _zz_255 = img_reg_array_30_17_imag;
        _zz_256 = img_reg_array_31_17_real;
        _zz_257 = img_reg_array_31_17_imag;
        _zz_258 = img_reg_array_32_17_real;
        _zz_259 = img_reg_array_32_17_imag;
        _zz_260 = img_reg_array_33_17_real;
        _zz_261 = img_reg_array_33_17_imag;
        _zz_262 = img_reg_array_34_17_real;
        _zz_263 = img_reg_array_34_17_imag;
        _zz_264 = img_reg_array_35_17_real;
        _zz_265 = img_reg_array_35_17_imag;
        _zz_266 = img_reg_array_36_17_real;
        _zz_267 = img_reg_array_36_17_imag;
        _zz_268 = img_reg_array_37_17_real;
        _zz_269 = img_reg_array_37_17_imag;
        _zz_270 = img_reg_array_38_17_real;
        _zz_271 = img_reg_array_38_17_imag;
        _zz_272 = img_reg_array_39_17_real;
        _zz_273 = img_reg_array_39_17_imag;
        _zz_274 = img_reg_array_40_17_real;
        _zz_275 = img_reg_array_40_17_imag;
        _zz_276 = img_reg_array_41_17_real;
        _zz_277 = img_reg_array_41_17_imag;
        _zz_278 = img_reg_array_42_17_real;
        _zz_279 = img_reg_array_42_17_imag;
        _zz_280 = img_reg_array_43_17_real;
        _zz_281 = img_reg_array_43_17_imag;
        _zz_282 = img_reg_array_44_17_real;
        _zz_283 = img_reg_array_44_17_imag;
        _zz_284 = img_reg_array_45_17_real;
        _zz_285 = img_reg_array_45_17_imag;
        _zz_286 = img_reg_array_46_17_real;
        _zz_287 = img_reg_array_46_17_imag;
        _zz_288 = img_reg_array_47_17_real;
        _zz_289 = img_reg_array_47_17_imag;
        _zz_290 = img_reg_array_48_17_real;
        _zz_291 = img_reg_array_48_17_imag;
        _zz_292 = img_reg_array_49_17_real;
        _zz_293 = img_reg_array_49_17_imag;
        _zz_294 = img_reg_array_50_17_real;
        _zz_295 = img_reg_array_50_17_imag;
        _zz_296 = img_reg_array_51_17_real;
        _zz_297 = img_reg_array_51_17_imag;
        _zz_298 = img_reg_array_52_17_real;
        _zz_299 = img_reg_array_52_17_imag;
        _zz_300 = img_reg_array_53_17_real;
        _zz_301 = img_reg_array_53_17_imag;
        _zz_302 = img_reg_array_54_17_real;
        _zz_303 = img_reg_array_54_17_imag;
        _zz_304 = img_reg_array_55_17_real;
        _zz_305 = img_reg_array_55_17_imag;
        _zz_306 = img_reg_array_56_17_real;
        _zz_307 = img_reg_array_56_17_imag;
        _zz_308 = img_reg_array_57_17_real;
        _zz_309 = img_reg_array_57_17_imag;
        _zz_310 = img_reg_array_58_17_real;
        _zz_311 = img_reg_array_58_17_imag;
        _zz_312 = img_reg_array_59_17_real;
        _zz_313 = img_reg_array_59_17_imag;
        _zz_314 = img_reg_array_60_17_real;
        _zz_315 = img_reg_array_60_17_imag;
        _zz_316 = img_reg_array_61_17_real;
        _zz_317 = img_reg_array_61_17_imag;
        _zz_318 = img_reg_array_62_17_real;
        _zz_319 = img_reg_array_62_17_imag;
        _zz_320 = img_reg_array_63_17_real;
        _zz_321 = img_reg_array_63_17_imag;
      end
      6'b010010 : begin
        _zz_194 = img_reg_array_0_18_real;
        _zz_195 = img_reg_array_0_18_imag;
        _zz_196 = img_reg_array_1_18_real;
        _zz_197 = img_reg_array_1_18_imag;
        _zz_198 = img_reg_array_2_18_real;
        _zz_199 = img_reg_array_2_18_imag;
        _zz_200 = img_reg_array_3_18_real;
        _zz_201 = img_reg_array_3_18_imag;
        _zz_202 = img_reg_array_4_18_real;
        _zz_203 = img_reg_array_4_18_imag;
        _zz_204 = img_reg_array_5_18_real;
        _zz_205 = img_reg_array_5_18_imag;
        _zz_206 = img_reg_array_6_18_real;
        _zz_207 = img_reg_array_6_18_imag;
        _zz_208 = img_reg_array_7_18_real;
        _zz_209 = img_reg_array_7_18_imag;
        _zz_210 = img_reg_array_8_18_real;
        _zz_211 = img_reg_array_8_18_imag;
        _zz_212 = img_reg_array_9_18_real;
        _zz_213 = img_reg_array_9_18_imag;
        _zz_214 = img_reg_array_10_18_real;
        _zz_215 = img_reg_array_10_18_imag;
        _zz_216 = img_reg_array_11_18_real;
        _zz_217 = img_reg_array_11_18_imag;
        _zz_218 = img_reg_array_12_18_real;
        _zz_219 = img_reg_array_12_18_imag;
        _zz_220 = img_reg_array_13_18_real;
        _zz_221 = img_reg_array_13_18_imag;
        _zz_222 = img_reg_array_14_18_real;
        _zz_223 = img_reg_array_14_18_imag;
        _zz_224 = img_reg_array_15_18_real;
        _zz_225 = img_reg_array_15_18_imag;
        _zz_226 = img_reg_array_16_18_real;
        _zz_227 = img_reg_array_16_18_imag;
        _zz_228 = img_reg_array_17_18_real;
        _zz_229 = img_reg_array_17_18_imag;
        _zz_230 = img_reg_array_18_18_real;
        _zz_231 = img_reg_array_18_18_imag;
        _zz_232 = img_reg_array_19_18_real;
        _zz_233 = img_reg_array_19_18_imag;
        _zz_234 = img_reg_array_20_18_real;
        _zz_235 = img_reg_array_20_18_imag;
        _zz_236 = img_reg_array_21_18_real;
        _zz_237 = img_reg_array_21_18_imag;
        _zz_238 = img_reg_array_22_18_real;
        _zz_239 = img_reg_array_22_18_imag;
        _zz_240 = img_reg_array_23_18_real;
        _zz_241 = img_reg_array_23_18_imag;
        _zz_242 = img_reg_array_24_18_real;
        _zz_243 = img_reg_array_24_18_imag;
        _zz_244 = img_reg_array_25_18_real;
        _zz_245 = img_reg_array_25_18_imag;
        _zz_246 = img_reg_array_26_18_real;
        _zz_247 = img_reg_array_26_18_imag;
        _zz_248 = img_reg_array_27_18_real;
        _zz_249 = img_reg_array_27_18_imag;
        _zz_250 = img_reg_array_28_18_real;
        _zz_251 = img_reg_array_28_18_imag;
        _zz_252 = img_reg_array_29_18_real;
        _zz_253 = img_reg_array_29_18_imag;
        _zz_254 = img_reg_array_30_18_real;
        _zz_255 = img_reg_array_30_18_imag;
        _zz_256 = img_reg_array_31_18_real;
        _zz_257 = img_reg_array_31_18_imag;
        _zz_258 = img_reg_array_32_18_real;
        _zz_259 = img_reg_array_32_18_imag;
        _zz_260 = img_reg_array_33_18_real;
        _zz_261 = img_reg_array_33_18_imag;
        _zz_262 = img_reg_array_34_18_real;
        _zz_263 = img_reg_array_34_18_imag;
        _zz_264 = img_reg_array_35_18_real;
        _zz_265 = img_reg_array_35_18_imag;
        _zz_266 = img_reg_array_36_18_real;
        _zz_267 = img_reg_array_36_18_imag;
        _zz_268 = img_reg_array_37_18_real;
        _zz_269 = img_reg_array_37_18_imag;
        _zz_270 = img_reg_array_38_18_real;
        _zz_271 = img_reg_array_38_18_imag;
        _zz_272 = img_reg_array_39_18_real;
        _zz_273 = img_reg_array_39_18_imag;
        _zz_274 = img_reg_array_40_18_real;
        _zz_275 = img_reg_array_40_18_imag;
        _zz_276 = img_reg_array_41_18_real;
        _zz_277 = img_reg_array_41_18_imag;
        _zz_278 = img_reg_array_42_18_real;
        _zz_279 = img_reg_array_42_18_imag;
        _zz_280 = img_reg_array_43_18_real;
        _zz_281 = img_reg_array_43_18_imag;
        _zz_282 = img_reg_array_44_18_real;
        _zz_283 = img_reg_array_44_18_imag;
        _zz_284 = img_reg_array_45_18_real;
        _zz_285 = img_reg_array_45_18_imag;
        _zz_286 = img_reg_array_46_18_real;
        _zz_287 = img_reg_array_46_18_imag;
        _zz_288 = img_reg_array_47_18_real;
        _zz_289 = img_reg_array_47_18_imag;
        _zz_290 = img_reg_array_48_18_real;
        _zz_291 = img_reg_array_48_18_imag;
        _zz_292 = img_reg_array_49_18_real;
        _zz_293 = img_reg_array_49_18_imag;
        _zz_294 = img_reg_array_50_18_real;
        _zz_295 = img_reg_array_50_18_imag;
        _zz_296 = img_reg_array_51_18_real;
        _zz_297 = img_reg_array_51_18_imag;
        _zz_298 = img_reg_array_52_18_real;
        _zz_299 = img_reg_array_52_18_imag;
        _zz_300 = img_reg_array_53_18_real;
        _zz_301 = img_reg_array_53_18_imag;
        _zz_302 = img_reg_array_54_18_real;
        _zz_303 = img_reg_array_54_18_imag;
        _zz_304 = img_reg_array_55_18_real;
        _zz_305 = img_reg_array_55_18_imag;
        _zz_306 = img_reg_array_56_18_real;
        _zz_307 = img_reg_array_56_18_imag;
        _zz_308 = img_reg_array_57_18_real;
        _zz_309 = img_reg_array_57_18_imag;
        _zz_310 = img_reg_array_58_18_real;
        _zz_311 = img_reg_array_58_18_imag;
        _zz_312 = img_reg_array_59_18_real;
        _zz_313 = img_reg_array_59_18_imag;
        _zz_314 = img_reg_array_60_18_real;
        _zz_315 = img_reg_array_60_18_imag;
        _zz_316 = img_reg_array_61_18_real;
        _zz_317 = img_reg_array_61_18_imag;
        _zz_318 = img_reg_array_62_18_real;
        _zz_319 = img_reg_array_62_18_imag;
        _zz_320 = img_reg_array_63_18_real;
        _zz_321 = img_reg_array_63_18_imag;
      end
      6'b010011 : begin
        _zz_194 = img_reg_array_0_19_real;
        _zz_195 = img_reg_array_0_19_imag;
        _zz_196 = img_reg_array_1_19_real;
        _zz_197 = img_reg_array_1_19_imag;
        _zz_198 = img_reg_array_2_19_real;
        _zz_199 = img_reg_array_2_19_imag;
        _zz_200 = img_reg_array_3_19_real;
        _zz_201 = img_reg_array_3_19_imag;
        _zz_202 = img_reg_array_4_19_real;
        _zz_203 = img_reg_array_4_19_imag;
        _zz_204 = img_reg_array_5_19_real;
        _zz_205 = img_reg_array_5_19_imag;
        _zz_206 = img_reg_array_6_19_real;
        _zz_207 = img_reg_array_6_19_imag;
        _zz_208 = img_reg_array_7_19_real;
        _zz_209 = img_reg_array_7_19_imag;
        _zz_210 = img_reg_array_8_19_real;
        _zz_211 = img_reg_array_8_19_imag;
        _zz_212 = img_reg_array_9_19_real;
        _zz_213 = img_reg_array_9_19_imag;
        _zz_214 = img_reg_array_10_19_real;
        _zz_215 = img_reg_array_10_19_imag;
        _zz_216 = img_reg_array_11_19_real;
        _zz_217 = img_reg_array_11_19_imag;
        _zz_218 = img_reg_array_12_19_real;
        _zz_219 = img_reg_array_12_19_imag;
        _zz_220 = img_reg_array_13_19_real;
        _zz_221 = img_reg_array_13_19_imag;
        _zz_222 = img_reg_array_14_19_real;
        _zz_223 = img_reg_array_14_19_imag;
        _zz_224 = img_reg_array_15_19_real;
        _zz_225 = img_reg_array_15_19_imag;
        _zz_226 = img_reg_array_16_19_real;
        _zz_227 = img_reg_array_16_19_imag;
        _zz_228 = img_reg_array_17_19_real;
        _zz_229 = img_reg_array_17_19_imag;
        _zz_230 = img_reg_array_18_19_real;
        _zz_231 = img_reg_array_18_19_imag;
        _zz_232 = img_reg_array_19_19_real;
        _zz_233 = img_reg_array_19_19_imag;
        _zz_234 = img_reg_array_20_19_real;
        _zz_235 = img_reg_array_20_19_imag;
        _zz_236 = img_reg_array_21_19_real;
        _zz_237 = img_reg_array_21_19_imag;
        _zz_238 = img_reg_array_22_19_real;
        _zz_239 = img_reg_array_22_19_imag;
        _zz_240 = img_reg_array_23_19_real;
        _zz_241 = img_reg_array_23_19_imag;
        _zz_242 = img_reg_array_24_19_real;
        _zz_243 = img_reg_array_24_19_imag;
        _zz_244 = img_reg_array_25_19_real;
        _zz_245 = img_reg_array_25_19_imag;
        _zz_246 = img_reg_array_26_19_real;
        _zz_247 = img_reg_array_26_19_imag;
        _zz_248 = img_reg_array_27_19_real;
        _zz_249 = img_reg_array_27_19_imag;
        _zz_250 = img_reg_array_28_19_real;
        _zz_251 = img_reg_array_28_19_imag;
        _zz_252 = img_reg_array_29_19_real;
        _zz_253 = img_reg_array_29_19_imag;
        _zz_254 = img_reg_array_30_19_real;
        _zz_255 = img_reg_array_30_19_imag;
        _zz_256 = img_reg_array_31_19_real;
        _zz_257 = img_reg_array_31_19_imag;
        _zz_258 = img_reg_array_32_19_real;
        _zz_259 = img_reg_array_32_19_imag;
        _zz_260 = img_reg_array_33_19_real;
        _zz_261 = img_reg_array_33_19_imag;
        _zz_262 = img_reg_array_34_19_real;
        _zz_263 = img_reg_array_34_19_imag;
        _zz_264 = img_reg_array_35_19_real;
        _zz_265 = img_reg_array_35_19_imag;
        _zz_266 = img_reg_array_36_19_real;
        _zz_267 = img_reg_array_36_19_imag;
        _zz_268 = img_reg_array_37_19_real;
        _zz_269 = img_reg_array_37_19_imag;
        _zz_270 = img_reg_array_38_19_real;
        _zz_271 = img_reg_array_38_19_imag;
        _zz_272 = img_reg_array_39_19_real;
        _zz_273 = img_reg_array_39_19_imag;
        _zz_274 = img_reg_array_40_19_real;
        _zz_275 = img_reg_array_40_19_imag;
        _zz_276 = img_reg_array_41_19_real;
        _zz_277 = img_reg_array_41_19_imag;
        _zz_278 = img_reg_array_42_19_real;
        _zz_279 = img_reg_array_42_19_imag;
        _zz_280 = img_reg_array_43_19_real;
        _zz_281 = img_reg_array_43_19_imag;
        _zz_282 = img_reg_array_44_19_real;
        _zz_283 = img_reg_array_44_19_imag;
        _zz_284 = img_reg_array_45_19_real;
        _zz_285 = img_reg_array_45_19_imag;
        _zz_286 = img_reg_array_46_19_real;
        _zz_287 = img_reg_array_46_19_imag;
        _zz_288 = img_reg_array_47_19_real;
        _zz_289 = img_reg_array_47_19_imag;
        _zz_290 = img_reg_array_48_19_real;
        _zz_291 = img_reg_array_48_19_imag;
        _zz_292 = img_reg_array_49_19_real;
        _zz_293 = img_reg_array_49_19_imag;
        _zz_294 = img_reg_array_50_19_real;
        _zz_295 = img_reg_array_50_19_imag;
        _zz_296 = img_reg_array_51_19_real;
        _zz_297 = img_reg_array_51_19_imag;
        _zz_298 = img_reg_array_52_19_real;
        _zz_299 = img_reg_array_52_19_imag;
        _zz_300 = img_reg_array_53_19_real;
        _zz_301 = img_reg_array_53_19_imag;
        _zz_302 = img_reg_array_54_19_real;
        _zz_303 = img_reg_array_54_19_imag;
        _zz_304 = img_reg_array_55_19_real;
        _zz_305 = img_reg_array_55_19_imag;
        _zz_306 = img_reg_array_56_19_real;
        _zz_307 = img_reg_array_56_19_imag;
        _zz_308 = img_reg_array_57_19_real;
        _zz_309 = img_reg_array_57_19_imag;
        _zz_310 = img_reg_array_58_19_real;
        _zz_311 = img_reg_array_58_19_imag;
        _zz_312 = img_reg_array_59_19_real;
        _zz_313 = img_reg_array_59_19_imag;
        _zz_314 = img_reg_array_60_19_real;
        _zz_315 = img_reg_array_60_19_imag;
        _zz_316 = img_reg_array_61_19_real;
        _zz_317 = img_reg_array_61_19_imag;
        _zz_318 = img_reg_array_62_19_real;
        _zz_319 = img_reg_array_62_19_imag;
        _zz_320 = img_reg_array_63_19_real;
        _zz_321 = img_reg_array_63_19_imag;
      end
      6'b010100 : begin
        _zz_194 = img_reg_array_0_20_real;
        _zz_195 = img_reg_array_0_20_imag;
        _zz_196 = img_reg_array_1_20_real;
        _zz_197 = img_reg_array_1_20_imag;
        _zz_198 = img_reg_array_2_20_real;
        _zz_199 = img_reg_array_2_20_imag;
        _zz_200 = img_reg_array_3_20_real;
        _zz_201 = img_reg_array_3_20_imag;
        _zz_202 = img_reg_array_4_20_real;
        _zz_203 = img_reg_array_4_20_imag;
        _zz_204 = img_reg_array_5_20_real;
        _zz_205 = img_reg_array_5_20_imag;
        _zz_206 = img_reg_array_6_20_real;
        _zz_207 = img_reg_array_6_20_imag;
        _zz_208 = img_reg_array_7_20_real;
        _zz_209 = img_reg_array_7_20_imag;
        _zz_210 = img_reg_array_8_20_real;
        _zz_211 = img_reg_array_8_20_imag;
        _zz_212 = img_reg_array_9_20_real;
        _zz_213 = img_reg_array_9_20_imag;
        _zz_214 = img_reg_array_10_20_real;
        _zz_215 = img_reg_array_10_20_imag;
        _zz_216 = img_reg_array_11_20_real;
        _zz_217 = img_reg_array_11_20_imag;
        _zz_218 = img_reg_array_12_20_real;
        _zz_219 = img_reg_array_12_20_imag;
        _zz_220 = img_reg_array_13_20_real;
        _zz_221 = img_reg_array_13_20_imag;
        _zz_222 = img_reg_array_14_20_real;
        _zz_223 = img_reg_array_14_20_imag;
        _zz_224 = img_reg_array_15_20_real;
        _zz_225 = img_reg_array_15_20_imag;
        _zz_226 = img_reg_array_16_20_real;
        _zz_227 = img_reg_array_16_20_imag;
        _zz_228 = img_reg_array_17_20_real;
        _zz_229 = img_reg_array_17_20_imag;
        _zz_230 = img_reg_array_18_20_real;
        _zz_231 = img_reg_array_18_20_imag;
        _zz_232 = img_reg_array_19_20_real;
        _zz_233 = img_reg_array_19_20_imag;
        _zz_234 = img_reg_array_20_20_real;
        _zz_235 = img_reg_array_20_20_imag;
        _zz_236 = img_reg_array_21_20_real;
        _zz_237 = img_reg_array_21_20_imag;
        _zz_238 = img_reg_array_22_20_real;
        _zz_239 = img_reg_array_22_20_imag;
        _zz_240 = img_reg_array_23_20_real;
        _zz_241 = img_reg_array_23_20_imag;
        _zz_242 = img_reg_array_24_20_real;
        _zz_243 = img_reg_array_24_20_imag;
        _zz_244 = img_reg_array_25_20_real;
        _zz_245 = img_reg_array_25_20_imag;
        _zz_246 = img_reg_array_26_20_real;
        _zz_247 = img_reg_array_26_20_imag;
        _zz_248 = img_reg_array_27_20_real;
        _zz_249 = img_reg_array_27_20_imag;
        _zz_250 = img_reg_array_28_20_real;
        _zz_251 = img_reg_array_28_20_imag;
        _zz_252 = img_reg_array_29_20_real;
        _zz_253 = img_reg_array_29_20_imag;
        _zz_254 = img_reg_array_30_20_real;
        _zz_255 = img_reg_array_30_20_imag;
        _zz_256 = img_reg_array_31_20_real;
        _zz_257 = img_reg_array_31_20_imag;
        _zz_258 = img_reg_array_32_20_real;
        _zz_259 = img_reg_array_32_20_imag;
        _zz_260 = img_reg_array_33_20_real;
        _zz_261 = img_reg_array_33_20_imag;
        _zz_262 = img_reg_array_34_20_real;
        _zz_263 = img_reg_array_34_20_imag;
        _zz_264 = img_reg_array_35_20_real;
        _zz_265 = img_reg_array_35_20_imag;
        _zz_266 = img_reg_array_36_20_real;
        _zz_267 = img_reg_array_36_20_imag;
        _zz_268 = img_reg_array_37_20_real;
        _zz_269 = img_reg_array_37_20_imag;
        _zz_270 = img_reg_array_38_20_real;
        _zz_271 = img_reg_array_38_20_imag;
        _zz_272 = img_reg_array_39_20_real;
        _zz_273 = img_reg_array_39_20_imag;
        _zz_274 = img_reg_array_40_20_real;
        _zz_275 = img_reg_array_40_20_imag;
        _zz_276 = img_reg_array_41_20_real;
        _zz_277 = img_reg_array_41_20_imag;
        _zz_278 = img_reg_array_42_20_real;
        _zz_279 = img_reg_array_42_20_imag;
        _zz_280 = img_reg_array_43_20_real;
        _zz_281 = img_reg_array_43_20_imag;
        _zz_282 = img_reg_array_44_20_real;
        _zz_283 = img_reg_array_44_20_imag;
        _zz_284 = img_reg_array_45_20_real;
        _zz_285 = img_reg_array_45_20_imag;
        _zz_286 = img_reg_array_46_20_real;
        _zz_287 = img_reg_array_46_20_imag;
        _zz_288 = img_reg_array_47_20_real;
        _zz_289 = img_reg_array_47_20_imag;
        _zz_290 = img_reg_array_48_20_real;
        _zz_291 = img_reg_array_48_20_imag;
        _zz_292 = img_reg_array_49_20_real;
        _zz_293 = img_reg_array_49_20_imag;
        _zz_294 = img_reg_array_50_20_real;
        _zz_295 = img_reg_array_50_20_imag;
        _zz_296 = img_reg_array_51_20_real;
        _zz_297 = img_reg_array_51_20_imag;
        _zz_298 = img_reg_array_52_20_real;
        _zz_299 = img_reg_array_52_20_imag;
        _zz_300 = img_reg_array_53_20_real;
        _zz_301 = img_reg_array_53_20_imag;
        _zz_302 = img_reg_array_54_20_real;
        _zz_303 = img_reg_array_54_20_imag;
        _zz_304 = img_reg_array_55_20_real;
        _zz_305 = img_reg_array_55_20_imag;
        _zz_306 = img_reg_array_56_20_real;
        _zz_307 = img_reg_array_56_20_imag;
        _zz_308 = img_reg_array_57_20_real;
        _zz_309 = img_reg_array_57_20_imag;
        _zz_310 = img_reg_array_58_20_real;
        _zz_311 = img_reg_array_58_20_imag;
        _zz_312 = img_reg_array_59_20_real;
        _zz_313 = img_reg_array_59_20_imag;
        _zz_314 = img_reg_array_60_20_real;
        _zz_315 = img_reg_array_60_20_imag;
        _zz_316 = img_reg_array_61_20_real;
        _zz_317 = img_reg_array_61_20_imag;
        _zz_318 = img_reg_array_62_20_real;
        _zz_319 = img_reg_array_62_20_imag;
        _zz_320 = img_reg_array_63_20_real;
        _zz_321 = img_reg_array_63_20_imag;
      end
      6'b010101 : begin
        _zz_194 = img_reg_array_0_21_real;
        _zz_195 = img_reg_array_0_21_imag;
        _zz_196 = img_reg_array_1_21_real;
        _zz_197 = img_reg_array_1_21_imag;
        _zz_198 = img_reg_array_2_21_real;
        _zz_199 = img_reg_array_2_21_imag;
        _zz_200 = img_reg_array_3_21_real;
        _zz_201 = img_reg_array_3_21_imag;
        _zz_202 = img_reg_array_4_21_real;
        _zz_203 = img_reg_array_4_21_imag;
        _zz_204 = img_reg_array_5_21_real;
        _zz_205 = img_reg_array_5_21_imag;
        _zz_206 = img_reg_array_6_21_real;
        _zz_207 = img_reg_array_6_21_imag;
        _zz_208 = img_reg_array_7_21_real;
        _zz_209 = img_reg_array_7_21_imag;
        _zz_210 = img_reg_array_8_21_real;
        _zz_211 = img_reg_array_8_21_imag;
        _zz_212 = img_reg_array_9_21_real;
        _zz_213 = img_reg_array_9_21_imag;
        _zz_214 = img_reg_array_10_21_real;
        _zz_215 = img_reg_array_10_21_imag;
        _zz_216 = img_reg_array_11_21_real;
        _zz_217 = img_reg_array_11_21_imag;
        _zz_218 = img_reg_array_12_21_real;
        _zz_219 = img_reg_array_12_21_imag;
        _zz_220 = img_reg_array_13_21_real;
        _zz_221 = img_reg_array_13_21_imag;
        _zz_222 = img_reg_array_14_21_real;
        _zz_223 = img_reg_array_14_21_imag;
        _zz_224 = img_reg_array_15_21_real;
        _zz_225 = img_reg_array_15_21_imag;
        _zz_226 = img_reg_array_16_21_real;
        _zz_227 = img_reg_array_16_21_imag;
        _zz_228 = img_reg_array_17_21_real;
        _zz_229 = img_reg_array_17_21_imag;
        _zz_230 = img_reg_array_18_21_real;
        _zz_231 = img_reg_array_18_21_imag;
        _zz_232 = img_reg_array_19_21_real;
        _zz_233 = img_reg_array_19_21_imag;
        _zz_234 = img_reg_array_20_21_real;
        _zz_235 = img_reg_array_20_21_imag;
        _zz_236 = img_reg_array_21_21_real;
        _zz_237 = img_reg_array_21_21_imag;
        _zz_238 = img_reg_array_22_21_real;
        _zz_239 = img_reg_array_22_21_imag;
        _zz_240 = img_reg_array_23_21_real;
        _zz_241 = img_reg_array_23_21_imag;
        _zz_242 = img_reg_array_24_21_real;
        _zz_243 = img_reg_array_24_21_imag;
        _zz_244 = img_reg_array_25_21_real;
        _zz_245 = img_reg_array_25_21_imag;
        _zz_246 = img_reg_array_26_21_real;
        _zz_247 = img_reg_array_26_21_imag;
        _zz_248 = img_reg_array_27_21_real;
        _zz_249 = img_reg_array_27_21_imag;
        _zz_250 = img_reg_array_28_21_real;
        _zz_251 = img_reg_array_28_21_imag;
        _zz_252 = img_reg_array_29_21_real;
        _zz_253 = img_reg_array_29_21_imag;
        _zz_254 = img_reg_array_30_21_real;
        _zz_255 = img_reg_array_30_21_imag;
        _zz_256 = img_reg_array_31_21_real;
        _zz_257 = img_reg_array_31_21_imag;
        _zz_258 = img_reg_array_32_21_real;
        _zz_259 = img_reg_array_32_21_imag;
        _zz_260 = img_reg_array_33_21_real;
        _zz_261 = img_reg_array_33_21_imag;
        _zz_262 = img_reg_array_34_21_real;
        _zz_263 = img_reg_array_34_21_imag;
        _zz_264 = img_reg_array_35_21_real;
        _zz_265 = img_reg_array_35_21_imag;
        _zz_266 = img_reg_array_36_21_real;
        _zz_267 = img_reg_array_36_21_imag;
        _zz_268 = img_reg_array_37_21_real;
        _zz_269 = img_reg_array_37_21_imag;
        _zz_270 = img_reg_array_38_21_real;
        _zz_271 = img_reg_array_38_21_imag;
        _zz_272 = img_reg_array_39_21_real;
        _zz_273 = img_reg_array_39_21_imag;
        _zz_274 = img_reg_array_40_21_real;
        _zz_275 = img_reg_array_40_21_imag;
        _zz_276 = img_reg_array_41_21_real;
        _zz_277 = img_reg_array_41_21_imag;
        _zz_278 = img_reg_array_42_21_real;
        _zz_279 = img_reg_array_42_21_imag;
        _zz_280 = img_reg_array_43_21_real;
        _zz_281 = img_reg_array_43_21_imag;
        _zz_282 = img_reg_array_44_21_real;
        _zz_283 = img_reg_array_44_21_imag;
        _zz_284 = img_reg_array_45_21_real;
        _zz_285 = img_reg_array_45_21_imag;
        _zz_286 = img_reg_array_46_21_real;
        _zz_287 = img_reg_array_46_21_imag;
        _zz_288 = img_reg_array_47_21_real;
        _zz_289 = img_reg_array_47_21_imag;
        _zz_290 = img_reg_array_48_21_real;
        _zz_291 = img_reg_array_48_21_imag;
        _zz_292 = img_reg_array_49_21_real;
        _zz_293 = img_reg_array_49_21_imag;
        _zz_294 = img_reg_array_50_21_real;
        _zz_295 = img_reg_array_50_21_imag;
        _zz_296 = img_reg_array_51_21_real;
        _zz_297 = img_reg_array_51_21_imag;
        _zz_298 = img_reg_array_52_21_real;
        _zz_299 = img_reg_array_52_21_imag;
        _zz_300 = img_reg_array_53_21_real;
        _zz_301 = img_reg_array_53_21_imag;
        _zz_302 = img_reg_array_54_21_real;
        _zz_303 = img_reg_array_54_21_imag;
        _zz_304 = img_reg_array_55_21_real;
        _zz_305 = img_reg_array_55_21_imag;
        _zz_306 = img_reg_array_56_21_real;
        _zz_307 = img_reg_array_56_21_imag;
        _zz_308 = img_reg_array_57_21_real;
        _zz_309 = img_reg_array_57_21_imag;
        _zz_310 = img_reg_array_58_21_real;
        _zz_311 = img_reg_array_58_21_imag;
        _zz_312 = img_reg_array_59_21_real;
        _zz_313 = img_reg_array_59_21_imag;
        _zz_314 = img_reg_array_60_21_real;
        _zz_315 = img_reg_array_60_21_imag;
        _zz_316 = img_reg_array_61_21_real;
        _zz_317 = img_reg_array_61_21_imag;
        _zz_318 = img_reg_array_62_21_real;
        _zz_319 = img_reg_array_62_21_imag;
        _zz_320 = img_reg_array_63_21_real;
        _zz_321 = img_reg_array_63_21_imag;
      end
      6'b010110 : begin
        _zz_194 = img_reg_array_0_22_real;
        _zz_195 = img_reg_array_0_22_imag;
        _zz_196 = img_reg_array_1_22_real;
        _zz_197 = img_reg_array_1_22_imag;
        _zz_198 = img_reg_array_2_22_real;
        _zz_199 = img_reg_array_2_22_imag;
        _zz_200 = img_reg_array_3_22_real;
        _zz_201 = img_reg_array_3_22_imag;
        _zz_202 = img_reg_array_4_22_real;
        _zz_203 = img_reg_array_4_22_imag;
        _zz_204 = img_reg_array_5_22_real;
        _zz_205 = img_reg_array_5_22_imag;
        _zz_206 = img_reg_array_6_22_real;
        _zz_207 = img_reg_array_6_22_imag;
        _zz_208 = img_reg_array_7_22_real;
        _zz_209 = img_reg_array_7_22_imag;
        _zz_210 = img_reg_array_8_22_real;
        _zz_211 = img_reg_array_8_22_imag;
        _zz_212 = img_reg_array_9_22_real;
        _zz_213 = img_reg_array_9_22_imag;
        _zz_214 = img_reg_array_10_22_real;
        _zz_215 = img_reg_array_10_22_imag;
        _zz_216 = img_reg_array_11_22_real;
        _zz_217 = img_reg_array_11_22_imag;
        _zz_218 = img_reg_array_12_22_real;
        _zz_219 = img_reg_array_12_22_imag;
        _zz_220 = img_reg_array_13_22_real;
        _zz_221 = img_reg_array_13_22_imag;
        _zz_222 = img_reg_array_14_22_real;
        _zz_223 = img_reg_array_14_22_imag;
        _zz_224 = img_reg_array_15_22_real;
        _zz_225 = img_reg_array_15_22_imag;
        _zz_226 = img_reg_array_16_22_real;
        _zz_227 = img_reg_array_16_22_imag;
        _zz_228 = img_reg_array_17_22_real;
        _zz_229 = img_reg_array_17_22_imag;
        _zz_230 = img_reg_array_18_22_real;
        _zz_231 = img_reg_array_18_22_imag;
        _zz_232 = img_reg_array_19_22_real;
        _zz_233 = img_reg_array_19_22_imag;
        _zz_234 = img_reg_array_20_22_real;
        _zz_235 = img_reg_array_20_22_imag;
        _zz_236 = img_reg_array_21_22_real;
        _zz_237 = img_reg_array_21_22_imag;
        _zz_238 = img_reg_array_22_22_real;
        _zz_239 = img_reg_array_22_22_imag;
        _zz_240 = img_reg_array_23_22_real;
        _zz_241 = img_reg_array_23_22_imag;
        _zz_242 = img_reg_array_24_22_real;
        _zz_243 = img_reg_array_24_22_imag;
        _zz_244 = img_reg_array_25_22_real;
        _zz_245 = img_reg_array_25_22_imag;
        _zz_246 = img_reg_array_26_22_real;
        _zz_247 = img_reg_array_26_22_imag;
        _zz_248 = img_reg_array_27_22_real;
        _zz_249 = img_reg_array_27_22_imag;
        _zz_250 = img_reg_array_28_22_real;
        _zz_251 = img_reg_array_28_22_imag;
        _zz_252 = img_reg_array_29_22_real;
        _zz_253 = img_reg_array_29_22_imag;
        _zz_254 = img_reg_array_30_22_real;
        _zz_255 = img_reg_array_30_22_imag;
        _zz_256 = img_reg_array_31_22_real;
        _zz_257 = img_reg_array_31_22_imag;
        _zz_258 = img_reg_array_32_22_real;
        _zz_259 = img_reg_array_32_22_imag;
        _zz_260 = img_reg_array_33_22_real;
        _zz_261 = img_reg_array_33_22_imag;
        _zz_262 = img_reg_array_34_22_real;
        _zz_263 = img_reg_array_34_22_imag;
        _zz_264 = img_reg_array_35_22_real;
        _zz_265 = img_reg_array_35_22_imag;
        _zz_266 = img_reg_array_36_22_real;
        _zz_267 = img_reg_array_36_22_imag;
        _zz_268 = img_reg_array_37_22_real;
        _zz_269 = img_reg_array_37_22_imag;
        _zz_270 = img_reg_array_38_22_real;
        _zz_271 = img_reg_array_38_22_imag;
        _zz_272 = img_reg_array_39_22_real;
        _zz_273 = img_reg_array_39_22_imag;
        _zz_274 = img_reg_array_40_22_real;
        _zz_275 = img_reg_array_40_22_imag;
        _zz_276 = img_reg_array_41_22_real;
        _zz_277 = img_reg_array_41_22_imag;
        _zz_278 = img_reg_array_42_22_real;
        _zz_279 = img_reg_array_42_22_imag;
        _zz_280 = img_reg_array_43_22_real;
        _zz_281 = img_reg_array_43_22_imag;
        _zz_282 = img_reg_array_44_22_real;
        _zz_283 = img_reg_array_44_22_imag;
        _zz_284 = img_reg_array_45_22_real;
        _zz_285 = img_reg_array_45_22_imag;
        _zz_286 = img_reg_array_46_22_real;
        _zz_287 = img_reg_array_46_22_imag;
        _zz_288 = img_reg_array_47_22_real;
        _zz_289 = img_reg_array_47_22_imag;
        _zz_290 = img_reg_array_48_22_real;
        _zz_291 = img_reg_array_48_22_imag;
        _zz_292 = img_reg_array_49_22_real;
        _zz_293 = img_reg_array_49_22_imag;
        _zz_294 = img_reg_array_50_22_real;
        _zz_295 = img_reg_array_50_22_imag;
        _zz_296 = img_reg_array_51_22_real;
        _zz_297 = img_reg_array_51_22_imag;
        _zz_298 = img_reg_array_52_22_real;
        _zz_299 = img_reg_array_52_22_imag;
        _zz_300 = img_reg_array_53_22_real;
        _zz_301 = img_reg_array_53_22_imag;
        _zz_302 = img_reg_array_54_22_real;
        _zz_303 = img_reg_array_54_22_imag;
        _zz_304 = img_reg_array_55_22_real;
        _zz_305 = img_reg_array_55_22_imag;
        _zz_306 = img_reg_array_56_22_real;
        _zz_307 = img_reg_array_56_22_imag;
        _zz_308 = img_reg_array_57_22_real;
        _zz_309 = img_reg_array_57_22_imag;
        _zz_310 = img_reg_array_58_22_real;
        _zz_311 = img_reg_array_58_22_imag;
        _zz_312 = img_reg_array_59_22_real;
        _zz_313 = img_reg_array_59_22_imag;
        _zz_314 = img_reg_array_60_22_real;
        _zz_315 = img_reg_array_60_22_imag;
        _zz_316 = img_reg_array_61_22_real;
        _zz_317 = img_reg_array_61_22_imag;
        _zz_318 = img_reg_array_62_22_real;
        _zz_319 = img_reg_array_62_22_imag;
        _zz_320 = img_reg_array_63_22_real;
        _zz_321 = img_reg_array_63_22_imag;
      end
      6'b010111 : begin
        _zz_194 = img_reg_array_0_23_real;
        _zz_195 = img_reg_array_0_23_imag;
        _zz_196 = img_reg_array_1_23_real;
        _zz_197 = img_reg_array_1_23_imag;
        _zz_198 = img_reg_array_2_23_real;
        _zz_199 = img_reg_array_2_23_imag;
        _zz_200 = img_reg_array_3_23_real;
        _zz_201 = img_reg_array_3_23_imag;
        _zz_202 = img_reg_array_4_23_real;
        _zz_203 = img_reg_array_4_23_imag;
        _zz_204 = img_reg_array_5_23_real;
        _zz_205 = img_reg_array_5_23_imag;
        _zz_206 = img_reg_array_6_23_real;
        _zz_207 = img_reg_array_6_23_imag;
        _zz_208 = img_reg_array_7_23_real;
        _zz_209 = img_reg_array_7_23_imag;
        _zz_210 = img_reg_array_8_23_real;
        _zz_211 = img_reg_array_8_23_imag;
        _zz_212 = img_reg_array_9_23_real;
        _zz_213 = img_reg_array_9_23_imag;
        _zz_214 = img_reg_array_10_23_real;
        _zz_215 = img_reg_array_10_23_imag;
        _zz_216 = img_reg_array_11_23_real;
        _zz_217 = img_reg_array_11_23_imag;
        _zz_218 = img_reg_array_12_23_real;
        _zz_219 = img_reg_array_12_23_imag;
        _zz_220 = img_reg_array_13_23_real;
        _zz_221 = img_reg_array_13_23_imag;
        _zz_222 = img_reg_array_14_23_real;
        _zz_223 = img_reg_array_14_23_imag;
        _zz_224 = img_reg_array_15_23_real;
        _zz_225 = img_reg_array_15_23_imag;
        _zz_226 = img_reg_array_16_23_real;
        _zz_227 = img_reg_array_16_23_imag;
        _zz_228 = img_reg_array_17_23_real;
        _zz_229 = img_reg_array_17_23_imag;
        _zz_230 = img_reg_array_18_23_real;
        _zz_231 = img_reg_array_18_23_imag;
        _zz_232 = img_reg_array_19_23_real;
        _zz_233 = img_reg_array_19_23_imag;
        _zz_234 = img_reg_array_20_23_real;
        _zz_235 = img_reg_array_20_23_imag;
        _zz_236 = img_reg_array_21_23_real;
        _zz_237 = img_reg_array_21_23_imag;
        _zz_238 = img_reg_array_22_23_real;
        _zz_239 = img_reg_array_22_23_imag;
        _zz_240 = img_reg_array_23_23_real;
        _zz_241 = img_reg_array_23_23_imag;
        _zz_242 = img_reg_array_24_23_real;
        _zz_243 = img_reg_array_24_23_imag;
        _zz_244 = img_reg_array_25_23_real;
        _zz_245 = img_reg_array_25_23_imag;
        _zz_246 = img_reg_array_26_23_real;
        _zz_247 = img_reg_array_26_23_imag;
        _zz_248 = img_reg_array_27_23_real;
        _zz_249 = img_reg_array_27_23_imag;
        _zz_250 = img_reg_array_28_23_real;
        _zz_251 = img_reg_array_28_23_imag;
        _zz_252 = img_reg_array_29_23_real;
        _zz_253 = img_reg_array_29_23_imag;
        _zz_254 = img_reg_array_30_23_real;
        _zz_255 = img_reg_array_30_23_imag;
        _zz_256 = img_reg_array_31_23_real;
        _zz_257 = img_reg_array_31_23_imag;
        _zz_258 = img_reg_array_32_23_real;
        _zz_259 = img_reg_array_32_23_imag;
        _zz_260 = img_reg_array_33_23_real;
        _zz_261 = img_reg_array_33_23_imag;
        _zz_262 = img_reg_array_34_23_real;
        _zz_263 = img_reg_array_34_23_imag;
        _zz_264 = img_reg_array_35_23_real;
        _zz_265 = img_reg_array_35_23_imag;
        _zz_266 = img_reg_array_36_23_real;
        _zz_267 = img_reg_array_36_23_imag;
        _zz_268 = img_reg_array_37_23_real;
        _zz_269 = img_reg_array_37_23_imag;
        _zz_270 = img_reg_array_38_23_real;
        _zz_271 = img_reg_array_38_23_imag;
        _zz_272 = img_reg_array_39_23_real;
        _zz_273 = img_reg_array_39_23_imag;
        _zz_274 = img_reg_array_40_23_real;
        _zz_275 = img_reg_array_40_23_imag;
        _zz_276 = img_reg_array_41_23_real;
        _zz_277 = img_reg_array_41_23_imag;
        _zz_278 = img_reg_array_42_23_real;
        _zz_279 = img_reg_array_42_23_imag;
        _zz_280 = img_reg_array_43_23_real;
        _zz_281 = img_reg_array_43_23_imag;
        _zz_282 = img_reg_array_44_23_real;
        _zz_283 = img_reg_array_44_23_imag;
        _zz_284 = img_reg_array_45_23_real;
        _zz_285 = img_reg_array_45_23_imag;
        _zz_286 = img_reg_array_46_23_real;
        _zz_287 = img_reg_array_46_23_imag;
        _zz_288 = img_reg_array_47_23_real;
        _zz_289 = img_reg_array_47_23_imag;
        _zz_290 = img_reg_array_48_23_real;
        _zz_291 = img_reg_array_48_23_imag;
        _zz_292 = img_reg_array_49_23_real;
        _zz_293 = img_reg_array_49_23_imag;
        _zz_294 = img_reg_array_50_23_real;
        _zz_295 = img_reg_array_50_23_imag;
        _zz_296 = img_reg_array_51_23_real;
        _zz_297 = img_reg_array_51_23_imag;
        _zz_298 = img_reg_array_52_23_real;
        _zz_299 = img_reg_array_52_23_imag;
        _zz_300 = img_reg_array_53_23_real;
        _zz_301 = img_reg_array_53_23_imag;
        _zz_302 = img_reg_array_54_23_real;
        _zz_303 = img_reg_array_54_23_imag;
        _zz_304 = img_reg_array_55_23_real;
        _zz_305 = img_reg_array_55_23_imag;
        _zz_306 = img_reg_array_56_23_real;
        _zz_307 = img_reg_array_56_23_imag;
        _zz_308 = img_reg_array_57_23_real;
        _zz_309 = img_reg_array_57_23_imag;
        _zz_310 = img_reg_array_58_23_real;
        _zz_311 = img_reg_array_58_23_imag;
        _zz_312 = img_reg_array_59_23_real;
        _zz_313 = img_reg_array_59_23_imag;
        _zz_314 = img_reg_array_60_23_real;
        _zz_315 = img_reg_array_60_23_imag;
        _zz_316 = img_reg_array_61_23_real;
        _zz_317 = img_reg_array_61_23_imag;
        _zz_318 = img_reg_array_62_23_real;
        _zz_319 = img_reg_array_62_23_imag;
        _zz_320 = img_reg_array_63_23_real;
        _zz_321 = img_reg_array_63_23_imag;
      end
      6'b011000 : begin
        _zz_194 = img_reg_array_0_24_real;
        _zz_195 = img_reg_array_0_24_imag;
        _zz_196 = img_reg_array_1_24_real;
        _zz_197 = img_reg_array_1_24_imag;
        _zz_198 = img_reg_array_2_24_real;
        _zz_199 = img_reg_array_2_24_imag;
        _zz_200 = img_reg_array_3_24_real;
        _zz_201 = img_reg_array_3_24_imag;
        _zz_202 = img_reg_array_4_24_real;
        _zz_203 = img_reg_array_4_24_imag;
        _zz_204 = img_reg_array_5_24_real;
        _zz_205 = img_reg_array_5_24_imag;
        _zz_206 = img_reg_array_6_24_real;
        _zz_207 = img_reg_array_6_24_imag;
        _zz_208 = img_reg_array_7_24_real;
        _zz_209 = img_reg_array_7_24_imag;
        _zz_210 = img_reg_array_8_24_real;
        _zz_211 = img_reg_array_8_24_imag;
        _zz_212 = img_reg_array_9_24_real;
        _zz_213 = img_reg_array_9_24_imag;
        _zz_214 = img_reg_array_10_24_real;
        _zz_215 = img_reg_array_10_24_imag;
        _zz_216 = img_reg_array_11_24_real;
        _zz_217 = img_reg_array_11_24_imag;
        _zz_218 = img_reg_array_12_24_real;
        _zz_219 = img_reg_array_12_24_imag;
        _zz_220 = img_reg_array_13_24_real;
        _zz_221 = img_reg_array_13_24_imag;
        _zz_222 = img_reg_array_14_24_real;
        _zz_223 = img_reg_array_14_24_imag;
        _zz_224 = img_reg_array_15_24_real;
        _zz_225 = img_reg_array_15_24_imag;
        _zz_226 = img_reg_array_16_24_real;
        _zz_227 = img_reg_array_16_24_imag;
        _zz_228 = img_reg_array_17_24_real;
        _zz_229 = img_reg_array_17_24_imag;
        _zz_230 = img_reg_array_18_24_real;
        _zz_231 = img_reg_array_18_24_imag;
        _zz_232 = img_reg_array_19_24_real;
        _zz_233 = img_reg_array_19_24_imag;
        _zz_234 = img_reg_array_20_24_real;
        _zz_235 = img_reg_array_20_24_imag;
        _zz_236 = img_reg_array_21_24_real;
        _zz_237 = img_reg_array_21_24_imag;
        _zz_238 = img_reg_array_22_24_real;
        _zz_239 = img_reg_array_22_24_imag;
        _zz_240 = img_reg_array_23_24_real;
        _zz_241 = img_reg_array_23_24_imag;
        _zz_242 = img_reg_array_24_24_real;
        _zz_243 = img_reg_array_24_24_imag;
        _zz_244 = img_reg_array_25_24_real;
        _zz_245 = img_reg_array_25_24_imag;
        _zz_246 = img_reg_array_26_24_real;
        _zz_247 = img_reg_array_26_24_imag;
        _zz_248 = img_reg_array_27_24_real;
        _zz_249 = img_reg_array_27_24_imag;
        _zz_250 = img_reg_array_28_24_real;
        _zz_251 = img_reg_array_28_24_imag;
        _zz_252 = img_reg_array_29_24_real;
        _zz_253 = img_reg_array_29_24_imag;
        _zz_254 = img_reg_array_30_24_real;
        _zz_255 = img_reg_array_30_24_imag;
        _zz_256 = img_reg_array_31_24_real;
        _zz_257 = img_reg_array_31_24_imag;
        _zz_258 = img_reg_array_32_24_real;
        _zz_259 = img_reg_array_32_24_imag;
        _zz_260 = img_reg_array_33_24_real;
        _zz_261 = img_reg_array_33_24_imag;
        _zz_262 = img_reg_array_34_24_real;
        _zz_263 = img_reg_array_34_24_imag;
        _zz_264 = img_reg_array_35_24_real;
        _zz_265 = img_reg_array_35_24_imag;
        _zz_266 = img_reg_array_36_24_real;
        _zz_267 = img_reg_array_36_24_imag;
        _zz_268 = img_reg_array_37_24_real;
        _zz_269 = img_reg_array_37_24_imag;
        _zz_270 = img_reg_array_38_24_real;
        _zz_271 = img_reg_array_38_24_imag;
        _zz_272 = img_reg_array_39_24_real;
        _zz_273 = img_reg_array_39_24_imag;
        _zz_274 = img_reg_array_40_24_real;
        _zz_275 = img_reg_array_40_24_imag;
        _zz_276 = img_reg_array_41_24_real;
        _zz_277 = img_reg_array_41_24_imag;
        _zz_278 = img_reg_array_42_24_real;
        _zz_279 = img_reg_array_42_24_imag;
        _zz_280 = img_reg_array_43_24_real;
        _zz_281 = img_reg_array_43_24_imag;
        _zz_282 = img_reg_array_44_24_real;
        _zz_283 = img_reg_array_44_24_imag;
        _zz_284 = img_reg_array_45_24_real;
        _zz_285 = img_reg_array_45_24_imag;
        _zz_286 = img_reg_array_46_24_real;
        _zz_287 = img_reg_array_46_24_imag;
        _zz_288 = img_reg_array_47_24_real;
        _zz_289 = img_reg_array_47_24_imag;
        _zz_290 = img_reg_array_48_24_real;
        _zz_291 = img_reg_array_48_24_imag;
        _zz_292 = img_reg_array_49_24_real;
        _zz_293 = img_reg_array_49_24_imag;
        _zz_294 = img_reg_array_50_24_real;
        _zz_295 = img_reg_array_50_24_imag;
        _zz_296 = img_reg_array_51_24_real;
        _zz_297 = img_reg_array_51_24_imag;
        _zz_298 = img_reg_array_52_24_real;
        _zz_299 = img_reg_array_52_24_imag;
        _zz_300 = img_reg_array_53_24_real;
        _zz_301 = img_reg_array_53_24_imag;
        _zz_302 = img_reg_array_54_24_real;
        _zz_303 = img_reg_array_54_24_imag;
        _zz_304 = img_reg_array_55_24_real;
        _zz_305 = img_reg_array_55_24_imag;
        _zz_306 = img_reg_array_56_24_real;
        _zz_307 = img_reg_array_56_24_imag;
        _zz_308 = img_reg_array_57_24_real;
        _zz_309 = img_reg_array_57_24_imag;
        _zz_310 = img_reg_array_58_24_real;
        _zz_311 = img_reg_array_58_24_imag;
        _zz_312 = img_reg_array_59_24_real;
        _zz_313 = img_reg_array_59_24_imag;
        _zz_314 = img_reg_array_60_24_real;
        _zz_315 = img_reg_array_60_24_imag;
        _zz_316 = img_reg_array_61_24_real;
        _zz_317 = img_reg_array_61_24_imag;
        _zz_318 = img_reg_array_62_24_real;
        _zz_319 = img_reg_array_62_24_imag;
        _zz_320 = img_reg_array_63_24_real;
        _zz_321 = img_reg_array_63_24_imag;
      end
      6'b011001 : begin
        _zz_194 = img_reg_array_0_25_real;
        _zz_195 = img_reg_array_0_25_imag;
        _zz_196 = img_reg_array_1_25_real;
        _zz_197 = img_reg_array_1_25_imag;
        _zz_198 = img_reg_array_2_25_real;
        _zz_199 = img_reg_array_2_25_imag;
        _zz_200 = img_reg_array_3_25_real;
        _zz_201 = img_reg_array_3_25_imag;
        _zz_202 = img_reg_array_4_25_real;
        _zz_203 = img_reg_array_4_25_imag;
        _zz_204 = img_reg_array_5_25_real;
        _zz_205 = img_reg_array_5_25_imag;
        _zz_206 = img_reg_array_6_25_real;
        _zz_207 = img_reg_array_6_25_imag;
        _zz_208 = img_reg_array_7_25_real;
        _zz_209 = img_reg_array_7_25_imag;
        _zz_210 = img_reg_array_8_25_real;
        _zz_211 = img_reg_array_8_25_imag;
        _zz_212 = img_reg_array_9_25_real;
        _zz_213 = img_reg_array_9_25_imag;
        _zz_214 = img_reg_array_10_25_real;
        _zz_215 = img_reg_array_10_25_imag;
        _zz_216 = img_reg_array_11_25_real;
        _zz_217 = img_reg_array_11_25_imag;
        _zz_218 = img_reg_array_12_25_real;
        _zz_219 = img_reg_array_12_25_imag;
        _zz_220 = img_reg_array_13_25_real;
        _zz_221 = img_reg_array_13_25_imag;
        _zz_222 = img_reg_array_14_25_real;
        _zz_223 = img_reg_array_14_25_imag;
        _zz_224 = img_reg_array_15_25_real;
        _zz_225 = img_reg_array_15_25_imag;
        _zz_226 = img_reg_array_16_25_real;
        _zz_227 = img_reg_array_16_25_imag;
        _zz_228 = img_reg_array_17_25_real;
        _zz_229 = img_reg_array_17_25_imag;
        _zz_230 = img_reg_array_18_25_real;
        _zz_231 = img_reg_array_18_25_imag;
        _zz_232 = img_reg_array_19_25_real;
        _zz_233 = img_reg_array_19_25_imag;
        _zz_234 = img_reg_array_20_25_real;
        _zz_235 = img_reg_array_20_25_imag;
        _zz_236 = img_reg_array_21_25_real;
        _zz_237 = img_reg_array_21_25_imag;
        _zz_238 = img_reg_array_22_25_real;
        _zz_239 = img_reg_array_22_25_imag;
        _zz_240 = img_reg_array_23_25_real;
        _zz_241 = img_reg_array_23_25_imag;
        _zz_242 = img_reg_array_24_25_real;
        _zz_243 = img_reg_array_24_25_imag;
        _zz_244 = img_reg_array_25_25_real;
        _zz_245 = img_reg_array_25_25_imag;
        _zz_246 = img_reg_array_26_25_real;
        _zz_247 = img_reg_array_26_25_imag;
        _zz_248 = img_reg_array_27_25_real;
        _zz_249 = img_reg_array_27_25_imag;
        _zz_250 = img_reg_array_28_25_real;
        _zz_251 = img_reg_array_28_25_imag;
        _zz_252 = img_reg_array_29_25_real;
        _zz_253 = img_reg_array_29_25_imag;
        _zz_254 = img_reg_array_30_25_real;
        _zz_255 = img_reg_array_30_25_imag;
        _zz_256 = img_reg_array_31_25_real;
        _zz_257 = img_reg_array_31_25_imag;
        _zz_258 = img_reg_array_32_25_real;
        _zz_259 = img_reg_array_32_25_imag;
        _zz_260 = img_reg_array_33_25_real;
        _zz_261 = img_reg_array_33_25_imag;
        _zz_262 = img_reg_array_34_25_real;
        _zz_263 = img_reg_array_34_25_imag;
        _zz_264 = img_reg_array_35_25_real;
        _zz_265 = img_reg_array_35_25_imag;
        _zz_266 = img_reg_array_36_25_real;
        _zz_267 = img_reg_array_36_25_imag;
        _zz_268 = img_reg_array_37_25_real;
        _zz_269 = img_reg_array_37_25_imag;
        _zz_270 = img_reg_array_38_25_real;
        _zz_271 = img_reg_array_38_25_imag;
        _zz_272 = img_reg_array_39_25_real;
        _zz_273 = img_reg_array_39_25_imag;
        _zz_274 = img_reg_array_40_25_real;
        _zz_275 = img_reg_array_40_25_imag;
        _zz_276 = img_reg_array_41_25_real;
        _zz_277 = img_reg_array_41_25_imag;
        _zz_278 = img_reg_array_42_25_real;
        _zz_279 = img_reg_array_42_25_imag;
        _zz_280 = img_reg_array_43_25_real;
        _zz_281 = img_reg_array_43_25_imag;
        _zz_282 = img_reg_array_44_25_real;
        _zz_283 = img_reg_array_44_25_imag;
        _zz_284 = img_reg_array_45_25_real;
        _zz_285 = img_reg_array_45_25_imag;
        _zz_286 = img_reg_array_46_25_real;
        _zz_287 = img_reg_array_46_25_imag;
        _zz_288 = img_reg_array_47_25_real;
        _zz_289 = img_reg_array_47_25_imag;
        _zz_290 = img_reg_array_48_25_real;
        _zz_291 = img_reg_array_48_25_imag;
        _zz_292 = img_reg_array_49_25_real;
        _zz_293 = img_reg_array_49_25_imag;
        _zz_294 = img_reg_array_50_25_real;
        _zz_295 = img_reg_array_50_25_imag;
        _zz_296 = img_reg_array_51_25_real;
        _zz_297 = img_reg_array_51_25_imag;
        _zz_298 = img_reg_array_52_25_real;
        _zz_299 = img_reg_array_52_25_imag;
        _zz_300 = img_reg_array_53_25_real;
        _zz_301 = img_reg_array_53_25_imag;
        _zz_302 = img_reg_array_54_25_real;
        _zz_303 = img_reg_array_54_25_imag;
        _zz_304 = img_reg_array_55_25_real;
        _zz_305 = img_reg_array_55_25_imag;
        _zz_306 = img_reg_array_56_25_real;
        _zz_307 = img_reg_array_56_25_imag;
        _zz_308 = img_reg_array_57_25_real;
        _zz_309 = img_reg_array_57_25_imag;
        _zz_310 = img_reg_array_58_25_real;
        _zz_311 = img_reg_array_58_25_imag;
        _zz_312 = img_reg_array_59_25_real;
        _zz_313 = img_reg_array_59_25_imag;
        _zz_314 = img_reg_array_60_25_real;
        _zz_315 = img_reg_array_60_25_imag;
        _zz_316 = img_reg_array_61_25_real;
        _zz_317 = img_reg_array_61_25_imag;
        _zz_318 = img_reg_array_62_25_real;
        _zz_319 = img_reg_array_62_25_imag;
        _zz_320 = img_reg_array_63_25_real;
        _zz_321 = img_reg_array_63_25_imag;
      end
      6'b011010 : begin
        _zz_194 = img_reg_array_0_26_real;
        _zz_195 = img_reg_array_0_26_imag;
        _zz_196 = img_reg_array_1_26_real;
        _zz_197 = img_reg_array_1_26_imag;
        _zz_198 = img_reg_array_2_26_real;
        _zz_199 = img_reg_array_2_26_imag;
        _zz_200 = img_reg_array_3_26_real;
        _zz_201 = img_reg_array_3_26_imag;
        _zz_202 = img_reg_array_4_26_real;
        _zz_203 = img_reg_array_4_26_imag;
        _zz_204 = img_reg_array_5_26_real;
        _zz_205 = img_reg_array_5_26_imag;
        _zz_206 = img_reg_array_6_26_real;
        _zz_207 = img_reg_array_6_26_imag;
        _zz_208 = img_reg_array_7_26_real;
        _zz_209 = img_reg_array_7_26_imag;
        _zz_210 = img_reg_array_8_26_real;
        _zz_211 = img_reg_array_8_26_imag;
        _zz_212 = img_reg_array_9_26_real;
        _zz_213 = img_reg_array_9_26_imag;
        _zz_214 = img_reg_array_10_26_real;
        _zz_215 = img_reg_array_10_26_imag;
        _zz_216 = img_reg_array_11_26_real;
        _zz_217 = img_reg_array_11_26_imag;
        _zz_218 = img_reg_array_12_26_real;
        _zz_219 = img_reg_array_12_26_imag;
        _zz_220 = img_reg_array_13_26_real;
        _zz_221 = img_reg_array_13_26_imag;
        _zz_222 = img_reg_array_14_26_real;
        _zz_223 = img_reg_array_14_26_imag;
        _zz_224 = img_reg_array_15_26_real;
        _zz_225 = img_reg_array_15_26_imag;
        _zz_226 = img_reg_array_16_26_real;
        _zz_227 = img_reg_array_16_26_imag;
        _zz_228 = img_reg_array_17_26_real;
        _zz_229 = img_reg_array_17_26_imag;
        _zz_230 = img_reg_array_18_26_real;
        _zz_231 = img_reg_array_18_26_imag;
        _zz_232 = img_reg_array_19_26_real;
        _zz_233 = img_reg_array_19_26_imag;
        _zz_234 = img_reg_array_20_26_real;
        _zz_235 = img_reg_array_20_26_imag;
        _zz_236 = img_reg_array_21_26_real;
        _zz_237 = img_reg_array_21_26_imag;
        _zz_238 = img_reg_array_22_26_real;
        _zz_239 = img_reg_array_22_26_imag;
        _zz_240 = img_reg_array_23_26_real;
        _zz_241 = img_reg_array_23_26_imag;
        _zz_242 = img_reg_array_24_26_real;
        _zz_243 = img_reg_array_24_26_imag;
        _zz_244 = img_reg_array_25_26_real;
        _zz_245 = img_reg_array_25_26_imag;
        _zz_246 = img_reg_array_26_26_real;
        _zz_247 = img_reg_array_26_26_imag;
        _zz_248 = img_reg_array_27_26_real;
        _zz_249 = img_reg_array_27_26_imag;
        _zz_250 = img_reg_array_28_26_real;
        _zz_251 = img_reg_array_28_26_imag;
        _zz_252 = img_reg_array_29_26_real;
        _zz_253 = img_reg_array_29_26_imag;
        _zz_254 = img_reg_array_30_26_real;
        _zz_255 = img_reg_array_30_26_imag;
        _zz_256 = img_reg_array_31_26_real;
        _zz_257 = img_reg_array_31_26_imag;
        _zz_258 = img_reg_array_32_26_real;
        _zz_259 = img_reg_array_32_26_imag;
        _zz_260 = img_reg_array_33_26_real;
        _zz_261 = img_reg_array_33_26_imag;
        _zz_262 = img_reg_array_34_26_real;
        _zz_263 = img_reg_array_34_26_imag;
        _zz_264 = img_reg_array_35_26_real;
        _zz_265 = img_reg_array_35_26_imag;
        _zz_266 = img_reg_array_36_26_real;
        _zz_267 = img_reg_array_36_26_imag;
        _zz_268 = img_reg_array_37_26_real;
        _zz_269 = img_reg_array_37_26_imag;
        _zz_270 = img_reg_array_38_26_real;
        _zz_271 = img_reg_array_38_26_imag;
        _zz_272 = img_reg_array_39_26_real;
        _zz_273 = img_reg_array_39_26_imag;
        _zz_274 = img_reg_array_40_26_real;
        _zz_275 = img_reg_array_40_26_imag;
        _zz_276 = img_reg_array_41_26_real;
        _zz_277 = img_reg_array_41_26_imag;
        _zz_278 = img_reg_array_42_26_real;
        _zz_279 = img_reg_array_42_26_imag;
        _zz_280 = img_reg_array_43_26_real;
        _zz_281 = img_reg_array_43_26_imag;
        _zz_282 = img_reg_array_44_26_real;
        _zz_283 = img_reg_array_44_26_imag;
        _zz_284 = img_reg_array_45_26_real;
        _zz_285 = img_reg_array_45_26_imag;
        _zz_286 = img_reg_array_46_26_real;
        _zz_287 = img_reg_array_46_26_imag;
        _zz_288 = img_reg_array_47_26_real;
        _zz_289 = img_reg_array_47_26_imag;
        _zz_290 = img_reg_array_48_26_real;
        _zz_291 = img_reg_array_48_26_imag;
        _zz_292 = img_reg_array_49_26_real;
        _zz_293 = img_reg_array_49_26_imag;
        _zz_294 = img_reg_array_50_26_real;
        _zz_295 = img_reg_array_50_26_imag;
        _zz_296 = img_reg_array_51_26_real;
        _zz_297 = img_reg_array_51_26_imag;
        _zz_298 = img_reg_array_52_26_real;
        _zz_299 = img_reg_array_52_26_imag;
        _zz_300 = img_reg_array_53_26_real;
        _zz_301 = img_reg_array_53_26_imag;
        _zz_302 = img_reg_array_54_26_real;
        _zz_303 = img_reg_array_54_26_imag;
        _zz_304 = img_reg_array_55_26_real;
        _zz_305 = img_reg_array_55_26_imag;
        _zz_306 = img_reg_array_56_26_real;
        _zz_307 = img_reg_array_56_26_imag;
        _zz_308 = img_reg_array_57_26_real;
        _zz_309 = img_reg_array_57_26_imag;
        _zz_310 = img_reg_array_58_26_real;
        _zz_311 = img_reg_array_58_26_imag;
        _zz_312 = img_reg_array_59_26_real;
        _zz_313 = img_reg_array_59_26_imag;
        _zz_314 = img_reg_array_60_26_real;
        _zz_315 = img_reg_array_60_26_imag;
        _zz_316 = img_reg_array_61_26_real;
        _zz_317 = img_reg_array_61_26_imag;
        _zz_318 = img_reg_array_62_26_real;
        _zz_319 = img_reg_array_62_26_imag;
        _zz_320 = img_reg_array_63_26_real;
        _zz_321 = img_reg_array_63_26_imag;
      end
      6'b011011 : begin
        _zz_194 = img_reg_array_0_27_real;
        _zz_195 = img_reg_array_0_27_imag;
        _zz_196 = img_reg_array_1_27_real;
        _zz_197 = img_reg_array_1_27_imag;
        _zz_198 = img_reg_array_2_27_real;
        _zz_199 = img_reg_array_2_27_imag;
        _zz_200 = img_reg_array_3_27_real;
        _zz_201 = img_reg_array_3_27_imag;
        _zz_202 = img_reg_array_4_27_real;
        _zz_203 = img_reg_array_4_27_imag;
        _zz_204 = img_reg_array_5_27_real;
        _zz_205 = img_reg_array_5_27_imag;
        _zz_206 = img_reg_array_6_27_real;
        _zz_207 = img_reg_array_6_27_imag;
        _zz_208 = img_reg_array_7_27_real;
        _zz_209 = img_reg_array_7_27_imag;
        _zz_210 = img_reg_array_8_27_real;
        _zz_211 = img_reg_array_8_27_imag;
        _zz_212 = img_reg_array_9_27_real;
        _zz_213 = img_reg_array_9_27_imag;
        _zz_214 = img_reg_array_10_27_real;
        _zz_215 = img_reg_array_10_27_imag;
        _zz_216 = img_reg_array_11_27_real;
        _zz_217 = img_reg_array_11_27_imag;
        _zz_218 = img_reg_array_12_27_real;
        _zz_219 = img_reg_array_12_27_imag;
        _zz_220 = img_reg_array_13_27_real;
        _zz_221 = img_reg_array_13_27_imag;
        _zz_222 = img_reg_array_14_27_real;
        _zz_223 = img_reg_array_14_27_imag;
        _zz_224 = img_reg_array_15_27_real;
        _zz_225 = img_reg_array_15_27_imag;
        _zz_226 = img_reg_array_16_27_real;
        _zz_227 = img_reg_array_16_27_imag;
        _zz_228 = img_reg_array_17_27_real;
        _zz_229 = img_reg_array_17_27_imag;
        _zz_230 = img_reg_array_18_27_real;
        _zz_231 = img_reg_array_18_27_imag;
        _zz_232 = img_reg_array_19_27_real;
        _zz_233 = img_reg_array_19_27_imag;
        _zz_234 = img_reg_array_20_27_real;
        _zz_235 = img_reg_array_20_27_imag;
        _zz_236 = img_reg_array_21_27_real;
        _zz_237 = img_reg_array_21_27_imag;
        _zz_238 = img_reg_array_22_27_real;
        _zz_239 = img_reg_array_22_27_imag;
        _zz_240 = img_reg_array_23_27_real;
        _zz_241 = img_reg_array_23_27_imag;
        _zz_242 = img_reg_array_24_27_real;
        _zz_243 = img_reg_array_24_27_imag;
        _zz_244 = img_reg_array_25_27_real;
        _zz_245 = img_reg_array_25_27_imag;
        _zz_246 = img_reg_array_26_27_real;
        _zz_247 = img_reg_array_26_27_imag;
        _zz_248 = img_reg_array_27_27_real;
        _zz_249 = img_reg_array_27_27_imag;
        _zz_250 = img_reg_array_28_27_real;
        _zz_251 = img_reg_array_28_27_imag;
        _zz_252 = img_reg_array_29_27_real;
        _zz_253 = img_reg_array_29_27_imag;
        _zz_254 = img_reg_array_30_27_real;
        _zz_255 = img_reg_array_30_27_imag;
        _zz_256 = img_reg_array_31_27_real;
        _zz_257 = img_reg_array_31_27_imag;
        _zz_258 = img_reg_array_32_27_real;
        _zz_259 = img_reg_array_32_27_imag;
        _zz_260 = img_reg_array_33_27_real;
        _zz_261 = img_reg_array_33_27_imag;
        _zz_262 = img_reg_array_34_27_real;
        _zz_263 = img_reg_array_34_27_imag;
        _zz_264 = img_reg_array_35_27_real;
        _zz_265 = img_reg_array_35_27_imag;
        _zz_266 = img_reg_array_36_27_real;
        _zz_267 = img_reg_array_36_27_imag;
        _zz_268 = img_reg_array_37_27_real;
        _zz_269 = img_reg_array_37_27_imag;
        _zz_270 = img_reg_array_38_27_real;
        _zz_271 = img_reg_array_38_27_imag;
        _zz_272 = img_reg_array_39_27_real;
        _zz_273 = img_reg_array_39_27_imag;
        _zz_274 = img_reg_array_40_27_real;
        _zz_275 = img_reg_array_40_27_imag;
        _zz_276 = img_reg_array_41_27_real;
        _zz_277 = img_reg_array_41_27_imag;
        _zz_278 = img_reg_array_42_27_real;
        _zz_279 = img_reg_array_42_27_imag;
        _zz_280 = img_reg_array_43_27_real;
        _zz_281 = img_reg_array_43_27_imag;
        _zz_282 = img_reg_array_44_27_real;
        _zz_283 = img_reg_array_44_27_imag;
        _zz_284 = img_reg_array_45_27_real;
        _zz_285 = img_reg_array_45_27_imag;
        _zz_286 = img_reg_array_46_27_real;
        _zz_287 = img_reg_array_46_27_imag;
        _zz_288 = img_reg_array_47_27_real;
        _zz_289 = img_reg_array_47_27_imag;
        _zz_290 = img_reg_array_48_27_real;
        _zz_291 = img_reg_array_48_27_imag;
        _zz_292 = img_reg_array_49_27_real;
        _zz_293 = img_reg_array_49_27_imag;
        _zz_294 = img_reg_array_50_27_real;
        _zz_295 = img_reg_array_50_27_imag;
        _zz_296 = img_reg_array_51_27_real;
        _zz_297 = img_reg_array_51_27_imag;
        _zz_298 = img_reg_array_52_27_real;
        _zz_299 = img_reg_array_52_27_imag;
        _zz_300 = img_reg_array_53_27_real;
        _zz_301 = img_reg_array_53_27_imag;
        _zz_302 = img_reg_array_54_27_real;
        _zz_303 = img_reg_array_54_27_imag;
        _zz_304 = img_reg_array_55_27_real;
        _zz_305 = img_reg_array_55_27_imag;
        _zz_306 = img_reg_array_56_27_real;
        _zz_307 = img_reg_array_56_27_imag;
        _zz_308 = img_reg_array_57_27_real;
        _zz_309 = img_reg_array_57_27_imag;
        _zz_310 = img_reg_array_58_27_real;
        _zz_311 = img_reg_array_58_27_imag;
        _zz_312 = img_reg_array_59_27_real;
        _zz_313 = img_reg_array_59_27_imag;
        _zz_314 = img_reg_array_60_27_real;
        _zz_315 = img_reg_array_60_27_imag;
        _zz_316 = img_reg_array_61_27_real;
        _zz_317 = img_reg_array_61_27_imag;
        _zz_318 = img_reg_array_62_27_real;
        _zz_319 = img_reg_array_62_27_imag;
        _zz_320 = img_reg_array_63_27_real;
        _zz_321 = img_reg_array_63_27_imag;
      end
      6'b011100 : begin
        _zz_194 = img_reg_array_0_28_real;
        _zz_195 = img_reg_array_0_28_imag;
        _zz_196 = img_reg_array_1_28_real;
        _zz_197 = img_reg_array_1_28_imag;
        _zz_198 = img_reg_array_2_28_real;
        _zz_199 = img_reg_array_2_28_imag;
        _zz_200 = img_reg_array_3_28_real;
        _zz_201 = img_reg_array_3_28_imag;
        _zz_202 = img_reg_array_4_28_real;
        _zz_203 = img_reg_array_4_28_imag;
        _zz_204 = img_reg_array_5_28_real;
        _zz_205 = img_reg_array_5_28_imag;
        _zz_206 = img_reg_array_6_28_real;
        _zz_207 = img_reg_array_6_28_imag;
        _zz_208 = img_reg_array_7_28_real;
        _zz_209 = img_reg_array_7_28_imag;
        _zz_210 = img_reg_array_8_28_real;
        _zz_211 = img_reg_array_8_28_imag;
        _zz_212 = img_reg_array_9_28_real;
        _zz_213 = img_reg_array_9_28_imag;
        _zz_214 = img_reg_array_10_28_real;
        _zz_215 = img_reg_array_10_28_imag;
        _zz_216 = img_reg_array_11_28_real;
        _zz_217 = img_reg_array_11_28_imag;
        _zz_218 = img_reg_array_12_28_real;
        _zz_219 = img_reg_array_12_28_imag;
        _zz_220 = img_reg_array_13_28_real;
        _zz_221 = img_reg_array_13_28_imag;
        _zz_222 = img_reg_array_14_28_real;
        _zz_223 = img_reg_array_14_28_imag;
        _zz_224 = img_reg_array_15_28_real;
        _zz_225 = img_reg_array_15_28_imag;
        _zz_226 = img_reg_array_16_28_real;
        _zz_227 = img_reg_array_16_28_imag;
        _zz_228 = img_reg_array_17_28_real;
        _zz_229 = img_reg_array_17_28_imag;
        _zz_230 = img_reg_array_18_28_real;
        _zz_231 = img_reg_array_18_28_imag;
        _zz_232 = img_reg_array_19_28_real;
        _zz_233 = img_reg_array_19_28_imag;
        _zz_234 = img_reg_array_20_28_real;
        _zz_235 = img_reg_array_20_28_imag;
        _zz_236 = img_reg_array_21_28_real;
        _zz_237 = img_reg_array_21_28_imag;
        _zz_238 = img_reg_array_22_28_real;
        _zz_239 = img_reg_array_22_28_imag;
        _zz_240 = img_reg_array_23_28_real;
        _zz_241 = img_reg_array_23_28_imag;
        _zz_242 = img_reg_array_24_28_real;
        _zz_243 = img_reg_array_24_28_imag;
        _zz_244 = img_reg_array_25_28_real;
        _zz_245 = img_reg_array_25_28_imag;
        _zz_246 = img_reg_array_26_28_real;
        _zz_247 = img_reg_array_26_28_imag;
        _zz_248 = img_reg_array_27_28_real;
        _zz_249 = img_reg_array_27_28_imag;
        _zz_250 = img_reg_array_28_28_real;
        _zz_251 = img_reg_array_28_28_imag;
        _zz_252 = img_reg_array_29_28_real;
        _zz_253 = img_reg_array_29_28_imag;
        _zz_254 = img_reg_array_30_28_real;
        _zz_255 = img_reg_array_30_28_imag;
        _zz_256 = img_reg_array_31_28_real;
        _zz_257 = img_reg_array_31_28_imag;
        _zz_258 = img_reg_array_32_28_real;
        _zz_259 = img_reg_array_32_28_imag;
        _zz_260 = img_reg_array_33_28_real;
        _zz_261 = img_reg_array_33_28_imag;
        _zz_262 = img_reg_array_34_28_real;
        _zz_263 = img_reg_array_34_28_imag;
        _zz_264 = img_reg_array_35_28_real;
        _zz_265 = img_reg_array_35_28_imag;
        _zz_266 = img_reg_array_36_28_real;
        _zz_267 = img_reg_array_36_28_imag;
        _zz_268 = img_reg_array_37_28_real;
        _zz_269 = img_reg_array_37_28_imag;
        _zz_270 = img_reg_array_38_28_real;
        _zz_271 = img_reg_array_38_28_imag;
        _zz_272 = img_reg_array_39_28_real;
        _zz_273 = img_reg_array_39_28_imag;
        _zz_274 = img_reg_array_40_28_real;
        _zz_275 = img_reg_array_40_28_imag;
        _zz_276 = img_reg_array_41_28_real;
        _zz_277 = img_reg_array_41_28_imag;
        _zz_278 = img_reg_array_42_28_real;
        _zz_279 = img_reg_array_42_28_imag;
        _zz_280 = img_reg_array_43_28_real;
        _zz_281 = img_reg_array_43_28_imag;
        _zz_282 = img_reg_array_44_28_real;
        _zz_283 = img_reg_array_44_28_imag;
        _zz_284 = img_reg_array_45_28_real;
        _zz_285 = img_reg_array_45_28_imag;
        _zz_286 = img_reg_array_46_28_real;
        _zz_287 = img_reg_array_46_28_imag;
        _zz_288 = img_reg_array_47_28_real;
        _zz_289 = img_reg_array_47_28_imag;
        _zz_290 = img_reg_array_48_28_real;
        _zz_291 = img_reg_array_48_28_imag;
        _zz_292 = img_reg_array_49_28_real;
        _zz_293 = img_reg_array_49_28_imag;
        _zz_294 = img_reg_array_50_28_real;
        _zz_295 = img_reg_array_50_28_imag;
        _zz_296 = img_reg_array_51_28_real;
        _zz_297 = img_reg_array_51_28_imag;
        _zz_298 = img_reg_array_52_28_real;
        _zz_299 = img_reg_array_52_28_imag;
        _zz_300 = img_reg_array_53_28_real;
        _zz_301 = img_reg_array_53_28_imag;
        _zz_302 = img_reg_array_54_28_real;
        _zz_303 = img_reg_array_54_28_imag;
        _zz_304 = img_reg_array_55_28_real;
        _zz_305 = img_reg_array_55_28_imag;
        _zz_306 = img_reg_array_56_28_real;
        _zz_307 = img_reg_array_56_28_imag;
        _zz_308 = img_reg_array_57_28_real;
        _zz_309 = img_reg_array_57_28_imag;
        _zz_310 = img_reg_array_58_28_real;
        _zz_311 = img_reg_array_58_28_imag;
        _zz_312 = img_reg_array_59_28_real;
        _zz_313 = img_reg_array_59_28_imag;
        _zz_314 = img_reg_array_60_28_real;
        _zz_315 = img_reg_array_60_28_imag;
        _zz_316 = img_reg_array_61_28_real;
        _zz_317 = img_reg_array_61_28_imag;
        _zz_318 = img_reg_array_62_28_real;
        _zz_319 = img_reg_array_62_28_imag;
        _zz_320 = img_reg_array_63_28_real;
        _zz_321 = img_reg_array_63_28_imag;
      end
      6'b011101 : begin
        _zz_194 = img_reg_array_0_29_real;
        _zz_195 = img_reg_array_0_29_imag;
        _zz_196 = img_reg_array_1_29_real;
        _zz_197 = img_reg_array_1_29_imag;
        _zz_198 = img_reg_array_2_29_real;
        _zz_199 = img_reg_array_2_29_imag;
        _zz_200 = img_reg_array_3_29_real;
        _zz_201 = img_reg_array_3_29_imag;
        _zz_202 = img_reg_array_4_29_real;
        _zz_203 = img_reg_array_4_29_imag;
        _zz_204 = img_reg_array_5_29_real;
        _zz_205 = img_reg_array_5_29_imag;
        _zz_206 = img_reg_array_6_29_real;
        _zz_207 = img_reg_array_6_29_imag;
        _zz_208 = img_reg_array_7_29_real;
        _zz_209 = img_reg_array_7_29_imag;
        _zz_210 = img_reg_array_8_29_real;
        _zz_211 = img_reg_array_8_29_imag;
        _zz_212 = img_reg_array_9_29_real;
        _zz_213 = img_reg_array_9_29_imag;
        _zz_214 = img_reg_array_10_29_real;
        _zz_215 = img_reg_array_10_29_imag;
        _zz_216 = img_reg_array_11_29_real;
        _zz_217 = img_reg_array_11_29_imag;
        _zz_218 = img_reg_array_12_29_real;
        _zz_219 = img_reg_array_12_29_imag;
        _zz_220 = img_reg_array_13_29_real;
        _zz_221 = img_reg_array_13_29_imag;
        _zz_222 = img_reg_array_14_29_real;
        _zz_223 = img_reg_array_14_29_imag;
        _zz_224 = img_reg_array_15_29_real;
        _zz_225 = img_reg_array_15_29_imag;
        _zz_226 = img_reg_array_16_29_real;
        _zz_227 = img_reg_array_16_29_imag;
        _zz_228 = img_reg_array_17_29_real;
        _zz_229 = img_reg_array_17_29_imag;
        _zz_230 = img_reg_array_18_29_real;
        _zz_231 = img_reg_array_18_29_imag;
        _zz_232 = img_reg_array_19_29_real;
        _zz_233 = img_reg_array_19_29_imag;
        _zz_234 = img_reg_array_20_29_real;
        _zz_235 = img_reg_array_20_29_imag;
        _zz_236 = img_reg_array_21_29_real;
        _zz_237 = img_reg_array_21_29_imag;
        _zz_238 = img_reg_array_22_29_real;
        _zz_239 = img_reg_array_22_29_imag;
        _zz_240 = img_reg_array_23_29_real;
        _zz_241 = img_reg_array_23_29_imag;
        _zz_242 = img_reg_array_24_29_real;
        _zz_243 = img_reg_array_24_29_imag;
        _zz_244 = img_reg_array_25_29_real;
        _zz_245 = img_reg_array_25_29_imag;
        _zz_246 = img_reg_array_26_29_real;
        _zz_247 = img_reg_array_26_29_imag;
        _zz_248 = img_reg_array_27_29_real;
        _zz_249 = img_reg_array_27_29_imag;
        _zz_250 = img_reg_array_28_29_real;
        _zz_251 = img_reg_array_28_29_imag;
        _zz_252 = img_reg_array_29_29_real;
        _zz_253 = img_reg_array_29_29_imag;
        _zz_254 = img_reg_array_30_29_real;
        _zz_255 = img_reg_array_30_29_imag;
        _zz_256 = img_reg_array_31_29_real;
        _zz_257 = img_reg_array_31_29_imag;
        _zz_258 = img_reg_array_32_29_real;
        _zz_259 = img_reg_array_32_29_imag;
        _zz_260 = img_reg_array_33_29_real;
        _zz_261 = img_reg_array_33_29_imag;
        _zz_262 = img_reg_array_34_29_real;
        _zz_263 = img_reg_array_34_29_imag;
        _zz_264 = img_reg_array_35_29_real;
        _zz_265 = img_reg_array_35_29_imag;
        _zz_266 = img_reg_array_36_29_real;
        _zz_267 = img_reg_array_36_29_imag;
        _zz_268 = img_reg_array_37_29_real;
        _zz_269 = img_reg_array_37_29_imag;
        _zz_270 = img_reg_array_38_29_real;
        _zz_271 = img_reg_array_38_29_imag;
        _zz_272 = img_reg_array_39_29_real;
        _zz_273 = img_reg_array_39_29_imag;
        _zz_274 = img_reg_array_40_29_real;
        _zz_275 = img_reg_array_40_29_imag;
        _zz_276 = img_reg_array_41_29_real;
        _zz_277 = img_reg_array_41_29_imag;
        _zz_278 = img_reg_array_42_29_real;
        _zz_279 = img_reg_array_42_29_imag;
        _zz_280 = img_reg_array_43_29_real;
        _zz_281 = img_reg_array_43_29_imag;
        _zz_282 = img_reg_array_44_29_real;
        _zz_283 = img_reg_array_44_29_imag;
        _zz_284 = img_reg_array_45_29_real;
        _zz_285 = img_reg_array_45_29_imag;
        _zz_286 = img_reg_array_46_29_real;
        _zz_287 = img_reg_array_46_29_imag;
        _zz_288 = img_reg_array_47_29_real;
        _zz_289 = img_reg_array_47_29_imag;
        _zz_290 = img_reg_array_48_29_real;
        _zz_291 = img_reg_array_48_29_imag;
        _zz_292 = img_reg_array_49_29_real;
        _zz_293 = img_reg_array_49_29_imag;
        _zz_294 = img_reg_array_50_29_real;
        _zz_295 = img_reg_array_50_29_imag;
        _zz_296 = img_reg_array_51_29_real;
        _zz_297 = img_reg_array_51_29_imag;
        _zz_298 = img_reg_array_52_29_real;
        _zz_299 = img_reg_array_52_29_imag;
        _zz_300 = img_reg_array_53_29_real;
        _zz_301 = img_reg_array_53_29_imag;
        _zz_302 = img_reg_array_54_29_real;
        _zz_303 = img_reg_array_54_29_imag;
        _zz_304 = img_reg_array_55_29_real;
        _zz_305 = img_reg_array_55_29_imag;
        _zz_306 = img_reg_array_56_29_real;
        _zz_307 = img_reg_array_56_29_imag;
        _zz_308 = img_reg_array_57_29_real;
        _zz_309 = img_reg_array_57_29_imag;
        _zz_310 = img_reg_array_58_29_real;
        _zz_311 = img_reg_array_58_29_imag;
        _zz_312 = img_reg_array_59_29_real;
        _zz_313 = img_reg_array_59_29_imag;
        _zz_314 = img_reg_array_60_29_real;
        _zz_315 = img_reg_array_60_29_imag;
        _zz_316 = img_reg_array_61_29_real;
        _zz_317 = img_reg_array_61_29_imag;
        _zz_318 = img_reg_array_62_29_real;
        _zz_319 = img_reg_array_62_29_imag;
        _zz_320 = img_reg_array_63_29_real;
        _zz_321 = img_reg_array_63_29_imag;
      end
      6'b011110 : begin
        _zz_194 = img_reg_array_0_30_real;
        _zz_195 = img_reg_array_0_30_imag;
        _zz_196 = img_reg_array_1_30_real;
        _zz_197 = img_reg_array_1_30_imag;
        _zz_198 = img_reg_array_2_30_real;
        _zz_199 = img_reg_array_2_30_imag;
        _zz_200 = img_reg_array_3_30_real;
        _zz_201 = img_reg_array_3_30_imag;
        _zz_202 = img_reg_array_4_30_real;
        _zz_203 = img_reg_array_4_30_imag;
        _zz_204 = img_reg_array_5_30_real;
        _zz_205 = img_reg_array_5_30_imag;
        _zz_206 = img_reg_array_6_30_real;
        _zz_207 = img_reg_array_6_30_imag;
        _zz_208 = img_reg_array_7_30_real;
        _zz_209 = img_reg_array_7_30_imag;
        _zz_210 = img_reg_array_8_30_real;
        _zz_211 = img_reg_array_8_30_imag;
        _zz_212 = img_reg_array_9_30_real;
        _zz_213 = img_reg_array_9_30_imag;
        _zz_214 = img_reg_array_10_30_real;
        _zz_215 = img_reg_array_10_30_imag;
        _zz_216 = img_reg_array_11_30_real;
        _zz_217 = img_reg_array_11_30_imag;
        _zz_218 = img_reg_array_12_30_real;
        _zz_219 = img_reg_array_12_30_imag;
        _zz_220 = img_reg_array_13_30_real;
        _zz_221 = img_reg_array_13_30_imag;
        _zz_222 = img_reg_array_14_30_real;
        _zz_223 = img_reg_array_14_30_imag;
        _zz_224 = img_reg_array_15_30_real;
        _zz_225 = img_reg_array_15_30_imag;
        _zz_226 = img_reg_array_16_30_real;
        _zz_227 = img_reg_array_16_30_imag;
        _zz_228 = img_reg_array_17_30_real;
        _zz_229 = img_reg_array_17_30_imag;
        _zz_230 = img_reg_array_18_30_real;
        _zz_231 = img_reg_array_18_30_imag;
        _zz_232 = img_reg_array_19_30_real;
        _zz_233 = img_reg_array_19_30_imag;
        _zz_234 = img_reg_array_20_30_real;
        _zz_235 = img_reg_array_20_30_imag;
        _zz_236 = img_reg_array_21_30_real;
        _zz_237 = img_reg_array_21_30_imag;
        _zz_238 = img_reg_array_22_30_real;
        _zz_239 = img_reg_array_22_30_imag;
        _zz_240 = img_reg_array_23_30_real;
        _zz_241 = img_reg_array_23_30_imag;
        _zz_242 = img_reg_array_24_30_real;
        _zz_243 = img_reg_array_24_30_imag;
        _zz_244 = img_reg_array_25_30_real;
        _zz_245 = img_reg_array_25_30_imag;
        _zz_246 = img_reg_array_26_30_real;
        _zz_247 = img_reg_array_26_30_imag;
        _zz_248 = img_reg_array_27_30_real;
        _zz_249 = img_reg_array_27_30_imag;
        _zz_250 = img_reg_array_28_30_real;
        _zz_251 = img_reg_array_28_30_imag;
        _zz_252 = img_reg_array_29_30_real;
        _zz_253 = img_reg_array_29_30_imag;
        _zz_254 = img_reg_array_30_30_real;
        _zz_255 = img_reg_array_30_30_imag;
        _zz_256 = img_reg_array_31_30_real;
        _zz_257 = img_reg_array_31_30_imag;
        _zz_258 = img_reg_array_32_30_real;
        _zz_259 = img_reg_array_32_30_imag;
        _zz_260 = img_reg_array_33_30_real;
        _zz_261 = img_reg_array_33_30_imag;
        _zz_262 = img_reg_array_34_30_real;
        _zz_263 = img_reg_array_34_30_imag;
        _zz_264 = img_reg_array_35_30_real;
        _zz_265 = img_reg_array_35_30_imag;
        _zz_266 = img_reg_array_36_30_real;
        _zz_267 = img_reg_array_36_30_imag;
        _zz_268 = img_reg_array_37_30_real;
        _zz_269 = img_reg_array_37_30_imag;
        _zz_270 = img_reg_array_38_30_real;
        _zz_271 = img_reg_array_38_30_imag;
        _zz_272 = img_reg_array_39_30_real;
        _zz_273 = img_reg_array_39_30_imag;
        _zz_274 = img_reg_array_40_30_real;
        _zz_275 = img_reg_array_40_30_imag;
        _zz_276 = img_reg_array_41_30_real;
        _zz_277 = img_reg_array_41_30_imag;
        _zz_278 = img_reg_array_42_30_real;
        _zz_279 = img_reg_array_42_30_imag;
        _zz_280 = img_reg_array_43_30_real;
        _zz_281 = img_reg_array_43_30_imag;
        _zz_282 = img_reg_array_44_30_real;
        _zz_283 = img_reg_array_44_30_imag;
        _zz_284 = img_reg_array_45_30_real;
        _zz_285 = img_reg_array_45_30_imag;
        _zz_286 = img_reg_array_46_30_real;
        _zz_287 = img_reg_array_46_30_imag;
        _zz_288 = img_reg_array_47_30_real;
        _zz_289 = img_reg_array_47_30_imag;
        _zz_290 = img_reg_array_48_30_real;
        _zz_291 = img_reg_array_48_30_imag;
        _zz_292 = img_reg_array_49_30_real;
        _zz_293 = img_reg_array_49_30_imag;
        _zz_294 = img_reg_array_50_30_real;
        _zz_295 = img_reg_array_50_30_imag;
        _zz_296 = img_reg_array_51_30_real;
        _zz_297 = img_reg_array_51_30_imag;
        _zz_298 = img_reg_array_52_30_real;
        _zz_299 = img_reg_array_52_30_imag;
        _zz_300 = img_reg_array_53_30_real;
        _zz_301 = img_reg_array_53_30_imag;
        _zz_302 = img_reg_array_54_30_real;
        _zz_303 = img_reg_array_54_30_imag;
        _zz_304 = img_reg_array_55_30_real;
        _zz_305 = img_reg_array_55_30_imag;
        _zz_306 = img_reg_array_56_30_real;
        _zz_307 = img_reg_array_56_30_imag;
        _zz_308 = img_reg_array_57_30_real;
        _zz_309 = img_reg_array_57_30_imag;
        _zz_310 = img_reg_array_58_30_real;
        _zz_311 = img_reg_array_58_30_imag;
        _zz_312 = img_reg_array_59_30_real;
        _zz_313 = img_reg_array_59_30_imag;
        _zz_314 = img_reg_array_60_30_real;
        _zz_315 = img_reg_array_60_30_imag;
        _zz_316 = img_reg_array_61_30_real;
        _zz_317 = img_reg_array_61_30_imag;
        _zz_318 = img_reg_array_62_30_real;
        _zz_319 = img_reg_array_62_30_imag;
        _zz_320 = img_reg_array_63_30_real;
        _zz_321 = img_reg_array_63_30_imag;
      end
      6'b011111 : begin
        _zz_194 = img_reg_array_0_31_real;
        _zz_195 = img_reg_array_0_31_imag;
        _zz_196 = img_reg_array_1_31_real;
        _zz_197 = img_reg_array_1_31_imag;
        _zz_198 = img_reg_array_2_31_real;
        _zz_199 = img_reg_array_2_31_imag;
        _zz_200 = img_reg_array_3_31_real;
        _zz_201 = img_reg_array_3_31_imag;
        _zz_202 = img_reg_array_4_31_real;
        _zz_203 = img_reg_array_4_31_imag;
        _zz_204 = img_reg_array_5_31_real;
        _zz_205 = img_reg_array_5_31_imag;
        _zz_206 = img_reg_array_6_31_real;
        _zz_207 = img_reg_array_6_31_imag;
        _zz_208 = img_reg_array_7_31_real;
        _zz_209 = img_reg_array_7_31_imag;
        _zz_210 = img_reg_array_8_31_real;
        _zz_211 = img_reg_array_8_31_imag;
        _zz_212 = img_reg_array_9_31_real;
        _zz_213 = img_reg_array_9_31_imag;
        _zz_214 = img_reg_array_10_31_real;
        _zz_215 = img_reg_array_10_31_imag;
        _zz_216 = img_reg_array_11_31_real;
        _zz_217 = img_reg_array_11_31_imag;
        _zz_218 = img_reg_array_12_31_real;
        _zz_219 = img_reg_array_12_31_imag;
        _zz_220 = img_reg_array_13_31_real;
        _zz_221 = img_reg_array_13_31_imag;
        _zz_222 = img_reg_array_14_31_real;
        _zz_223 = img_reg_array_14_31_imag;
        _zz_224 = img_reg_array_15_31_real;
        _zz_225 = img_reg_array_15_31_imag;
        _zz_226 = img_reg_array_16_31_real;
        _zz_227 = img_reg_array_16_31_imag;
        _zz_228 = img_reg_array_17_31_real;
        _zz_229 = img_reg_array_17_31_imag;
        _zz_230 = img_reg_array_18_31_real;
        _zz_231 = img_reg_array_18_31_imag;
        _zz_232 = img_reg_array_19_31_real;
        _zz_233 = img_reg_array_19_31_imag;
        _zz_234 = img_reg_array_20_31_real;
        _zz_235 = img_reg_array_20_31_imag;
        _zz_236 = img_reg_array_21_31_real;
        _zz_237 = img_reg_array_21_31_imag;
        _zz_238 = img_reg_array_22_31_real;
        _zz_239 = img_reg_array_22_31_imag;
        _zz_240 = img_reg_array_23_31_real;
        _zz_241 = img_reg_array_23_31_imag;
        _zz_242 = img_reg_array_24_31_real;
        _zz_243 = img_reg_array_24_31_imag;
        _zz_244 = img_reg_array_25_31_real;
        _zz_245 = img_reg_array_25_31_imag;
        _zz_246 = img_reg_array_26_31_real;
        _zz_247 = img_reg_array_26_31_imag;
        _zz_248 = img_reg_array_27_31_real;
        _zz_249 = img_reg_array_27_31_imag;
        _zz_250 = img_reg_array_28_31_real;
        _zz_251 = img_reg_array_28_31_imag;
        _zz_252 = img_reg_array_29_31_real;
        _zz_253 = img_reg_array_29_31_imag;
        _zz_254 = img_reg_array_30_31_real;
        _zz_255 = img_reg_array_30_31_imag;
        _zz_256 = img_reg_array_31_31_real;
        _zz_257 = img_reg_array_31_31_imag;
        _zz_258 = img_reg_array_32_31_real;
        _zz_259 = img_reg_array_32_31_imag;
        _zz_260 = img_reg_array_33_31_real;
        _zz_261 = img_reg_array_33_31_imag;
        _zz_262 = img_reg_array_34_31_real;
        _zz_263 = img_reg_array_34_31_imag;
        _zz_264 = img_reg_array_35_31_real;
        _zz_265 = img_reg_array_35_31_imag;
        _zz_266 = img_reg_array_36_31_real;
        _zz_267 = img_reg_array_36_31_imag;
        _zz_268 = img_reg_array_37_31_real;
        _zz_269 = img_reg_array_37_31_imag;
        _zz_270 = img_reg_array_38_31_real;
        _zz_271 = img_reg_array_38_31_imag;
        _zz_272 = img_reg_array_39_31_real;
        _zz_273 = img_reg_array_39_31_imag;
        _zz_274 = img_reg_array_40_31_real;
        _zz_275 = img_reg_array_40_31_imag;
        _zz_276 = img_reg_array_41_31_real;
        _zz_277 = img_reg_array_41_31_imag;
        _zz_278 = img_reg_array_42_31_real;
        _zz_279 = img_reg_array_42_31_imag;
        _zz_280 = img_reg_array_43_31_real;
        _zz_281 = img_reg_array_43_31_imag;
        _zz_282 = img_reg_array_44_31_real;
        _zz_283 = img_reg_array_44_31_imag;
        _zz_284 = img_reg_array_45_31_real;
        _zz_285 = img_reg_array_45_31_imag;
        _zz_286 = img_reg_array_46_31_real;
        _zz_287 = img_reg_array_46_31_imag;
        _zz_288 = img_reg_array_47_31_real;
        _zz_289 = img_reg_array_47_31_imag;
        _zz_290 = img_reg_array_48_31_real;
        _zz_291 = img_reg_array_48_31_imag;
        _zz_292 = img_reg_array_49_31_real;
        _zz_293 = img_reg_array_49_31_imag;
        _zz_294 = img_reg_array_50_31_real;
        _zz_295 = img_reg_array_50_31_imag;
        _zz_296 = img_reg_array_51_31_real;
        _zz_297 = img_reg_array_51_31_imag;
        _zz_298 = img_reg_array_52_31_real;
        _zz_299 = img_reg_array_52_31_imag;
        _zz_300 = img_reg_array_53_31_real;
        _zz_301 = img_reg_array_53_31_imag;
        _zz_302 = img_reg_array_54_31_real;
        _zz_303 = img_reg_array_54_31_imag;
        _zz_304 = img_reg_array_55_31_real;
        _zz_305 = img_reg_array_55_31_imag;
        _zz_306 = img_reg_array_56_31_real;
        _zz_307 = img_reg_array_56_31_imag;
        _zz_308 = img_reg_array_57_31_real;
        _zz_309 = img_reg_array_57_31_imag;
        _zz_310 = img_reg_array_58_31_real;
        _zz_311 = img_reg_array_58_31_imag;
        _zz_312 = img_reg_array_59_31_real;
        _zz_313 = img_reg_array_59_31_imag;
        _zz_314 = img_reg_array_60_31_real;
        _zz_315 = img_reg_array_60_31_imag;
        _zz_316 = img_reg_array_61_31_real;
        _zz_317 = img_reg_array_61_31_imag;
        _zz_318 = img_reg_array_62_31_real;
        _zz_319 = img_reg_array_62_31_imag;
        _zz_320 = img_reg_array_63_31_real;
        _zz_321 = img_reg_array_63_31_imag;
      end
      6'b100000 : begin
        _zz_194 = img_reg_array_0_32_real;
        _zz_195 = img_reg_array_0_32_imag;
        _zz_196 = img_reg_array_1_32_real;
        _zz_197 = img_reg_array_1_32_imag;
        _zz_198 = img_reg_array_2_32_real;
        _zz_199 = img_reg_array_2_32_imag;
        _zz_200 = img_reg_array_3_32_real;
        _zz_201 = img_reg_array_3_32_imag;
        _zz_202 = img_reg_array_4_32_real;
        _zz_203 = img_reg_array_4_32_imag;
        _zz_204 = img_reg_array_5_32_real;
        _zz_205 = img_reg_array_5_32_imag;
        _zz_206 = img_reg_array_6_32_real;
        _zz_207 = img_reg_array_6_32_imag;
        _zz_208 = img_reg_array_7_32_real;
        _zz_209 = img_reg_array_7_32_imag;
        _zz_210 = img_reg_array_8_32_real;
        _zz_211 = img_reg_array_8_32_imag;
        _zz_212 = img_reg_array_9_32_real;
        _zz_213 = img_reg_array_9_32_imag;
        _zz_214 = img_reg_array_10_32_real;
        _zz_215 = img_reg_array_10_32_imag;
        _zz_216 = img_reg_array_11_32_real;
        _zz_217 = img_reg_array_11_32_imag;
        _zz_218 = img_reg_array_12_32_real;
        _zz_219 = img_reg_array_12_32_imag;
        _zz_220 = img_reg_array_13_32_real;
        _zz_221 = img_reg_array_13_32_imag;
        _zz_222 = img_reg_array_14_32_real;
        _zz_223 = img_reg_array_14_32_imag;
        _zz_224 = img_reg_array_15_32_real;
        _zz_225 = img_reg_array_15_32_imag;
        _zz_226 = img_reg_array_16_32_real;
        _zz_227 = img_reg_array_16_32_imag;
        _zz_228 = img_reg_array_17_32_real;
        _zz_229 = img_reg_array_17_32_imag;
        _zz_230 = img_reg_array_18_32_real;
        _zz_231 = img_reg_array_18_32_imag;
        _zz_232 = img_reg_array_19_32_real;
        _zz_233 = img_reg_array_19_32_imag;
        _zz_234 = img_reg_array_20_32_real;
        _zz_235 = img_reg_array_20_32_imag;
        _zz_236 = img_reg_array_21_32_real;
        _zz_237 = img_reg_array_21_32_imag;
        _zz_238 = img_reg_array_22_32_real;
        _zz_239 = img_reg_array_22_32_imag;
        _zz_240 = img_reg_array_23_32_real;
        _zz_241 = img_reg_array_23_32_imag;
        _zz_242 = img_reg_array_24_32_real;
        _zz_243 = img_reg_array_24_32_imag;
        _zz_244 = img_reg_array_25_32_real;
        _zz_245 = img_reg_array_25_32_imag;
        _zz_246 = img_reg_array_26_32_real;
        _zz_247 = img_reg_array_26_32_imag;
        _zz_248 = img_reg_array_27_32_real;
        _zz_249 = img_reg_array_27_32_imag;
        _zz_250 = img_reg_array_28_32_real;
        _zz_251 = img_reg_array_28_32_imag;
        _zz_252 = img_reg_array_29_32_real;
        _zz_253 = img_reg_array_29_32_imag;
        _zz_254 = img_reg_array_30_32_real;
        _zz_255 = img_reg_array_30_32_imag;
        _zz_256 = img_reg_array_31_32_real;
        _zz_257 = img_reg_array_31_32_imag;
        _zz_258 = img_reg_array_32_32_real;
        _zz_259 = img_reg_array_32_32_imag;
        _zz_260 = img_reg_array_33_32_real;
        _zz_261 = img_reg_array_33_32_imag;
        _zz_262 = img_reg_array_34_32_real;
        _zz_263 = img_reg_array_34_32_imag;
        _zz_264 = img_reg_array_35_32_real;
        _zz_265 = img_reg_array_35_32_imag;
        _zz_266 = img_reg_array_36_32_real;
        _zz_267 = img_reg_array_36_32_imag;
        _zz_268 = img_reg_array_37_32_real;
        _zz_269 = img_reg_array_37_32_imag;
        _zz_270 = img_reg_array_38_32_real;
        _zz_271 = img_reg_array_38_32_imag;
        _zz_272 = img_reg_array_39_32_real;
        _zz_273 = img_reg_array_39_32_imag;
        _zz_274 = img_reg_array_40_32_real;
        _zz_275 = img_reg_array_40_32_imag;
        _zz_276 = img_reg_array_41_32_real;
        _zz_277 = img_reg_array_41_32_imag;
        _zz_278 = img_reg_array_42_32_real;
        _zz_279 = img_reg_array_42_32_imag;
        _zz_280 = img_reg_array_43_32_real;
        _zz_281 = img_reg_array_43_32_imag;
        _zz_282 = img_reg_array_44_32_real;
        _zz_283 = img_reg_array_44_32_imag;
        _zz_284 = img_reg_array_45_32_real;
        _zz_285 = img_reg_array_45_32_imag;
        _zz_286 = img_reg_array_46_32_real;
        _zz_287 = img_reg_array_46_32_imag;
        _zz_288 = img_reg_array_47_32_real;
        _zz_289 = img_reg_array_47_32_imag;
        _zz_290 = img_reg_array_48_32_real;
        _zz_291 = img_reg_array_48_32_imag;
        _zz_292 = img_reg_array_49_32_real;
        _zz_293 = img_reg_array_49_32_imag;
        _zz_294 = img_reg_array_50_32_real;
        _zz_295 = img_reg_array_50_32_imag;
        _zz_296 = img_reg_array_51_32_real;
        _zz_297 = img_reg_array_51_32_imag;
        _zz_298 = img_reg_array_52_32_real;
        _zz_299 = img_reg_array_52_32_imag;
        _zz_300 = img_reg_array_53_32_real;
        _zz_301 = img_reg_array_53_32_imag;
        _zz_302 = img_reg_array_54_32_real;
        _zz_303 = img_reg_array_54_32_imag;
        _zz_304 = img_reg_array_55_32_real;
        _zz_305 = img_reg_array_55_32_imag;
        _zz_306 = img_reg_array_56_32_real;
        _zz_307 = img_reg_array_56_32_imag;
        _zz_308 = img_reg_array_57_32_real;
        _zz_309 = img_reg_array_57_32_imag;
        _zz_310 = img_reg_array_58_32_real;
        _zz_311 = img_reg_array_58_32_imag;
        _zz_312 = img_reg_array_59_32_real;
        _zz_313 = img_reg_array_59_32_imag;
        _zz_314 = img_reg_array_60_32_real;
        _zz_315 = img_reg_array_60_32_imag;
        _zz_316 = img_reg_array_61_32_real;
        _zz_317 = img_reg_array_61_32_imag;
        _zz_318 = img_reg_array_62_32_real;
        _zz_319 = img_reg_array_62_32_imag;
        _zz_320 = img_reg_array_63_32_real;
        _zz_321 = img_reg_array_63_32_imag;
      end
      6'b100001 : begin
        _zz_194 = img_reg_array_0_33_real;
        _zz_195 = img_reg_array_0_33_imag;
        _zz_196 = img_reg_array_1_33_real;
        _zz_197 = img_reg_array_1_33_imag;
        _zz_198 = img_reg_array_2_33_real;
        _zz_199 = img_reg_array_2_33_imag;
        _zz_200 = img_reg_array_3_33_real;
        _zz_201 = img_reg_array_3_33_imag;
        _zz_202 = img_reg_array_4_33_real;
        _zz_203 = img_reg_array_4_33_imag;
        _zz_204 = img_reg_array_5_33_real;
        _zz_205 = img_reg_array_5_33_imag;
        _zz_206 = img_reg_array_6_33_real;
        _zz_207 = img_reg_array_6_33_imag;
        _zz_208 = img_reg_array_7_33_real;
        _zz_209 = img_reg_array_7_33_imag;
        _zz_210 = img_reg_array_8_33_real;
        _zz_211 = img_reg_array_8_33_imag;
        _zz_212 = img_reg_array_9_33_real;
        _zz_213 = img_reg_array_9_33_imag;
        _zz_214 = img_reg_array_10_33_real;
        _zz_215 = img_reg_array_10_33_imag;
        _zz_216 = img_reg_array_11_33_real;
        _zz_217 = img_reg_array_11_33_imag;
        _zz_218 = img_reg_array_12_33_real;
        _zz_219 = img_reg_array_12_33_imag;
        _zz_220 = img_reg_array_13_33_real;
        _zz_221 = img_reg_array_13_33_imag;
        _zz_222 = img_reg_array_14_33_real;
        _zz_223 = img_reg_array_14_33_imag;
        _zz_224 = img_reg_array_15_33_real;
        _zz_225 = img_reg_array_15_33_imag;
        _zz_226 = img_reg_array_16_33_real;
        _zz_227 = img_reg_array_16_33_imag;
        _zz_228 = img_reg_array_17_33_real;
        _zz_229 = img_reg_array_17_33_imag;
        _zz_230 = img_reg_array_18_33_real;
        _zz_231 = img_reg_array_18_33_imag;
        _zz_232 = img_reg_array_19_33_real;
        _zz_233 = img_reg_array_19_33_imag;
        _zz_234 = img_reg_array_20_33_real;
        _zz_235 = img_reg_array_20_33_imag;
        _zz_236 = img_reg_array_21_33_real;
        _zz_237 = img_reg_array_21_33_imag;
        _zz_238 = img_reg_array_22_33_real;
        _zz_239 = img_reg_array_22_33_imag;
        _zz_240 = img_reg_array_23_33_real;
        _zz_241 = img_reg_array_23_33_imag;
        _zz_242 = img_reg_array_24_33_real;
        _zz_243 = img_reg_array_24_33_imag;
        _zz_244 = img_reg_array_25_33_real;
        _zz_245 = img_reg_array_25_33_imag;
        _zz_246 = img_reg_array_26_33_real;
        _zz_247 = img_reg_array_26_33_imag;
        _zz_248 = img_reg_array_27_33_real;
        _zz_249 = img_reg_array_27_33_imag;
        _zz_250 = img_reg_array_28_33_real;
        _zz_251 = img_reg_array_28_33_imag;
        _zz_252 = img_reg_array_29_33_real;
        _zz_253 = img_reg_array_29_33_imag;
        _zz_254 = img_reg_array_30_33_real;
        _zz_255 = img_reg_array_30_33_imag;
        _zz_256 = img_reg_array_31_33_real;
        _zz_257 = img_reg_array_31_33_imag;
        _zz_258 = img_reg_array_32_33_real;
        _zz_259 = img_reg_array_32_33_imag;
        _zz_260 = img_reg_array_33_33_real;
        _zz_261 = img_reg_array_33_33_imag;
        _zz_262 = img_reg_array_34_33_real;
        _zz_263 = img_reg_array_34_33_imag;
        _zz_264 = img_reg_array_35_33_real;
        _zz_265 = img_reg_array_35_33_imag;
        _zz_266 = img_reg_array_36_33_real;
        _zz_267 = img_reg_array_36_33_imag;
        _zz_268 = img_reg_array_37_33_real;
        _zz_269 = img_reg_array_37_33_imag;
        _zz_270 = img_reg_array_38_33_real;
        _zz_271 = img_reg_array_38_33_imag;
        _zz_272 = img_reg_array_39_33_real;
        _zz_273 = img_reg_array_39_33_imag;
        _zz_274 = img_reg_array_40_33_real;
        _zz_275 = img_reg_array_40_33_imag;
        _zz_276 = img_reg_array_41_33_real;
        _zz_277 = img_reg_array_41_33_imag;
        _zz_278 = img_reg_array_42_33_real;
        _zz_279 = img_reg_array_42_33_imag;
        _zz_280 = img_reg_array_43_33_real;
        _zz_281 = img_reg_array_43_33_imag;
        _zz_282 = img_reg_array_44_33_real;
        _zz_283 = img_reg_array_44_33_imag;
        _zz_284 = img_reg_array_45_33_real;
        _zz_285 = img_reg_array_45_33_imag;
        _zz_286 = img_reg_array_46_33_real;
        _zz_287 = img_reg_array_46_33_imag;
        _zz_288 = img_reg_array_47_33_real;
        _zz_289 = img_reg_array_47_33_imag;
        _zz_290 = img_reg_array_48_33_real;
        _zz_291 = img_reg_array_48_33_imag;
        _zz_292 = img_reg_array_49_33_real;
        _zz_293 = img_reg_array_49_33_imag;
        _zz_294 = img_reg_array_50_33_real;
        _zz_295 = img_reg_array_50_33_imag;
        _zz_296 = img_reg_array_51_33_real;
        _zz_297 = img_reg_array_51_33_imag;
        _zz_298 = img_reg_array_52_33_real;
        _zz_299 = img_reg_array_52_33_imag;
        _zz_300 = img_reg_array_53_33_real;
        _zz_301 = img_reg_array_53_33_imag;
        _zz_302 = img_reg_array_54_33_real;
        _zz_303 = img_reg_array_54_33_imag;
        _zz_304 = img_reg_array_55_33_real;
        _zz_305 = img_reg_array_55_33_imag;
        _zz_306 = img_reg_array_56_33_real;
        _zz_307 = img_reg_array_56_33_imag;
        _zz_308 = img_reg_array_57_33_real;
        _zz_309 = img_reg_array_57_33_imag;
        _zz_310 = img_reg_array_58_33_real;
        _zz_311 = img_reg_array_58_33_imag;
        _zz_312 = img_reg_array_59_33_real;
        _zz_313 = img_reg_array_59_33_imag;
        _zz_314 = img_reg_array_60_33_real;
        _zz_315 = img_reg_array_60_33_imag;
        _zz_316 = img_reg_array_61_33_real;
        _zz_317 = img_reg_array_61_33_imag;
        _zz_318 = img_reg_array_62_33_real;
        _zz_319 = img_reg_array_62_33_imag;
        _zz_320 = img_reg_array_63_33_real;
        _zz_321 = img_reg_array_63_33_imag;
      end
      6'b100010 : begin
        _zz_194 = img_reg_array_0_34_real;
        _zz_195 = img_reg_array_0_34_imag;
        _zz_196 = img_reg_array_1_34_real;
        _zz_197 = img_reg_array_1_34_imag;
        _zz_198 = img_reg_array_2_34_real;
        _zz_199 = img_reg_array_2_34_imag;
        _zz_200 = img_reg_array_3_34_real;
        _zz_201 = img_reg_array_3_34_imag;
        _zz_202 = img_reg_array_4_34_real;
        _zz_203 = img_reg_array_4_34_imag;
        _zz_204 = img_reg_array_5_34_real;
        _zz_205 = img_reg_array_5_34_imag;
        _zz_206 = img_reg_array_6_34_real;
        _zz_207 = img_reg_array_6_34_imag;
        _zz_208 = img_reg_array_7_34_real;
        _zz_209 = img_reg_array_7_34_imag;
        _zz_210 = img_reg_array_8_34_real;
        _zz_211 = img_reg_array_8_34_imag;
        _zz_212 = img_reg_array_9_34_real;
        _zz_213 = img_reg_array_9_34_imag;
        _zz_214 = img_reg_array_10_34_real;
        _zz_215 = img_reg_array_10_34_imag;
        _zz_216 = img_reg_array_11_34_real;
        _zz_217 = img_reg_array_11_34_imag;
        _zz_218 = img_reg_array_12_34_real;
        _zz_219 = img_reg_array_12_34_imag;
        _zz_220 = img_reg_array_13_34_real;
        _zz_221 = img_reg_array_13_34_imag;
        _zz_222 = img_reg_array_14_34_real;
        _zz_223 = img_reg_array_14_34_imag;
        _zz_224 = img_reg_array_15_34_real;
        _zz_225 = img_reg_array_15_34_imag;
        _zz_226 = img_reg_array_16_34_real;
        _zz_227 = img_reg_array_16_34_imag;
        _zz_228 = img_reg_array_17_34_real;
        _zz_229 = img_reg_array_17_34_imag;
        _zz_230 = img_reg_array_18_34_real;
        _zz_231 = img_reg_array_18_34_imag;
        _zz_232 = img_reg_array_19_34_real;
        _zz_233 = img_reg_array_19_34_imag;
        _zz_234 = img_reg_array_20_34_real;
        _zz_235 = img_reg_array_20_34_imag;
        _zz_236 = img_reg_array_21_34_real;
        _zz_237 = img_reg_array_21_34_imag;
        _zz_238 = img_reg_array_22_34_real;
        _zz_239 = img_reg_array_22_34_imag;
        _zz_240 = img_reg_array_23_34_real;
        _zz_241 = img_reg_array_23_34_imag;
        _zz_242 = img_reg_array_24_34_real;
        _zz_243 = img_reg_array_24_34_imag;
        _zz_244 = img_reg_array_25_34_real;
        _zz_245 = img_reg_array_25_34_imag;
        _zz_246 = img_reg_array_26_34_real;
        _zz_247 = img_reg_array_26_34_imag;
        _zz_248 = img_reg_array_27_34_real;
        _zz_249 = img_reg_array_27_34_imag;
        _zz_250 = img_reg_array_28_34_real;
        _zz_251 = img_reg_array_28_34_imag;
        _zz_252 = img_reg_array_29_34_real;
        _zz_253 = img_reg_array_29_34_imag;
        _zz_254 = img_reg_array_30_34_real;
        _zz_255 = img_reg_array_30_34_imag;
        _zz_256 = img_reg_array_31_34_real;
        _zz_257 = img_reg_array_31_34_imag;
        _zz_258 = img_reg_array_32_34_real;
        _zz_259 = img_reg_array_32_34_imag;
        _zz_260 = img_reg_array_33_34_real;
        _zz_261 = img_reg_array_33_34_imag;
        _zz_262 = img_reg_array_34_34_real;
        _zz_263 = img_reg_array_34_34_imag;
        _zz_264 = img_reg_array_35_34_real;
        _zz_265 = img_reg_array_35_34_imag;
        _zz_266 = img_reg_array_36_34_real;
        _zz_267 = img_reg_array_36_34_imag;
        _zz_268 = img_reg_array_37_34_real;
        _zz_269 = img_reg_array_37_34_imag;
        _zz_270 = img_reg_array_38_34_real;
        _zz_271 = img_reg_array_38_34_imag;
        _zz_272 = img_reg_array_39_34_real;
        _zz_273 = img_reg_array_39_34_imag;
        _zz_274 = img_reg_array_40_34_real;
        _zz_275 = img_reg_array_40_34_imag;
        _zz_276 = img_reg_array_41_34_real;
        _zz_277 = img_reg_array_41_34_imag;
        _zz_278 = img_reg_array_42_34_real;
        _zz_279 = img_reg_array_42_34_imag;
        _zz_280 = img_reg_array_43_34_real;
        _zz_281 = img_reg_array_43_34_imag;
        _zz_282 = img_reg_array_44_34_real;
        _zz_283 = img_reg_array_44_34_imag;
        _zz_284 = img_reg_array_45_34_real;
        _zz_285 = img_reg_array_45_34_imag;
        _zz_286 = img_reg_array_46_34_real;
        _zz_287 = img_reg_array_46_34_imag;
        _zz_288 = img_reg_array_47_34_real;
        _zz_289 = img_reg_array_47_34_imag;
        _zz_290 = img_reg_array_48_34_real;
        _zz_291 = img_reg_array_48_34_imag;
        _zz_292 = img_reg_array_49_34_real;
        _zz_293 = img_reg_array_49_34_imag;
        _zz_294 = img_reg_array_50_34_real;
        _zz_295 = img_reg_array_50_34_imag;
        _zz_296 = img_reg_array_51_34_real;
        _zz_297 = img_reg_array_51_34_imag;
        _zz_298 = img_reg_array_52_34_real;
        _zz_299 = img_reg_array_52_34_imag;
        _zz_300 = img_reg_array_53_34_real;
        _zz_301 = img_reg_array_53_34_imag;
        _zz_302 = img_reg_array_54_34_real;
        _zz_303 = img_reg_array_54_34_imag;
        _zz_304 = img_reg_array_55_34_real;
        _zz_305 = img_reg_array_55_34_imag;
        _zz_306 = img_reg_array_56_34_real;
        _zz_307 = img_reg_array_56_34_imag;
        _zz_308 = img_reg_array_57_34_real;
        _zz_309 = img_reg_array_57_34_imag;
        _zz_310 = img_reg_array_58_34_real;
        _zz_311 = img_reg_array_58_34_imag;
        _zz_312 = img_reg_array_59_34_real;
        _zz_313 = img_reg_array_59_34_imag;
        _zz_314 = img_reg_array_60_34_real;
        _zz_315 = img_reg_array_60_34_imag;
        _zz_316 = img_reg_array_61_34_real;
        _zz_317 = img_reg_array_61_34_imag;
        _zz_318 = img_reg_array_62_34_real;
        _zz_319 = img_reg_array_62_34_imag;
        _zz_320 = img_reg_array_63_34_real;
        _zz_321 = img_reg_array_63_34_imag;
      end
      6'b100011 : begin
        _zz_194 = img_reg_array_0_35_real;
        _zz_195 = img_reg_array_0_35_imag;
        _zz_196 = img_reg_array_1_35_real;
        _zz_197 = img_reg_array_1_35_imag;
        _zz_198 = img_reg_array_2_35_real;
        _zz_199 = img_reg_array_2_35_imag;
        _zz_200 = img_reg_array_3_35_real;
        _zz_201 = img_reg_array_3_35_imag;
        _zz_202 = img_reg_array_4_35_real;
        _zz_203 = img_reg_array_4_35_imag;
        _zz_204 = img_reg_array_5_35_real;
        _zz_205 = img_reg_array_5_35_imag;
        _zz_206 = img_reg_array_6_35_real;
        _zz_207 = img_reg_array_6_35_imag;
        _zz_208 = img_reg_array_7_35_real;
        _zz_209 = img_reg_array_7_35_imag;
        _zz_210 = img_reg_array_8_35_real;
        _zz_211 = img_reg_array_8_35_imag;
        _zz_212 = img_reg_array_9_35_real;
        _zz_213 = img_reg_array_9_35_imag;
        _zz_214 = img_reg_array_10_35_real;
        _zz_215 = img_reg_array_10_35_imag;
        _zz_216 = img_reg_array_11_35_real;
        _zz_217 = img_reg_array_11_35_imag;
        _zz_218 = img_reg_array_12_35_real;
        _zz_219 = img_reg_array_12_35_imag;
        _zz_220 = img_reg_array_13_35_real;
        _zz_221 = img_reg_array_13_35_imag;
        _zz_222 = img_reg_array_14_35_real;
        _zz_223 = img_reg_array_14_35_imag;
        _zz_224 = img_reg_array_15_35_real;
        _zz_225 = img_reg_array_15_35_imag;
        _zz_226 = img_reg_array_16_35_real;
        _zz_227 = img_reg_array_16_35_imag;
        _zz_228 = img_reg_array_17_35_real;
        _zz_229 = img_reg_array_17_35_imag;
        _zz_230 = img_reg_array_18_35_real;
        _zz_231 = img_reg_array_18_35_imag;
        _zz_232 = img_reg_array_19_35_real;
        _zz_233 = img_reg_array_19_35_imag;
        _zz_234 = img_reg_array_20_35_real;
        _zz_235 = img_reg_array_20_35_imag;
        _zz_236 = img_reg_array_21_35_real;
        _zz_237 = img_reg_array_21_35_imag;
        _zz_238 = img_reg_array_22_35_real;
        _zz_239 = img_reg_array_22_35_imag;
        _zz_240 = img_reg_array_23_35_real;
        _zz_241 = img_reg_array_23_35_imag;
        _zz_242 = img_reg_array_24_35_real;
        _zz_243 = img_reg_array_24_35_imag;
        _zz_244 = img_reg_array_25_35_real;
        _zz_245 = img_reg_array_25_35_imag;
        _zz_246 = img_reg_array_26_35_real;
        _zz_247 = img_reg_array_26_35_imag;
        _zz_248 = img_reg_array_27_35_real;
        _zz_249 = img_reg_array_27_35_imag;
        _zz_250 = img_reg_array_28_35_real;
        _zz_251 = img_reg_array_28_35_imag;
        _zz_252 = img_reg_array_29_35_real;
        _zz_253 = img_reg_array_29_35_imag;
        _zz_254 = img_reg_array_30_35_real;
        _zz_255 = img_reg_array_30_35_imag;
        _zz_256 = img_reg_array_31_35_real;
        _zz_257 = img_reg_array_31_35_imag;
        _zz_258 = img_reg_array_32_35_real;
        _zz_259 = img_reg_array_32_35_imag;
        _zz_260 = img_reg_array_33_35_real;
        _zz_261 = img_reg_array_33_35_imag;
        _zz_262 = img_reg_array_34_35_real;
        _zz_263 = img_reg_array_34_35_imag;
        _zz_264 = img_reg_array_35_35_real;
        _zz_265 = img_reg_array_35_35_imag;
        _zz_266 = img_reg_array_36_35_real;
        _zz_267 = img_reg_array_36_35_imag;
        _zz_268 = img_reg_array_37_35_real;
        _zz_269 = img_reg_array_37_35_imag;
        _zz_270 = img_reg_array_38_35_real;
        _zz_271 = img_reg_array_38_35_imag;
        _zz_272 = img_reg_array_39_35_real;
        _zz_273 = img_reg_array_39_35_imag;
        _zz_274 = img_reg_array_40_35_real;
        _zz_275 = img_reg_array_40_35_imag;
        _zz_276 = img_reg_array_41_35_real;
        _zz_277 = img_reg_array_41_35_imag;
        _zz_278 = img_reg_array_42_35_real;
        _zz_279 = img_reg_array_42_35_imag;
        _zz_280 = img_reg_array_43_35_real;
        _zz_281 = img_reg_array_43_35_imag;
        _zz_282 = img_reg_array_44_35_real;
        _zz_283 = img_reg_array_44_35_imag;
        _zz_284 = img_reg_array_45_35_real;
        _zz_285 = img_reg_array_45_35_imag;
        _zz_286 = img_reg_array_46_35_real;
        _zz_287 = img_reg_array_46_35_imag;
        _zz_288 = img_reg_array_47_35_real;
        _zz_289 = img_reg_array_47_35_imag;
        _zz_290 = img_reg_array_48_35_real;
        _zz_291 = img_reg_array_48_35_imag;
        _zz_292 = img_reg_array_49_35_real;
        _zz_293 = img_reg_array_49_35_imag;
        _zz_294 = img_reg_array_50_35_real;
        _zz_295 = img_reg_array_50_35_imag;
        _zz_296 = img_reg_array_51_35_real;
        _zz_297 = img_reg_array_51_35_imag;
        _zz_298 = img_reg_array_52_35_real;
        _zz_299 = img_reg_array_52_35_imag;
        _zz_300 = img_reg_array_53_35_real;
        _zz_301 = img_reg_array_53_35_imag;
        _zz_302 = img_reg_array_54_35_real;
        _zz_303 = img_reg_array_54_35_imag;
        _zz_304 = img_reg_array_55_35_real;
        _zz_305 = img_reg_array_55_35_imag;
        _zz_306 = img_reg_array_56_35_real;
        _zz_307 = img_reg_array_56_35_imag;
        _zz_308 = img_reg_array_57_35_real;
        _zz_309 = img_reg_array_57_35_imag;
        _zz_310 = img_reg_array_58_35_real;
        _zz_311 = img_reg_array_58_35_imag;
        _zz_312 = img_reg_array_59_35_real;
        _zz_313 = img_reg_array_59_35_imag;
        _zz_314 = img_reg_array_60_35_real;
        _zz_315 = img_reg_array_60_35_imag;
        _zz_316 = img_reg_array_61_35_real;
        _zz_317 = img_reg_array_61_35_imag;
        _zz_318 = img_reg_array_62_35_real;
        _zz_319 = img_reg_array_62_35_imag;
        _zz_320 = img_reg_array_63_35_real;
        _zz_321 = img_reg_array_63_35_imag;
      end
      6'b100100 : begin
        _zz_194 = img_reg_array_0_36_real;
        _zz_195 = img_reg_array_0_36_imag;
        _zz_196 = img_reg_array_1_36_real;
        _zz_197 = img_reg_array_1_36_imag;
        _zz_198 = img_reg_array_2_36_real;
        _zz_199 = img_reg_array_2_36_imag;
        _zz_200 = img_reg_array_3_36_real;
        _zz_201 = img_reg_array_3_36_imag;
        _zz_202 = img_reg_array_4_36_real;
        _zz_203 = img_reg_array_4_36_imag;
        _zz_204 = img_reg_array_5_36_real;
        _zz_205 = img_reg_array_5_36_imag;
        _zz_206 = img_reg_array_6_36_real;
        _zz_207 = img_reg_array_6_36_imag;
        _zz_208 = img_reg_array_7_36_real;
        _zz_209 = img_reg_array_7_36_imag;
        _zz_210 = img_reg_array_8_36_real;
        _zz_211 = img_reg_array_8_36_imag;
        _zz_212 = img_reg_array_9_36_real;
        _zz_213 = img_reg_array_9_36_imag;
        _zz_214 = img_reg_array_10_36_real;
        _zz_215 = img_reg_array_10_36_imag;
        _zz_216 = img_reg_array_11_36_real;
        _zz_217 = img_reg_array_11_36_imag;
        _zz_218 = img_reg_array_12_36_real;
        _zz_219 = img_reg_array_12_36_imag;
        _zz_220 = img_reg_array_13_36_real;
        _zz_221 = img_reg_array_13_36_imag;
        _zz_222 = img_reg_array_14_36_real;
        _zz_223 = img_reg_array_14_36_imag;
        _zz_224 = img_reg_array_15_36_real;
        _zz_225 = img_reg_array_15_36_imag;
        _zz_226 = img_reg_array_16_36_real;
        _zz_227 = img_reg_array_16_36_imag;
        _zz_228 = img_reg_array_17_36_real;
        _zz_229 = img_reg_array_17_36_imag;
        _zz_230 = img_reg_array_18_36_real;
        _zz_231 = img_reg_array_18_36_imag;
        _zz_232 = img_reg_array_19_36_real;
        _zz_233 = img_reg_array_19_36_imag;
        _zz_234 = img_reg_array_20_36_real;
        _zz_235 = img_reg_array_20_36_imag;
        _zz_236 = img_reg_array_21_36_real;
        _zz_237 = img_reg_array_21_36_imag;
        _zz_238 = img_reg_array_22_36_real;
        _zz_239 = img_reg_array_22_36_imag;
        _zz_240 = img_reg_array_23_36_real;
        _zz_241 = img_reg_array_23_36_imag;
        _zz_242 = img_reg_array_24_36_real;
        _zz_243 = img_reg_array_24_36_imag;
        _zz_244 = img_reg_array_25_36_real;
        _zz_245 = img_reg_array_25_36_imag;
        _zz_246 = img_reg_array_26_36_real;
        _zz_247 = img_reg_array_26_36_imag;
        _zz_248 = img_reg_array_27_36_real;
        _zz_249 = img_reg_array_27_36_imag;
        _zz_250 = img_reg_array_28_36_real;
        _zz_251 = img_reg_array_28_36_imag;
        _zz_252 = img_reg_array_29_36_real;
        _zz_253 = img_reg_array_29_36_imag;
        _zz_254 = img_reg_array_30_36_real;
        _zz_255 = img_reg_array_30_36_imag;
        _zz_256 = img_reg_array_31_36_real;
        _zz_257 = img_reg_array_31_36_imag;
        _zz_258 = img_reg_array_32_36_real;
        _zz_259 = img_reg_array_32_36_imag;
        _zz_260 = img_reg_array_33_36_real;
        _zz_261 = img_reg_array_33_36_imag;
        _zz_262 = img_reg_array_34_36_real;
        _zz_263 = img_reg_array_34_36_imag;
        _zz_264 = img_reg_array_35_36_real;
        _zz_265 = img_reg_array_35_36_imag;
        _zz_266 = img_reg_array_36_36_real;
        _zz_267 = img_reg_array_36_36_imag;
        _zz_268 = img_reg_array_37_36_real;
        _zz_269 = img_reg_array_37_36_imag;
        _zz_270 = img_reg_array_38_36_real;
        _zz_271 = img_reg_array_38_36_imag;
        _zz_272 = img_reg_array_39_36_real;
        _zz_273 = img_reg_array_39_36_imag;
        _zz_274 = img_reg_array_40_36_real;
        _zz_275 = img_reg_array_40_36_imag;
        _zz_276 = img_reg_array_41_36_real;
        _zz_277 = img_reg_array_41_36_imag;
        _zz_278 = img_reg_array_42_36_real;
        _zz_279 = img_reg_array_42_36_imag;
        _zz_280 = img_reg_array_43_36_real;
        _zz_281 = img_reg_array_43_36_imag;
        _zz_282 = img_reg_array_44_36_real;
        _zz_283 = img_reg_array_44_36_imag;
        _zz_284 = img_reg_array_45_36_real;
        _zz_285 = img_reg_array_45_36_imag;
        _zz_286 = img_reg_array_46_36_real;
        _zz_287 = img_reg_array_46_36_imag;
        _zz_288 = img_reg_array_47_36_real;
        _zz_289 = img_reg_array_47_36_imag;
        _zz_290 = img_reg_array_48_36_real;
        _zz_291 = img_reg_array_48_36_imag;
        _zz_292 = img_reg_array_49_36_real;
        _zz_293 = img_reg_array_49_36_imag;
        _zz_294 = img_reg_array_50_36_real;
        _zz_295 = img_reg_array_50_36_imag;
        _zz_296 = img_reg_array_51_36_real;
        _zz_297 = img_reg_array_51_36_imag;
        _zz_298 = img_reg_array_52_36_real;
        _zz_299 = img_reg_array_52_36_imag;
        _zz_300 = img_reg_array_53_36_real;
        _zz_301 = img_reg_array_53_36_imag;
        _zz_302 = img_reg_array_54_36_real;
        _zz_303 = img_reg_array_54_36_imag;
        _zz_304 = img_reg_array_55_36_real;
        _zz_305 = img_reg_array_55_36_imag;
        _zz_306 = img_reg_array_56_36_real;
        _zz_307 = img_reg_array_56_36_imag;
        _zz_308 = img_reg_array_57_36_real;
        _zz_309 = img_reg_array_57_36_imag;
        _zz_310 = img_reg_array_58_36_real;
        _zz_311 = img_reg_array_58_36_imag;
        _zz_312 = img_reg_array_59_36_real;
        _zz_313 = img_reg_array_59_36_imag;
        _zz_314 = img_reg_array_60_36_real;
        _zz_315 = img_reg_array_60_36_imag;
        _zz_316 = img_reg_array_61_36_real;
        _zz_317 = img_reg_array_61_36_imag;
        _zz_318 = img_reg_array_62_36_real;
        _zz_319 = img_reg_array_62_36_imag;
        _zz_320 = img_reg_array_63_36_real;
        _zz_321 = img_reg_array_63_36_imag;
      end
      6'b100101 : begin
        _zz_194 = img_reg_array_0_37_real;
        _zz_195 = img_reg_array_0_37_imag;
        _zz_196 = img_reg_array_1_37_real;
        _zz_197 = img_reg_array_1_37_imag;
        _zz_198 = img_reg_array_2_37_real;
        _zz_199 = img_reg_array_2_37_imag;
        _zz_200 = img_reg_array_3_37_real;
        _zz_201 = img_reg_array_3_37_imag;
        _zz_202 = img_reg_array_4_37_real;
        _zz_203 = img_reg_array_4_37_imag;
        _zz_204 = img_reg_array_5_37_real;
        _zz_205 = img_reg_array_5_37_imag;
        _zz_206 = img_reg_array_6_37_real;
        _zz_207 = img_reg_array_6_37_imag;
        _zz_208 = img_reg_array_7_37_real;
        _zz_209 = img_reg_array_7_37_imag;
        _zz_210 = img_reg_array_8_37_real;
        _zz_211 = img_reg_array_8_37_imag;
        _zz_212 = img_reg_array_9_37_real;
        _zz_213 = img_reg_array_9_37_imag;
        _zz_214 = img_reg_array_10_37_real;
        _zz_215 = img_reg_array_10_37_imag;
        _zz_216 = img_reg_array_11_37_real;
        _zz_217 = img_reg_array_11_37_imag;
        _zz_218 = img_reg_array_12_37_real;
        _zz_219 = img_reg_array_12_37_imag;
        _zz_220 = img_reg_array_13_37_real;
        _zz_221 = img_reg_array_13_37_imag;
        _zz_222 = img_reg_array_14_37_real;
        _zz_223 = img_reg_array_14_37_imag;
        _zz_224 = img_reg_array_15_37_real;
        _zz_225 = img_reg_array_15_37_imag;
        _zz_226 = img_reg_array_16_37_real;
        _zz_227 = img_reg_array_16_37_imag;
        _zz_228 = img_reg_array_17_37_real;
        _zz_229 = img_reg_array_17_37_imag;
        _zz_230 = img_reg_array_18_37_real;
        _zz_231 = img_reg_array_18_37_imag;
        _zz_232 = img_reg_array_19_37_real;
        _zz_233 = img_reg_array_19_37_imag;
        _zz_234 = img_reg_array_20_37_real;
        _zz_235 = img_reg_array_20_37_imag;
        _zz_236 = img_reg_array_21_37_real;
        _zz_237 = img_reg_array_21_37_imag;
        _zz_238 = img_reg_array_22_37_real;
        _zz_239 = img_reg_array_22_37_imag;
        _zz_240 = img_reg_array_23_37_real;
        _zz_241 = img_reg_array_23_37_imag;
        _zz_242 = img_reg_array_24_37_real;
        _zz_243 = img_reg_array_24_37_imag;
        _zz_244 = img_reg_array_25_37_real;
        _zz_245 = img_reg_array_25_37_imag;
        _zz_246 = img_reg_array_26_37_real;
        _zz_247 = img_reg_array_26_37_imag;
        _zz_248 = img_reg_array_27_37_real;
        _zz_249 = img_reg_array_27_37_imag;
        _zz_250 = img_reg_array_28_37_real;
        _zz_251 = img_reg_array_28_37_imag;
        _zz_252 = img_reg_array_29_37_real;
        _zz_253 = img_reg_array_29_37_imag;
        _zz_254 = img_reg_array_30_37_real;
        _zz_255 = img_reg_array_30_37_imag;
        _zz_256 = img_reg_array_31_37_real;
        _zz_257 = img_reg_array_31_37_imag;
        _zz_258 = img_reg_array_32_37_real;
        _zz_259 = img_reg_array_32_37_imag;
        _zz_260 = img_reg_array_33_37_real;
        _zz_261 = img_reg_array_33_37_imag;
        _zz_262 = img_reg_array_34_37_real;
        _zz_263 = img_reg_array_34_37_imag;
        _zz_264 = img_reg_array_35_37_real;
        _zz_265 = img_reg_array_35_37_imag;
        _zz_266 = img_reg_array_36_37_real;
        _zz_267 = img_reg_array_36_37_imag;
        _zz_268 = img_reg_array_37_37_real;
        _zz_269 = img_reg_array_37_37_imag;
        _zz_270 = img_reg_array_38_37_real;
        _zz_271 = img_reg_array_38_37_imag;
        _zz_272 = img_reg_array_39_37_real;
        _zz_273 = img_reg_array_39_37_imag;
        _zz_274 = img_reg_array_40_37_real;
        _zz_275 = img_reg_array_40_37_imag;
        _zz_276 = img_reg_array_41_37_real;
        _zz_277 = img_reg_array_41_37_imag;
        _zz_278 = img_reg_array_42_37_real;
        _zz_279 = img_reg_array_42_37_imag;
        _zz_280 = img_reg_array_43_37_real;
        _zz_281 = img_reg_array_43_37_imag;
        _zz_282 = img_reg_array_44_37_real;
        _zz_283 = img_reg_array_44_37_imag;
        _zz_284 = img_reg_array_45_37_real;
        _zz_285 = img_reg_array_45_37_imag;
        _zz_286 = img_reg_array_46_37_real;
        _zz_287 = img_reg_array_46_37_imag;
        _zz_288 = img_reg_array_47_37_real;
        _zz_289 = img_reg_array_47_37_imag;
        _zz_290 = img_reg_array_48_37_real;
        _zz_291 = img_reg_array_48_37_imag;
        _zz_292 = img_reg_array_49_37_real;
        _zz_293 = img_reg_array_49_37_imag;
        _zz_294 = img_reg_array_50_37_real;
        _zz_295 = img_reg_array_50_37_imag;
        _zz_296 = img_reg_array_51_37_real;
        _zz_297 = img_reg_array_51_37_imag;
        _zz_298 = img_reg_array_52_37_real;
        _zz_299 = img_reg_array_52_37_imag;
        _zz_300 = img_reg_array_53_37_real;
        _zz_301 = img_reg_array_53_37_imag;
        _zz_302 = img_reg_array_54_37_real;
        _zz_303 = img_reg_array_54_37_imag;
        _zz_304 = img_reg_array_55_37_real;
        _zz_305 = img_reg_array_55_37_imag;
        _zz_306 = img_reg_array_56_37_real;
        _zz_307 = img_reg_array_56_37_imag;
        _zz_308 = img_reg_array_57_37_real;
        _zz_309 = img_reg_array_57_37_imag;
        _zz_310 = img_reg_array_58_37_real;
        _zz_311 = img_reg_array_58_37_imag;
        _zz_312 = img_reg_array_59_37_real;
        _zz_313 = img_reg_array_59_37_imag;
        _zz_314 = img_reg_array_60_37_real;
        _zz_315 = img_reg_array_60_37_imag;
        _zz_316 = img_reg_array_61_37_real;
        _zz_317 = img_reg_array_61_37_imag;
        _zz_318 = img_reg_array_62_37_real;
        _zz_319 = img_reg_array_62_37_imag;
        _zz_320 = img_reg_array_63_37_real;
        _zz_321 = img_reg_array_63_37_imag;
      end
      6'b100110 : begin
        _zz_194 = img_reg_array_0_38_real;
        _zz_195 = img_reg_array_0_38_imag;
        _zz_196 = img_reg_array_1_38_real;
        _zz_197 = img_reg_array_1_38_imag;
        _zz_198 = img_reg_array_2_38_real;
        _zz_199 = img_reg_array_2_38_imag;
        _zz_200 = img_reg_array_3_38_real;
        _zz_201 = img_reg_array_3_38_imag;
        _zz_202 = img_reg_array_4_38_real;
        _zz_203 = img_reg_array_4_38_imag;
        _zz_204 = img_reg_array_5_38_real;
        _zz_205 = img_reg_array_5_38_imag;
        _zz_206 = img_reg_array_6_38_real;
        _zz_207 = img_reg_array_6_38_imag;
        _zz_208 = img_reg_array_7_38_real;
        _zz_209 = img_reg_array_7_38_imag;
        _zz_210 = img_reg_array_8_38_real;
        _zz_211 = img_reg_array_8_38_imag;
        _zz_212 = img_reg_array_9_38_real;
        _zz_213 = img_reg_array_9_38_imag;
        _zz_214 = img_reg_array_10_38_real;
        _zz_215 = img_reg_array_10_38_imag;
        _zz_216 = img_reg_array_11_38_real;
        _zz_217 = img_reg_array_11_38_imag;
        _zz_218 = img_reg_array_12_38_real;
        _zz_219 = img_reg_array_12_38_imag;
        _zz_220 = img_reg_array_13_38_real;
        _zz_221 = img_reg_array_13_38_imag;
        _zz_222 = img_reg_array_14_38_real;
        _zz_223 = img_reg_array_14_38_imag;
        _zz_224 = img_reg_array_15_38_real;
        _zz_225 = img_reg_array_15_38_imag;
        _zz_226 = img_reg_array_16_38_real;
        _zz_227 = img_reg_array_16_38_imag;
        _zz_228 = img_reg_array_17_38_real;
        _zz_229 = img_reg_array_17_38_imag;
        _zz_230 = img_reg_array_18_38_real;
        _zz_231 = img_reg_array_18_38_imag;
        _zz_232 = img_reg_array_19_38_real;
        _zz_233 = img_reg_array_19_38_imag;
        _zz_234 = img_reg_array_20_38_real;
        _zz_235 = img_reg_array_20_38_imag;
        _zz_236 = img_reg_array_21_38_real;
        _zz_237 = img_reg_array_21_38_imag;
        _zz_238 = img_reg_array_22_38_real;
        _zz_239 = img_reg_array_22_38_imag;
        _zz_240 = img_reg_array_23_38_real;
        _zz_241 = img_reg_array_23_38_imag;
        _zz_242 = img_reg_array_24_38_real;
        _zz_243 = img_reg_array_24_38_imag;
        _zz_244 = img_reg_array_25_38_real;
        _zz_245 = img_reg_array_25_38_imag;
        _zz_246 = img_reg_array_26_38_real;
        _zz_247 = img_reg_array_26_38_imag;
        _zz_248 = img_reg_array_27_38_real;
        _zz_249 = img_reg_array_27_38_imag;
        _zz_250 = img_reg_array_28_38_real;
        _zz_251 = img_reg_array_28_38_imag;
        _zz_252 = img_reg_array_29_38_real;
        _zz_253 = img_reg_array_29_38_imag;
        _zz_254 = img_reg_array_30_38_real;
        _zz_255 = img_reg_array_30_38_imag;
        _zz_256 = img_reg_array_31_38_real;
        _zz_257 = img_reg_array_31_38_imag;
        _zz_258 = img_reg_array_32_38_real;
        _zz_259 = img_reg_array_32_38_imag;
        _zz_260 = img_reg_array_33_38_real;
        _zz_261 = img_reg_array_33_38_imag;
        _zz_262 = img_reg_array_34_38_real;
        _zz_263 = img_reg_array_34_38_imag;
        _zz_264 = img_reg_array_35_38_real;
        _zz_265 = img_reg_array_35_38_imag;
        _zz_266 = img_reg_array_36_38_real;
        _zz_267 = img_reg_array_36_38_imag;
        _zz_268 = img_reg_array_37_38_real;
        _zz_269 = img_reg_array_37_38_imag;
        _zz_270 = img_reg_array_38_38_real;
        _zz_271 = img_reg_array_38_38_imag;
        _zz_272 = img_reg_array_39_38_real;
        _zz_273 = img_reg_array_39_38_imag;
        _zz_274 = img_reg_array_40_38_real;
        _zz_275 = img_reg_array_40_38_imag;
        _zz_276 = img_reg_array_41_38_real;
        _zz_277 = img_reg_array_41_38_imag;
        _zz_278 = img_reg_array_42_38_real;
        _zz_279 = img_reg_array_42_38_imag;
        _zz_280 = img_reg_array_43_38_real;
        _zz_281 = img_reg_array_43_38_imag;
        _zz_282 = img_reg_array_44_38_real;
        _zz_283 = img_reg_array_44_38_imag;
        _zz_284 = img_reg_array_45_38_real;
        _zz_285 = img_reg_array_45_38_imag;
        _zz_286 = img_reg_array_46_38_real;
        _zz_287 = img_reg_array_46_38_imag;
        _zz_288 = img_reg_array_47_38_real;
        _zz_289 = img_reg_array_47_38_imag;
        _zz_290 = img_reg_array_48_38_real;
        _zz_291 = img_reg_array_48_38_imag;
        _zz_292 = img_reg_array_49_38_real;
        _zz_293 = img_reg_array_49_38_imag;
        _zz_294 = img_reg_array_50_38_real;
        _zz_295 = img_reg_array_50_38_imag;
        _zz_296 = img_reg_array_51_38_real;
        _zz_297 = img_reg_array_51_38_imag;
        _zz_298 = img_reg_array_52_38_real;
        _zz_299 = img_reg_array_52_38_imag;
        _zz_300 = img_reg_array_53_38_real;
        _zz_301 = img_reg_array_53_38_imag;
        _zz_302 = img_reg_array_54_38_real;
        _zz_303 = img_reg_array_54_38_imag;
        _zz_304 = img_reg_array_55_38_real;
        _zz_305 = img_reg_array_55_38_imag;
        _zz_306 = img_reg_array_56_38_real;
        _zz_307 = img_reg_array_56_38_imag;
        _zz_308 = img_reg_array_57_38_real;
        _zz_309 = img_reg_array_57_38_imag;
        _zz_310 = img_reg_array_58_38_real;
        _zz_311 = img_reg_array_58_38_imag;
        _zz_312 = img_reg_array_59_38_real;
        _zz_313 = img_reg_array_59_38_imag;
        _zz_314 = img_reg_array_60_38_real;
        _zz_315 = img_reg_array_60_38_imag;
        _zz_316 = img_reg_array_61_38_real;
        _zz_317 = img_reg_array_61_38_imag;
        _zz_318 = img_reg_array_62_38_real;
        _zz_319 = img_reg_array_62_38_imag;
        _zz_320 = img_reg_array_63_38_real;
        _zz_321 = img_reg_array_63_38_imag;
      end
      6'b100111 : begin
        _zz_194 = img_reg_array_0_39_real;
        _zz_195 = img_reg_array_0_39_imag;
        _zz_196 = img_reg_array_1_39_real;
        _zz_197 = img_reg_array_1_39_imag;
        _zz_198 = img_reg_array_2_39_real;
        _zz_199 = img_reg_array_2_39_imag;
        _zz_200 = img_reg_array_3_39_real;
        _zz_201 = img_reg_array_3_39_imag;
        _zz_202 = img_reg_array_4_39_real;
        _zz_203 = img_reg_array_4_39_imag;
        _zz_204 = img_reg_array_5_39_real;
        _zz_205 = img_reg_array_5_39_imag;
        _zz_206 = img_reg_array_6_39_real;
        _zz_207 = img_reg_array_6_39_imag;
        _zz_208 = img_reg_array_7_39_real;
        _zz_209 = img_reg_array_7_39_imag;
        _zz_210 = img_reg_array_8_39_real;
        _zz_211 = img_reg_array_8_39_imag;
        _zz_212 = img_reg_array_9_39_real;
        _zz_213 = img_reg_array_9_39_imag;
        _zz_214 = img_reg_array_10_39_real;
        _zz_215 = img_reg_array_10_39_imag;
        _zz_216 = img_reg_array_11_39_real;
        _zz_217 = img_reg_array_11_39_imag;
        _zz_218 = img_reg_array_12_39_real;
        _zz_219 = img_reg_array_12_39_imag;
        _zz_220 = img_reg_array_13_39_real;
        _zz_221 = img_reg_array_13_39_imag;
        _zz_222 = img_reg_array_14_39_real;
        _zz_223 = img_reg_array_14_39_imag;
        _zz_224 = img_reg_array_15_39_real;
        _zz_225 = img_reg_array_15_39_imag;
        _zz_226 = img_reg_array_16_39_real;
        _zz_227 = img_reg_array_16_39_imag;
        _zz_228 = img_reg_array_17_39_real;
        _zz_229 = img_reg_array_17_39_imag;
        _zz_230 = img_reg_array_18_39_real;
        _zz_231 = img_reg_array_18_39_imag;
        _zz_232 = img_reg_array_19_39_real;
        _zz_233 = img_reg_array_19_39_imag;
        _zz_234 = img_reg_array_20_39_real;
        _zz_235 = img_reg_array_20_39_imag;
        _zz_236 = img_reg_array_21_39_real;
        _zz_237 = img_reg_array_21_39_imag;
        _zz_238 = img_reg_array_22_39_real;
        _zz_239 = img_reg_array_22_39_imag;
        _zz_240 = img_reg_array_23_39_real;
        _zz_241 = img_reg_array_23_39_imag;
        _zz_242 = img_reg_array_24_39_real;
        _zz_243 = img_reg_array_24_39_imag;
        _zz_244 = img_reg_array_25_39_real;
        _zz_245 = img_reg_array_25_39_imag;
        _zz_246 = img_reg_array_26_39_real;
        _zz_247 = img_reg_array_26_39_imag;
        _zz_248 = img_reg_array_27_39_real;
        _zz_249 = img_reg_array_27_39_imag;
        _zz_250 = img_reg_array_28_39_real;
        _zz_251 = img_reg_array_28_39_imag;
        _zz_252 = img_reg_array_29_39_real;
        _zz_253 = img_reg_array_29_39_imag;
        _zz_254 = img_reg_array_30_39_real;
        _zz_255 = img_reg_array_30_39_imag;
        _zz_256 = img_reg_array_31_39_real;
        _zz_257 = img_reg_array_31_39_imag;
        _zz_258 = img_reg_array_32_39_real;
        _zz_259 = img_reg_array_32_39_imag;
        _zz_260 = img_reg_array_33_39_real;
        _zz_261 = img_reg_array_33_39_imag;
        _zz_262 = img_reg_array_34_39_real;
        _zz_263 = img_reg_array_34_39_imag;
        _zz_264 = img_reg_array_35_39_real;
        _zz_265 = img_reg_array_35_39_imag;
        _zz_266 = img_reg_array_36_39_real;
        _zz_267 = img_reg_array_36_39_imag;
        _zz_268 = img_reg_array_37_39_real;
        _zz_269 = img_reg_array_37_39_imag;
        _zz_270 = img_reg_array_38_39_real;
        _zz_271 = img_reg_array_38_39_imag;
        _zz_272 = img_reg_array_39_39_real;
        _zz_273 = img_reg_array_39_39_imag;
        _zz_274 = img_reg_array_40_39_real;
        _zz_275 = img_reg_array_40_39_imag;
        _zz_276 = img_reg_array_41_39_real;
        _zz_277 = img_reg_array_41_39_imag;
        _zz_278 = img_reg_array_42_39_real;
        _zz_279 = img_reg_array_42_39_imag;
        _zz_280 = img_reg_array_43_39_real;
        _zz_281 = img_reg_array_43_39_imag;
        _zz_282 = img_reg_array_44_39_real;
        _zz_283 = img_reg_array_44_39_imag;
        _zz_284 = img_reg_array_45_39_real;
        _zz_285 = img_reg_array_45_39_imag;
        _zz_286 = img_reg_array_46_39_real;
        _zz_287 = img_reg_array_46_39_imag;
        _zz_288 = img_reg_array_47_39_real;
        _zz_289 = img_reg_array_47_39_imag;
        _zz_290 = img_reg_array_48_39_real;
        _zz_291 = img_reg_array_48_39_imag;
        _zz_292 = img_reg_array_49_39_real;
        _zz_293 = img_reg_array_49_39_imag;
        _zz_294 = img_reg_array_50_39_real;
        _zz_295 = img_reg_array_50_39_imag;
        _zz_296 = img_reg_array_51_39_real;
        _zz_297 = img_reg_array_51_39_imag;
        _zz_298 = img_reg_array_52_39_real;
        _zz_299 = img_reg_array_52_39_imag;
        _zz_300 = img_reg_array_53_39_real;
        _zz_301 = img_reg_array_53_39_imag;
        _zz_302 = img_reg_array_54_39_real;
        _zz_303 = img_reg_array_54_39_imag;
        _zz_304 = img_reg_array_55_39_real;
        _zz_305 = img_reg_array_55_39_imag;
        _zz_306 = img_reg_array_56_39_real;
        _zz_307 = img_reg_array_56_39_imag;
        _zz_308 = img_reg_array_57_39_real;
        _zz_309 = img_reg_array_57_39_imag;
        _zz_310 = img_reg_array_58_39_real;
        _zz_311 = img_reg_array_58_39_imag;
        _zz_312 = img_reg_array_59_39_real;
        _zz_313 = img_reg_array_59_39_imag;
        _zz_314 = img_reg_array_60_39_real;
        _zz_315 = img_reg_array_60_39_imag;
        _zz_316 = img_reg_array_61_39_real;
        _zz_317 = img_reg_array_61_39_imag;
        _zz_318 = img_reg_array_62_39_real;
        _zz_319 = img_reg_array_62_39_imag;
        _zz_320 = img_reg_array_63_39_real;
        _zz_321 = img_reg_array_63_39_imag;
      end
      6'b101000 : begin
        _zz_194 = img_reg_array_0_40_real;
        _zz_195 = img_reg_array_0_40_imag;
        _zz_196 = img_reg_array_1_40_real;
        _zz_197 = img_reg_array_1_40_imag;
        _zz_198 = img_reg_array_2_40_real;
        _zz_199 = img_reg_array_2_40_imag;
        _zz_200 = img_reg_array_3_40_real;
        _zz_201 = img_reg_array_3_40_imag;
        _zz_202 = img_reg_array_4_40_real;
        _zz_203 = img_reg_array_4_40_imag;
        _zz_204 = img_reg_array_5_40_real;
        _zz_205 = img_reg_array_5_40_imag;
        _zz_206 = img_reg_array_6_40_real;
        _zz_207 = img_reg_array_6_40_imag;
        _zz_208 = img_reg_array_7_40_real;
        _zz_209 = img_reg_array_7_40_imag;
        _zz_210 = img_reg_array_8_40_real;
        _zz_211 = img_reg_array_8_40_imag;
        _zz_212 = img_reg_array_9_40_real;
        _zz_213 = img_reg_array_9_40_imag;
        _zz_214 = img_reg_array_10_40_real;
        _zz_215 = img_reg_array_10_40_imag;
        _zz_216 = img_reg_array_11_40_real;
        _zz_217 = img_reg_array_11_40_imag;
        _zz_218 = img_reg_array_12_40_real;
        _zz_219 = img_reg_array_12_40_imag;
        _zz_220 = img_reg_array_13_40_real;
        _zz_221 = img_reg_array_13_40_imag;
        _zz_222 = img_reg_array_14_40_real;
        _zz_223 = img_reg_array_14_40_imag;
        _zz_224 = img_reg_array_15_40_real;
        _zz_225 = img_reg_array_15_40_imag;
        _zz_226 = img_reg_array_16_40_real;
        _zz_227 = img_reg_array_16_40_imag;
        _zz_228 = img_reg_array_17_40_real;
        _zz_229 = img_reg_array_17_40_imag;
        _zz_230 = img_reg_array_18_40_real;
        _zz_231 = img_reg_array_18_40_imag;
        _zz_232 = img_reg_array_19_40_real;
        _zz_233 = img_reg_array_19_40_imag;
        _zz_234 = img_reg_array_20_40_real;
        _zz_235 = img_reg_array_20_40_imag;
        _zz_236 = img_reg_array_21_40_real;
        _zz_237 = img_reg_array_21_40_imag;
        _zz_238 = img_reg_array_22_40_real;
        _zz_239 = img_reg_array_22_40_imag;
        _zz_240 = img_reg_array_23_40_real;
        _zz_241 = img_reg_array_23_40_imag;
        _zz_242 = img_reg_array_24_40_real;
        _zz_243 = img_reg_array_24_40_imag;
        _zz_244 = img_reg_array_25_40_real;
        _zz_245 = img_reg_array_25_40_imag;
        _zz_246 = img_reg_array_26_40_real;
        _zz_247 = img_reg_array_26_40_imag;
        _zz_248 = img_reg_array_27_40_real;
        _zz_249 = img_reg_array_27_40_imag;
        _zz_250 = img_reg_array_28_40_real;
        _zz_251 = img_reg_array_28_40_imag;
        _zz_252 = img_reg_array_29_40_real;
        _zz_253 = img_reg_array_29_40_imag;
        _zz_254 = img_reg_array_30_40_real;
        _zz_255 = img_reg_array_30_40_imag;
        _zz_256 = img_reg_array_31_40_real;
        _zz_257 = img_reg_array_31_40_imag;
        _zz_258 = img_reg_array_32_40_real;
        _zz_259 = img_reg_array_32_40_imag;
        _zz_260 = img_reg_array_33_40_real;
        _zz_261 = img_reg_array_33_40_imag;
        _zz_262 = img_reg_array_34_40_real;
        _zz_263 = img_reg_array_34_40_imag;
        _zz_264 = img_reg_array_35_40_real;
        _zz_265 = img_reg_array_35_40_imag;
        _zz_266 = img_reg_array_36_40_real;
        _zz_267 = img_reg_array_36_40_imag;
        _zz_268 = img_reg_array_37_40_real;
        _zz_269 = img_reg_array_37_40_imag;
        _zz_270 = img_reg_array_38_40_real;
        _zz_271 = img_reg_array_38_40_imag;
        _zz_272 = img_reg_array_39_40_real;
        _zz_273 = img_reg_array_39_40_imag;
        _zz_274 = img_reg_array_40_40_real;
        _zz_275 = img_reg_array_40_40_imag;
        _zz_276 = img_reg_array_41_40_real;
        _zz_277 = img_reg_array_41_40_imag;
        _zz_278 = img_reg_array_42_40_real;
        _zz_279 = img_reg_array_42_40_imag;
        _zz_280 = img_reg_array_43_40_real;
        _zz_281 = img_reg_array_43_40_imag;
        _zz_282 = img_reg_array_44_40_real;
        _zz_283 = img_reg_array_44_40_imag;
        _zz_284 = img_reg_array_45_40_real;
        _zz_285 = img_reg_array_45_40_imag;
        _zz_286 = img_reg_array_46_40_real;
        _zz_287 = img_reg_array_46_40_imag;
        _zz_288 = img_reg_array_47_40_real;
        _zz_289 = img_reg_array_47_40_imag;
        _zz_290 = img_reg_array_48_40_real;
        _zz_291 = img_reg_array_48_40_imag;
        _zz_292 = img_reg_array_49_40_real;
        _zz_293 = img_reg_array_49_40_imag;
        _zz_294 = img_reg_array_50_40_real;
        _zz_295 = img_reg_array_50_40_imag;
        _zz_296 = img_reg_array_51_40_real;
        _zz_297 = img_reg_array_51_40_imag;
        _zz_298 = img_reg_array_52_40_real;
        _zz_299 = img_reg_array_52_40_imag;
        _zz_300 = img_reg_array_53_40_real;
        _zz_301 = img_reg_array_53_40_imag;
        _zz_302 = img_reg_array_54_40_real;
        _zz_303 = img_reg_array_54_40_imag;
        _zz_304 = img_reg_array_55_40_real;
        _zz_305 = img_reg_array_55_40_imag;
        _zz_306 = img_reg_array_56_40_real;
        _zz_307 = img_reg_array_56_40_imag;
        _zz_308 = img_reg_array_57_40_real;
        _zz_309 = img_reg_array_57_40_imag;
        _zz_310 = img_reg_array_58_40_real;
        _zz_311 = img_reg_array_58_40_imag;
        _zz_312 = img_reg_array_59_40_real;
        _zz_313 = img_reg_array_59_40_imag;
        _zz_314 = img_reg_array_60_40_real;
        _zz_315 = img_reg_array_60_40_imag;
        _zz_316 = img_reg_array_61_40_real;
        _zz_317 = img_reg_array_61_40_imag;
        _zz_318 = img_reg_array_62_40_real;
        _zz_319 = img_reg_array_62_40_imag;
        _zz_320 = img_reg_array_63_40_real;
        _zz_321 = img_reg_array_63_40_imag;
      end
      6'b101001 : begin
        _zz_194 = img_reg_array_0_41_real;
        _zz_195 = img_reg_array_0_41_imag;
        _zz_196 = img_reg_array_1_41_real;
        _zz_197 = img_reg_array_1_41_imag;
        _zz_198 = img_reg_array_2_41_real;
        _zz_199 = img_reg_array_2_41_imag;
        _zz_200 = img_reg_array_3_41_real;
        _zz_201 = img_reg_array_3_41_imag;
        _zz_202 = img_reg_array_4_41_real;
        _zz_203 = img_reg_array_4_41_imag;
        _zz_204 = img_reg_array_5_41_real;
        _zz_205 = img_reg_array_5_41_imag;
        _zz_206 = img_reg_array_6_41_real;
        _zz_207 = img_reg_array_6_41_imag;
        _zz_208 = img_reg_array_7_41_real;
        _zz_209 = img_reg_array_7_41_imag;
        _zz_210 = img_reg_array_8_41_real;
        _zz_211 = img_reg_array_8_41_imag;
        _zz_212 = img_reg_array_9_41_real;
        _zz_213 = img_reg_array_9_41_imag;
        _zz_214 = img_reg_array_10_41_real;
        _zz_215 = img_reg_array_10_41_imag;
        _zz_216 = img_reg_array_11_41_real;
        _zz_217 = img_reg_array_11_41_imag;
        _zz_218 = img_reg_array_12_41_real;
        _zz_219 = img_reg_array_12_41_imag;
        _zz_220 = img_reg_array_13_41_real;
        _zz_221 = img_reg_array_13_41_imag;
        _zz_222 = img_reg_array_14_41_real;
        _zz_223 = img_reg_array_14_41_imag;
        _zz_224 = img_reg_array_15_41_real;
        _zz_225 = img_reg_array_15_41_imag;
        _zz_226 = img_reg_array_16_41_real;
        _zz_227 = img_reg_array_16_41_imag;
        _zz_228 = img_reg_array_17_41_real;
        _zz_229 = img_reg_array_17_41_imag;
        _zz_230 = img_reg_array_18_41_real;
        _zz_231 = img_reg_array_18_41_imag;
        _zz_232 = img_reg_array_19_41_real;
        _zz_233 = img_reg_array_19_41_imag;
        _zz_234 = img_reg_array_20_41_real;
        _zz_235 = img_reg_array_20_41_imag;
        _zz_236 = img_reg_array_21_41_real;
        _zz_237 = img_reg_array_21_41_imag;
        _zz_238 = img_reg_array_22_41_real;
        _zz_239 = img_reg_array_22_41_imag;
        _zz_240 = img_reg_array_23_41_real;
        _zz_241 = img_reg_array_23_41_imag;
        _zz_242 = img_reg_array_24_41_real;
        _zz_243 = img_reg_array_24_41_imag;
        _zz_244 = img_reg_array_25_41_real;
        _zz_245 = img_reg_array_25_41_imag;
        _zz_246 = img_reg_array_26_41_real;
        _zz_247 = img_reg_array_26_41_imag;
        _zz_248 = img_reg_array_27_41_real;
        _zz_249 = img_reg_array_27_41_imag;
        _zz_250 = img_reg_array_28_41_real;
        _zz_251 = img_reg_array_28_41_imag;
        _zz_252 = img_reg_array_29_41_real;
        _zz_253 = img_reg_array_29_41_imag;
        _zz_254 = img_reg_array_30_41_real;
        _zz_255 = img_reg_array_30_41_imag;
        _zz_256 = img_reg_array_31_41_real;
        _zz_257 = img_reg_array_31_41_imag;
        _zz_258 = img_reg_array_32_41_real;
        _zz_259 = img_reg_array_32_41_imag;
        _zz_260 = img_reg_array_33_41_real;
        _zz_261 = img_reg_array_33_41_imag;
        _zz_262 = img_reg_array_34_41_real;
        _zz_263 = img_reg_array_34_41_imag;
        _zz_264 = img_reg_array_35_41_real;
        _zz_265 = img_reg_array_35_41_imag;
        _zz_266 = img_reg_array_36_41_real;
        _zz_267 = img_reg_array_36_41_imag;
        _zz_268 = img_reg_array_37_41_real;
        _zz_269 = img_reg_array_37_41_imag;
        _zz_270 = img_reg_array_38_41_real;
        _zz_271 = img_reg_array_38_41_imag;
        _zz_272 = img_reg_array_39_41_real;
        _zz_273 = img_reg_array_39_41_imag;
        _zz_274 = img_reg_array_40_41_real;
        _zz_275 = img_reg_array_40_41_imag;
        _zz_276 = img_reg_array_41_41_real;
        _zz_277 = img_reg_array_41_41_imag;
        _zz_278 = img_reg_array_42_41_real;
        _zz_279 = img_reg_array_42_41_imag;
        _zz_280 = img_reg_array_43_41_real;
        _zz_281 = img_reg_array_43_41_imag;
        _zz_282 = img_reg_array_44_41_real;
        _zz_283 = img_reg_array_44_41_imag;
        _zz_284 = img_reg_array_45_41_real;
        _zz_285 = img_reg_array_45_41_imag;
        _zz_286 = img_reg_array_46_41_real;
        _zz_287 = img_reg_array_46_41_imag;
        _zz_288 = img_reg_array_47_41_real;
        _zz_289 = img_reg_array_47_41_imag;
        _zz_290 = img_reg_array_48_41_real;
        _zz_291 = img_reg_array_48_41_imag;
        _zz_292 = img_reg_array_49_41_real;
        _zz_293 = img_reg_array_49_41_imag;
        _zz_294 = img_reg_array_50_41_real;
        _zz_295 = img_reg_array_50_41_imag;
        _zz_296 = img_reg_array_51_41_real;
        _zz_297 = img_reg_array_51_41_imag;
        _zz_298 = img_reg_array_52_41_real;
        _zz_299 = img_reg_array_52_41_imag;
        _zz_300 = img_reg_array_53_41_real;
        _zz_301 = img_reg_array_53_41_imag;
        _zz_302 = img_reg_array_54_41_real;
        _zz_303 = img_reg_array_54_41_imag;
        _zz_304 = img_reg_array_55_41_real;
        _zz_305 = img_reg_array_55_41_imag;
        _zz_306 = img_reg_array_56_41_real;
        _zz_307 = img_reg_array_56_41_imag;
        _zz_308 = img_reg_array_57_41_real;
        _zz_309 = img_reg_array_57_41_imag;
        _zz_310 = img_reg_array_58_41_real;
        _zz_311 = img_reg_array_58_41_imag;
        _zz_312 = img_reg_array_59_41_real;
        _zz_313 = img_reg_array_59_41_imag;
        _zz_314 = img_reg_array_60_41_real;
        _zz_315 = img_reg_array_60_41_imag;
        _zz_316 = img_reg_array_61_41_real;
        _zz_317 = img_reg_array_61_41_imag;
        _zz_318 = img_reg_array_62_41_real;
        _zz_319 = img_reg_array_62_41_imag;
        _zz_320 = img_reg_array_63_41_real;
        _zz_321 = img_reg_array_63_41_imag;
      end
      6'b101010 : begin
        _zz_194 = img_reg_array_0_42_real;
        _zz_195 = img_reg_array_0_42_imag;
        _zz_196 = img_reg_array_1_42_real;
        _zz_197 = img_reg_array_1_42_imag;
        _zz_198 = img_reg_array_2_42_real;
        _zz_199 = img_reg_array_2_42_imag;
        _zz_200 = img_reg_array_3_42_real;
        _zz_201 = img_reg_array_3_42_imag;
        _zz_202 = img_reg_array_4_42_real;
        _zz_203 = img_reg_array_4_42_imag;
        _zz_204 = img_reg_array_5_42_real;
        _zz_205 = img_reg_array_5_42_imag;
        _zz_206 = img_reg_array_6_42_real;
        _zz_207 = img_reg_array_6_42_imag;
        _zz_208 = img_reg_array_7_42_real;
        _zz_209 = img_reg_array_7_42_imag;
        _zz_210 = img_reg_array_8_42_real;
        _zz_211 = img_reg_array_8_42_imag;
        _zz_212 = img_reg_array_9_42_real;
        _zz_213 = img_reg_array_9_42_imag;
        _zz_214 = img_reg_array_10_42_real;
        _zz_215 = img_reg_array_10_42_imag;
        _zz_216 = img_reg_array_11_42_real;
        _zz_217 = img_reg_array_11_42_imag;
        _zz_218 = img_reg_array_12_42_real;
        _zz_219 = img_reg_array_12_42_imag;
        _zz_220 = img_reg_array_13_42_real;
        _zz_221 = img_reg_array_13_42_imag;
        _zz_222 = img_reg_array_14_42_real;
        _zz_223 = img_reg_array_14_42_imag;
        _zz_224 = img_reg_array_15_42_real;
        _zz_225 = img_reg_array_15_42_imag;
        _zz_226 = img_reg_array_16_42_real;
        _zz_227 = img_reg_array_16_42_imag;
        _zz_228 = img_reg_array_17_42_real;
        _zz_229 = img_reg_array_17_42_imag;
        _zz_230 = img_reg_array_18_42_real;
        _zz_231 = img_reg_array_18_42_imag;
        _zz_232 = img_reg_array_19_42_real;
        _zz_233 = img_reg_array_19_42_imag;
        _zz_234 = img_reg_array_20_42_real;
        _zz_235 = img_reg_array_20_42_imag;
        _zz_236 = img_reg_array_21_42_real;
        _zz_237 = img_reg_array_21_42_imag;
        _zz_238 = img_reg_array_22_42_real;
        _zz_239 = img_reg_array_22_42_imag;
        _zz_240 = img_reg_array_23_42_real;
        _zz_241 = img_reg_array_23_42_imag;
        _zz_242 = img_reg_array_24_42_real;
        _zz_243 = img_reg_array_24_42_imag;
        _zz_244 = img_reg_array_25_42_real;
        _zz_245 = img_reg_array_25_42_imag;
        _zz_246 = img_reg_array_26_42_real;
        _zz_247 = img_reg_array_26_42_imag;
        _zz_248 = img_reg_array_27_42_real;
        _zz_249 = img_reg_array_27_42_imag;
        _zz_250 = img_reg_array_28_42_real;
        _zz_251 = img_reg_array_28_42_imag;
        _zz_252 = img_reg_array_29_42_real;
        _zz_253 = img_reg_array_29_42_imag;
        _zz_254 = img_reg_array_30_42_real;
        _zz_255 = img_reg_array_30_42_imag;
        _zz_256 = img_reg_array_31_42_real;
        _zz_257 = img_reg_array_31_42_imag;
        _zz_258 = img_reg_array_32_42_real;
        _zz_259 = img_reg_array_32_42_imag;
        _zz_260 = img_reg_array_33_42_real;
        _zz_261 = img_reg_array_33_42_imag;
        _zz_262 = img_reg_array_34_42_real;
        _zz_263 = img_reg_array_34_42_imag;
        _zz_264 = img_reg_array_35_42_real;
        _zz_265 = img_reg_array_35_42_imag;
        _zz_266 = img_reg_array_36_42_real;
        _zz_267 = img_reg_array_36_42_imag;
        _zz_268 = img_reg_array_37_42_real;
        _zz_269 = img_reg_array_37_42_imag;
        _zz_270 = img_reg_array_38_42_real;
        _zz_271 = img_reg_array_38_42_imag;
        _zz_272 = img_reg_array_39_42_real;
        _zz_273 = img_reg_array_39_42_imag;
        _zz_274 = img_reg_array_40_42_real;
        _zz_275 = img_reg_array_40_42_imag;
        _zz_276 = img_reg_array_41_42_real;
        _zz_277 = img_reg_array_41_42_imag;
        _zz_278 = img_reg_array_42_42_real;
        _zz_279 = img_reg_array_42_42_imag;
        _zz_280 = img_reg_array_43_42_real;
        _zz_281 = img_reg_array_43_42_imag;
        _zz_282 = img_reg_array_44_42_real;
        _zz_283 = img_reg_array_44_42_imag;
        _zz_284 = img_reg_array_45_42_real;
        _zz_285 = img_reg_array_45_42_imag;
        _zz_286 = img_reg_array_46_42_real;
        _zz_287 = img_reg_array_46_42_imag;
        _zz_288 = img_reg_array_47_42_real;
        _zz_289 = img_reg_array_47_42_imag;
        _zz_290 = img_reg_array_48_42_real;
        _zz_291 = img_reg_array_48_42_imag;
        _zz_292 = img_reg_array_49_42_real;
        _zz_293 = img_reg_array_49_42_imag;
        _zz_294 = img_reg_array_50_42_real;
        _zz_295 = img_reg_array_50_42_imag;
        _zz_296 = img_reg_array_51_42_real;
        _zz_297 = img_reg_array_51_42_imag;
        _zz_298 = img_reg_array_52_42_real;
        _zz_299 = img_reg_array_52_42_imag;
        _zz_300 = img_reg_array_53_42_real;
        _zz_301 = img_reg_array_53_42_imag;
        _zz_302 = img_reg_array_54_42_real;
        _zz_303 = img_reg_array_54_42_imag;
        _zz_304 = img_reg_array_55_42_real;
        _zz_305 = img_reg_array_55_42_imag;
        _zz_306 = img_reg_array_56_42_real;
        _zz_307 = img_reg_array_56_42_imag;
        _zz_308 = img_reg_array_57_42_real;
        _zz_309 = img_reg_array_57_42_imag;
        _zz_310 = img_reg_array_58_42_real;
        _zz_311 = img_reg_array_58_42_imag;
        _zz_312 = img_reg_array_59_42_real;
        _zz_313 = img_reg_array_59_42_imag;
        _zz_314 = img_reg_array_60_42_real;
        _zz_315 = img_reg_array_60_42_imag;
        _zz_316 = img_reg_array_61_42_real;
        _zz_317 = img_reg_array_61_42_imag;
        _zz_318 = img_reg_array_62_42_real;
        _zz_319 = img_reg_array_62_42_imag;
        _zz_320 = img_reg_array_63_42_real;
        _zz_321 = img_reg_array_63_42_imag;
      end
      6'b101011 : begin
        _zz_194 = img_reg_array_0_43_real;
        _zz_195 = img_reg_array_0_43_imag;
        _zz_196 = img_reg_array_1_43_real;
        _zz_197 = img_reg_array_1_43_imag;
        _zz_198 = img_reg_array_2_43_real;
        _zz_199 = img_reg_array_2_43_imag;
        _zz_200 = img_reg_array_3_43_real;
        _zz_201 = img_reg_array_3_43_imag;
        _zz_202 = img_reg_array_4_43_real;
        _zz_203 = img_reg_array_4_43_imag;
        _zz_204 = img_reg_array_5_43_real;
        _zz_205 = img_reg_array_5_43_imag;
        _zz_206 = img_reg_array_6_43_real;
        _zz_207 = img_reg_array_6_43_imag;
        _zz_208 = img_reg_array_7_43_real;
        _zz_209 = img_reg_array_7_43_imag;
        _zz_210 = img_reg_array_8_43_real;
        _zz_211 = img_reg_array_8_43_imag;
        _zz_212 = img_reg_array_9_43_real;
        _zz_213 = img_reg_array_9_43_imag;
        _zz_214 = img_reg_array_10_43_real;
        _zz_215 = img_reg_array_10_43_imag;
        _zz_216 = img_reg_array_11_43_real;
        _zz_217 = img_reg_array_11_43_imag;
        _zz_218 = img_reg_array_12_43_real;
        _zz_219 = img_reg_array_12_43_imag;
        _zz_220 = img_reg_array_13_43_real;
        _zz_221 = img_reg_array_13_43_imag;
        _zz_222 = img_reg_array_14_43_real;
        _zz_223 = img_reg_array_14_43_imag;
        _zz_224 = img_reg_array_15_43_real;
        _zz_225 = img_reg_array_15_43_imag;
        _zz_226 = img_reg_array_16_43_real;
        _zz_227 = img_reg_array_16_43_imag;
        _zz_228 = img_reg_array_17_43_real;
        _zz_229 = img_reg_array_17_43_imag;
        _zz_230 = img_reg_array_18_43_real;
        _zz_231 = img_reg_array_18_43_imag;
        _zz_232 = img_reg_array_19_43_real;
        _zz_233 = img_reg_array_19_43_imag;
        _zz_234 = img_reg_array_20_43_real;
        _zz_235 = img_reg_array_20_43_imag;
        _zz_236 = img_reg_array_21_43_real;
        _zz_237 = img_reg_array_21_43_imag;
        _zz_238 = img_reg_array_22_43_real;
        _zz_239 = img_reg_array_22_43_imag;
        _zz_240 = img_reg_array_23_43_real;
        _zz_241 = img_reg_array_23_43_imag;
        _zz_242 = img_reg_array_24_43_real;
        _zz_243 = img_reg_array_24_43_imag;
        _zz_244 = img_reg_array_25_43_real;
        _zz_245 = img_reg_array_25_43_imag;
        _zz_246 = img_reg_array_26_43_real;
        _zz_247 = img_reg_array_26_43_imag;
        _zz_248 = img_reg_array_27_43_real;
        _zz_249 = img_reg_array_27_43_imag;
        _zz_250 = img_reg_array_28_43_real;
        _zz_251 = img_reg_array_28_43_imag;
        _zz_252 = img_reg_array_29_43_real;
        _zz_253 = img_reg_array_29_43_imag;
        _zz_254 = img_reg_array_30_43_real;
        _zz_255 = img_reg_array_30_43_imag;
        _zz_256 = img_reg_array_31_43_real;
        _zz_257 = img_reg_array_31_43_imag;
        _zz_258 = img_reg_array_32_43_real;
        _zz_259 = img_reg_array_32_43_imag;
        _zz_260 = img_reg_array_33_43_real;
        _zz_261 = img_reg_array_33_43_imag;
        _zz_262 = img_reg_array_34_43_real;
        _zz_263 = img_reg_array_34_43_imag;
        _zz_264 = img_reg_array_35_43_real;
        _zz_265 = img_reg_array_35_43_imag;
        _zz_266 = img_reg_array_36_43_real;
        _zz_267 = img_reg_array_36_43_imag;
        _zz_268 = img_reg_array_37_43_real;
        _zz_269 = img_reg_array_37_43_imag;
        _zz_270 = img_reg_array_38_43_real;
        _zz_271 = img_reg_array_38_43_imag;
        _zz_272 = img_reg_array_39_43_real;
        _zz_273 = img_reg_array_39_43_imag;
        _zz_274 = img_reg_array_40_43_real;
        _zz_275 = img_reg_array_40_43_imag;
        _zz_276 = img_reg_array_41_43_real;
        _zz_277 = img_reg_array_41_43_imag;
        _zz_278 = img_reg_array_42_43_real;
        _zz_279 = img_reg_array_42_43_imag;
        _zz_280 = img_reg_array_43_43_real;
        _zz_281 = img_reg_array_43_43_imag;
        _zz_282 = img_reg_array_44_43_real;
        _zz_283 = img_reg_array_44_43_imag;
        _zz_284 = img_reg_array_45_43_real;
        _zz_285 = img_reg_array_45_43_imag;
        _zz_286 = img_reg_array_46_43_real;
        _zz_287 = img_reg_array_46_43_imag;
        _zz_288 = img_reg_array_47_43_real;
        _zz_289 = img_reg_array_47_43_imag;
        _zz_290 = img_reg_array_48_43_real;
        _zz_291 = img_reg_array_48_43_imag;
        _zz_292 = img_reg_array_49_43_real;
        _zz_293 = img_reg_array_49_43_imag;
        _zz_294 = img_reg_array_50_43_real;
        _zz_295 = img_reg_array_50_43_imag;
        _zz_296 = img_reg_array_51_43_real;
        _zz_297 = img_reg_array_51_43_imag;
        _zz_298 = img_reg_array_52_43_real;
        _zz_299 = img_reg_array_52_43_imag;
        _zz_300 = img_reg_array_53_43_real;
        _zz_301 = img_reg_array_53_43_imag;
        _zz_302 = img_reg_array_54_43_real;
        _zz_303 = img_reg_array_54_43_imag;
        _zz_304 = img_reg_array_55_43_real;
        _zz_305 = img_reg_array_55_43_imag;
        _zz_306 = img_reg_array_56_43_real;
        _zz_307 = img_reg_array_56_43_imag;
        _zz_308 = img_reg_array_57_43_real;
        _zz_309 = img_reg_array_57_43_imag;
        _zz_310 = img_reg_array_58_43_real;
        _zz_311 = img_reg_array_58_43_imag;
        _zz_312 = img_reg_array_59_43_real;
        _zz_313 = img_reg_array_59_43_imag;
        _zz_314 = img_reg_array_60_43_real;
        _zz_315 = img_reg_array_60_43_imag;
        _zz_316 = img_reg_array_61_43_real;
        _zz_317 = img_reg_array_61_43_imag;
        _zz_318 = img_reg_array_62_43_real;
        _zz_319 = img_reg_array_62_43_imag;
        _zz_320 = img_reg_array_63_43_real;
        _zz_321 = img_reg_array_63_43_imag;
      end
      6'b101100 : begin
        _zz_194 = img_reg_array_0_44_real;
        _zz_195 = img_reg_array_0_44_imag;
        _zz_196 = img_reg_array_1_44_real;
        _zz_197 = img_reg_array_1_44_imag;
        _zz_198 = img_reg_array_2_44_real;
        _zz_199 = img_reg_array_2_44_imag;
        _zz_200 = img_reg_array_3_44_real;
        _zz_201 = img_reg_array_3_44_imag;
        _zz_202 = img_reg_array_4_44_real;
        _zz_203 = img_reg_array_4_44_imag;
        _zz_204 = img_reg_array_5_44_real;
        _zz_205 = img_reg_array_5_44_imag;
        _zz_206 = img_reg_array_6_44_real;
        _zz_207 = img_reg_array_6_44_imag;
        _zz_208 = img_reg_array_7_44_real;
        _zz_209 = img_reg_array_7_44_imag;
        _zz_210 = img_reg_array_8_44_real;
        _zz_211 = img_reg_array_8_44_imag;
        _zz_212 = img_reg_array_9_44_real;
        _zz_213 = img_reg_array_9_44_imag;
        _zz_214 = img_reg_array_10_44_real;
        _zz_215 = img_reg_array_10_44_imag;
        _zz_216 = img_reg_array_11_44_real;
        _zz_217 = img_reg_array_11_44_imag;
        _zz_218 = img_reg_array_12_44_real;
        _zz_219 = img_reg_array_12_44_imag;
        _zz_220 = img_reg_array_13_44_real;
        _zz_221 = img_reg_array_13_44_imag;
        _zz_222 = img_reg_array_14_44_real;
        _zz_223 = img_reg_array_14_44_imag;
        _zz_224 = img_reg_array_15_44_real;
        _zz_225 = img_reg_array_15_44_imag;
        _zz_226 = img_reg_array_16_44_real;
        _zz_227 = img_reg_array_16_44_imag;
        _zz_228 = img_reg_array_17_44_real;
        _zz_229 = img_reg_array_17_44_imag;
        _zz_230 = img_reg_array_18_44_real;
        _zz_231 = img_reg_array_18_44_imag;
        _zz_232 = img_reg_array_19_44_real;
        _zz_233 = img_reg_array_19_44_imag;
        _zz_234 = img_reg_array_20_44_real;
        _zz_235 = img_reg_array_20_44_imag;
        _zz_236 = img_reg_array_21_44_real;
        _zz_237 = img_reg_array_21_44_imag;
        _zz_238 = img_reg_array_22_44_real;
        _zz_239 = img_reg_array_22_44_imag;
        _zz_240 = img_reg_array_23_44_real;
        _zz_241 = img_reg_array_23_44_imag;
        _zz_242 = img_reg_array_24_44_real;
        _zz_243 = img_reg_array_24_44_imag;
        _zz_244 = img_reg_array_25_44_real;
        _zz_245 = img_reg_array_25_44_imag;
        _zz_246 = img_reg_array_26_44_real;
        _zz_247 = img_reg_array_26_44_imag;
        _zz_248 = img_reg_array_27_44_real;
        _zz_249 = img_reg_array_27_44_imag;
        _zz_250 = img_reg_array_28_44_real;
        _zz_251 = img_reg_array_28_44_imag;
        _zz_252 = img_reg_array_29_44_real;
        _zz_253 = img_reg_array_29_44_imag;
        _zz_254 = img_reg_array_30_44_real;
        _zz_255 = img_reg_array_30_44_imag;
        _zz_256 = img_reg_array_31_44_real;
        _zz_257 = img_reg_array_31_44_imag;
        _zz_258 = img_reg_array_32_44_real;
        _zz_259 = img_reg_array_32_44_imag;
        _zz_260 = img_reg_array_33_44_real;
        _zz_261 = img_reg_array_33_44_imag;
        _zz_262 = img_reg_array_34_44_real;
        _zz_263 = img_reg_array_34_44_imag;
        _zz_264 = img_reg_array_35_44_real;
        _zz_265 = img_reg_array_35_44_imag;
        _zz_266 = img_reg_array_36_44_real;
        _zz_267 = img_reg_array_36_44_imag;
        _zz_268 = img_reg_array_37_44_real;
        _zz_269 = img_reg_array_37_44_imag;
        _zz_270 = img_reg_array_38_44_real;
        _zz_271 = img_reg_array_38_44_imag;
        _zz_272 = img_reg_array_39_44_real;
        _zz_273 = img_reg_array_39_44_imag;
        _zz_274 = img_reg_array_40_44_real;
        _zz_275 = img_reg_array_40_44_imag;
        _zz_276 = img_reg_array_41_44_real;
        _zz_277 = img_reg_array_41_44_imag;
        _zz_278 = img_reg_array_42_44_real;
        _zz_279 = img_reg_array_42_44_imag;
        _zz_280 = img_reg_array_43_44_real;
        _zz_281 = img_reg_array_43_44_imag;
        _zz_282 = img_reg_array_44_44_real;
        _zz_283 = img_reg_array_44_44_imag;
        _zz_284 = img_reg_array_45_44_real;
        _zz_285 = img_reg_array_45_44_imag;
        _zz_286 = img_reg_array_46_44_real;
        _zz_287 = img_reg_array_46_44_imag;
        _zz_288 = img_reg_array_47_44_real;
        _zz_289 = img_reg_array_47_44_imag;
        _zz_290 = img_reg_array_48_44_real;
        _zz_291 = img_reg_array_48_44_imag;
        _zz_292 = img_reg_array_49_44_real;
        _zz_293 = img_reg_array_49_44_imag;
        _zz_294 = img_reg_array_50_44_real;
        _zz_295 = img_reg_array_50_44_imag;
        _zz_296 = img_reg_array_51_44_real;
        _zz_297 = img_reg_array_51_44_imag;
        _zz_298 = img_reg_array_52_44_real;
        _zz_299 = img_reg_array_52_44_imag;
        _zz_300 = img_reg_array_53_44_real;
        _zz_301 = img_reg_array_53_44_imag;
        _zz_302 = img_reg_array_54_44_real;
        _zz_303 = img_reg_array_54_44_imag;
        _zz_304 = img_reg_array_55_44_real;
        _zz_305 = img_reg_array_55_44_imag;
        _zz_306 = img_reg_array_56_44_real;
        _zz_307 = img_reg_array_56_44_imag;
        _zz_308 = img_reg_array_57_44_real;
        _zz_309 = img_reg_array_57_44_imag;
        _zz_310 = img_reg_array_58_44_real;
        _zz_311 = img_reg_array_58_44_imag;
        _zz_312 = img_reg_array_59_44_real;
        _zz_313 = img_reg_array_59_44_imag;
        _zz_314 = img_reg_array_60_44_real;
        _zz_315 = img_reg_array_60_44_imag;
        _zz_316 = img_reg_array_61_44_real;
        _zz_317 = img_reg_array_61_44_imag;
        _zz_318 = img_reg_array_62_44_real;
        _zz_319 = img_reg_array_62_44_imag;
        _zz_320 = img_reg_array_63_44_real;
        _zz_321 = img_reg_array_63_44_imag;
      end
      6'b101101 : begin
        _zz_194 = img_reg_array_0_45_real;
        _zz_195 = img_reg_array_0_45_imag;
        _zz_196 = img_reg_array_1_45_real;
        _zz_197 = img_reg_array_1_45_imag;
        _zz_198 = img_reg_array_2_45_real;
        _zz_199 = img_reg_array_2_45_imag;
        _zz_200 = img_reg_array_3_45_real;
        _zz_201 = img_reg_array_3_45_imag;
        _zz_202 = img_reg_array_4_45_real;
        _zz_203 = img_reg_array_4_45_imag;
        _zz_204 = img_reg_array_5_45_real;
        _zz_205 = img_reg_array_5_45_imag;
        _zz_206 = img_reg_array_6_45_real;
        _zz_207 = img_reg_array_6_45_imag;
        _zz_208 = img_reg_array_7_45_real;
        _zz_209 = img_reg_array_7_45_imag;
        _zz_210 = img_reg_array_8_45_real;
        _zz_211 = img_reg_array_8_45_imag;
        _zz_212 = img_reg_array_9_45_real;
        _zz_213 = img_reg_array_9_45_imag;
        _zz_214 = img_reg_array_10_45_real;
        _zz_215 = img_reg_array_10_45_imag;
        _zz_216 = img_reg_array_11_45_real;
        _zz_217 = img_reg_array_11_45_imag;
        _zz_218 = img_reg_array_12_45_real;
        _zz_219 = img_reg_array_12_45_imag;
        _zz_220 = img_reg_array_13_45_real;
        _zz_221 = img_reg_array_13_45_imag;
        _zz_222 = img_reg_array_14_45_real;
        _zz_223 = img_reg_array_14_45_imag;
        _zz_224 = img_reg_array_15_45_real;
        _zz_225 = img_reg_array_15_45_imag;
        _zz_226 = img_reg_array_16_45_real;
        _zz_227 = img_reg_array_16_45_imag;
        _zz_228 = img_reg_array_17_45_real;
        _zz_229 = img_reg_array_17_45_imag;
        _zz_230 = img_reg_array_18_45_real;
        _zz_231 = img_reg_array_18_45_imag;
        _zz_232 = img_reg_array_19_45_real;
        _zz_233 = img_reg_array_19_45_imag;
        _zz_234 = img_reg_array_20_45_real;
        _zz_235 = img_reg_array_20_45_imag;
        _zz_236 = img_reg_array_21_45_real;
        _zz_237 = img_reg_array_21_45_imag;
        _zz_238 = img_reg_array_22_45_real;
        _zz_239 = img_reg_array_22_45_imag;
        _zz_240 = img_reg_array_23_45_real;
        _zz_241 = img_reg_array_23_45_imag;
        _zz_242 = img_reg_array_24_45_real;
        _zz_243 = img_reg_array_24_45_imag;
        _zz_244 = img_reg_array_25_45_real;
        _zz_245 = img_reg_array_25_45_imag;
        _zz_246 = img_reg_array_26_45_real;
        _zz_247 = img_reg_array_26_45_imag;
        _zz_248 = img_reg_array_27_45_real;
        _zz_249 = img_reg_array_27_45_imag;
        _zz_250 = img_reg_array_28_45_real;
        _zz_251 = img_reg_array_28_45_imag;
        _zz_252 = img_reg_array_29_45_real;
        _zz_253 = img_reg_array_29_45_imag;
        _zz_254 = img_reg_array_30_45_real;
        _zz_255 = img_reg_array_30_45_imag;
        _zz_256 = img_reg_array_31_45_real;
        _zz_257 = img_reg_array_31_45_imag;
        _zz_258 = img_reg_array_32_45_real;
        _zz_259 = img_reg_array_32_45_imag;
        _zz_260 = img_reg_array_33_45_real;
        _zz_261 = img_reg_array_33_45_imag;
        _zz_262 = img_reg_array_34_45_real;
        _zz_263 = img_reg_array_34_45_imag;
        _zz_264 = img_reg_array_35_45_real;
        _zz_265 = img_reg_array_35_45_imag;
        _zz_266 = img_reg_array_36_45_real;
        _zz_267 = img_reg_array_36_45_imag;
        _zz_268 = img_reg_array_37_45_real;
        _zz_269 = img_reg_array_37_45_imag;
        _zz_270 = img_reg_array_38_45_real;
        _zz_271 = img_reg_array_38_45_imag;
        _zz_272 = img_reg_array_39_45_real;
        _zz_273 = img_reg_array_39_45_imag;
        _zz_274 = img_reg_array_40_45_real;
        _zz_275 = img_reg_array_40_45_imag;
        _zz_276 = img_reg_array_41_45_real;
        _zz_277 = img_reg_array_41_45_imag;
        _zz_278 = img_reg_array_42_45_real;
        _zz_279 = img_reg_array_42_45_imag;
        _zz_280 = img_reg_array_43_45_real;
        _zz_281 = img_reg_array_43_45_imag;
        _zz_282 = img_reg_array_44_45_real;
        _zz_283 = img_reg_array_44_45_imag;
        _zz_284 = img_reg_array_45_45_real;
        _zz_285 = img_reg_array_45_45_imag;
        _zz_286 = img_reg_array_46_45_real;
        _zz_287 = img_reg_array_46_45_imag;
        _zz_288 = img_reg_array_47_45_real;
        _zz_289 = img_reg_array_47_45_imag;
        _zz_290 = img_reg_array_48_45_real;
        _zz_291 = img_reg_array_48_45_imag;
        _zz_292 = img_reg_array_49_45_real;
        _zz_293 = img_reg_array_49_45_imag;
        _zz_294 = img_reg_array_50_45_real;
        _zz_295 = img_reg_array_50_45_imag;
        _zz_296 = img_reg_array_51_45_real;
        _zz_297 = img_reg_array_51_45_imag;
        _zz_298 = img_reg_array_52_45_real;
        _zz_299 = img_reg_array_52_45_imag;
        _zz_300 = img_reg_array_53_45_real;
        _zz_301 = img_reg_array_53_45_imag;
        _zz_302 = img_reg_array_54_45_real;
        _zz_303 = img_reg_array_54_45_imag;
        _zz_304 = img_reg_array_55_45_real;
        _zz_305 = img_reg_array_55_45_imag;
        _zz_306 = img_reg_array_56_45_real;
        _zz_307 = img_reg_array_56_45_imag;
        _zz_308 = img_reg_array_57_45_real;
        _zz_309 = img_reg_array_57_45_imag;
        _zz_310 = img_reg_array_58_45_real;
        _zz_311 = img_reg_array_58_45_imag;
        _zz_312 = img_reg_array_59_45_real;
        _zz_313 = img_reg_array_59_45_imag;
        _zz_314 = img_reg_array_60_45_real;
        _zz_315 = img_reg_array_60_45_imag;
        _zz_316 = img_reg_array_61_45_real;
        _zz_317 = img_reg_array_61_45_imag;
        _zz_318 = img_reg_array_62_45_real;
        _zz_319 = img_reg_array_62_45_imag;
        _zz_320 = img_reg_array_63_45_real;
        _zz_321 = img_reg_array_63_45_imag;
      end
      6'b101110 : begin
        _zz_194 = img_reg_array_0_46_real;
        _zz_195 = img_reg_array_0_46_imag;
        _zz_196 = img_reg_array_1_46_real;
        _zz_197 = img_reg_array_1_46_imag;
        _zz_198 = img_reg_array_2_46_real;
        _zz_199 = img_reg_array_2_46_imag;
        _zz_200 = img_reg_array_3_46_real;
        _zz_201 = img_reg_array_3_46_imag;
        _zz_202 = img_reg_array_4_46_real;
        _zz_203 = img_reg_array_4_46_imag;
        _zz_204 = img_reg_array_5_46_real;
        _zz_205 = img_reg_array_5_46_imag;
        _zz_206 = img_reg_array_6_46_real;
        _zz_207 = img_reg_array_6_46_imag;
        _zz_208 = img_reg_array_7_46_real;
        _zz_209 = img_reg_array_7_46_imag;
        _zz_210 = img_reg_array_8_46_real;
        _zz_211 = img_reg_array_8_46_imag;
        _zz_212 = img_reg_array_9_46_real;
        _zz_213 = img_reg_array_9_46_imag;
        _zz_214 = img_reg_array_10_46_real;
        _zz_215 = img_reg_array_10_46_imag;
        _zz_216 = img_reg_array_11_46_real;
        _zz_217 = img_reg_array_11_46_imag;
        _zz_218 = img_reg_array_12_46_real;
        _zz_219 = img_reg_array_12_46_imag;
        _zz_220 = img_reg_array_13_46_real;
        _zz_221 = img_reg_array_13_46_imag;
        _zz_222 = img_reg_array_14_46_real;
        _zz_223 = img_reg_array_14_46_imag;
        _zz_224 = img_reg_array_15_46_real;
        _zz_225 = img_reg_array_15_46_imag;
        _zz_226 = img_reg_array_16_46_real;
        _zz_227 = img_reg_array_16_46_imag;
        _zz_228 = img_reg_array_17_46_real;
        _zz_229 = img_reg_array_17_46_imag;
        _zz_230 = img_reg_array_18_46_real;
        _zz_231 = img_reg_array_18_46_imag;
        _zz_232 = img_reg_array_19_46_real;
        _zz_233 = img_reg_array_19_46_imag;
        _zz_234 = img_reg_array_20_46_real;
        _zz_235 = img_reg_array_20_46_imag;
        _zz_236 = img_reg_array_21_46_real;
        _zz_237 = img_reg_array_21_46_imag;
        _zz_238 = img_reg_array_22_46_real;
        _zz_239 = img_reg_array_22_46_imag;
        _zz_240 = img_reg_array_23_46_real;
        _zz_241 = img_reg_array_23_46_imag;
        _zz_242 = img_reg_array_24_46_real;
        _zz_243 = img_reg_array_24_46_imag;
        _zz_244 = img_reg_array_25_46_real;
        _zz_245 = img_reg_array_25_46_imag;
        _zz_246 = img_reg_array_26_46_real;
        _zz_247 = img_reg_array_26_46_imag;
        _zz_248 = img_reg_array_27_46_real;
        _zz_249 = img_reg_array_27_46_imag;
        _zz_250 = img_reg_array_28_46_real;
        _zz_251 = img_reg_array_28_46_imag;
        _zz_252 = img_reg_array_29_46_real;
        _zz_253 = img_reg_array_29_46_imag;
        _zz_254 = img_reg_array_30_46_real;
        _zz_255 = img_reg_array_30_46_imag;
        _zz_256 = img_reg_array_31_46_real;
        _zz_257 = img_reg_array_31_46_imag;
        _zz_258 = img_reg_array_32_46_real;
        _zz_259 = img_reg_array_32_46_imag;
        _zz_260 = img_reg_array_33_46_real;
        _zz_261 = img_reg_array_33_46_imag;
        _zz_262 = img_reg_array_34_46_real;
        _zz_263 = img_reg_array_34_46_imag;
        _zz_264 = img_reg_array_35_46_real;
        _zz_265 = img_reg_array_35_46_imag;
        _zz_266 = img_reg_array_36_46_real;
        _zz_267 = img_reg_array_36_46_imag;
        _zz_268 = img_reg_array_37_46_real;
        _zz_269 = img_reg_array_37_46_imag;
        _zz_270 = img_reg_array_38_46_real;
        _zz_271 = img_reg_array_38_46_imag;
        _zz_272 = img_reg_array_39_46_real;
        _zz_273 = img_reg_array_39_46_imag;
        _zz_274 = img_reg_array_40_46_real;
        _zz_275 = img_reg_array_40_46_imag;
        _zz_276 = img_reg_array_41_46_real;
        _zz_277 = img_reg_array_41_46_imag;
        _zz_278 = img_reg_array_42_46_real;
        _zz_279 = img_reg_array_42_46_imag;
        _zz_280 = img_reg_array_43_46_real;
        _zz_281 = img_reg_array_43_46_imag;
        _zz_282 = img_reg_array_44_46_real;
        _zz_283 = img_reg_array_44_46_imag;
        _zz_284 = img_reg_array_45_46_real;
        _zz_285 = img_reg_array_45_46_imag;
        _zz_286 = img_reg_array_46_46_real;
        _zz_287 = img_reg_array_46_46_imag;
        _zz_288 = img_reg_array_47_46_real;
        _zz_289 = img_reg_array_47_46_imag;
        _zz_290 = img_reg_array_48_46_real;
        _zz_291 = img_reg_array_48_46_imag;
        _zz_292 = img_reg_array_49_46_real;
        _zz_293 = img_reg_array_49_46_imag;
        _zz_294 = img_reg_array_50_46_real;
        _zz_295 = img_reg_array_50_46_imag;
        _zz_296 = img_reg_array_51_46_real;
        _zz_297 = img_reg_array_51_46_imag;
        _zz_298 = img_reg_array_52_46_real;
        _zz_299 = img_reg_array_52_46_imag;
        _zz_300 = img_reg_array_53_46_real;
        _zz_301 = img_reg_array_53_46_imag;
        _zz_302 = img_reg_array_54_46_real;
        _zz_303 = img_reg_array_54_46_imag;
        _zz_304 = img_reg_array_55_46_real;
        _zz_305 = img_reg_array_55_46_imag;
        _zz_306 = img_reg_array_56_46_real;
        _zz_307 = img_reg_array_56_46_imag;
        _zz_308 = img_reg_array_57_46_real;
        _zz_309 = img_reg_array_57_46_imag;
        _zz_310 = img_reg_array_58_46_real;
        _zz_311 = img_reg_array_58_46_imag;
        _zz_312 = img_reg_array_59_46_real;
        _zz_313 = img_reg_array_59_46_imag;
        _zz_314 = img_reg_array_60_46_real;
        _zz_315 = img_reg_array_60_46_imag;
        _zz_316 = img_reg_array_61_46_real;
        _zz_317 = img_reg_array_61_46_imag;
        _zz_318 = img_reg_array_62_46_real;
        _zz_319 = img_reg_array_62_46_imag;
        _zz_320 = img_reg_array_63_46_real;
        _zz_321 = img_reg_array_63_46_imag;
      end
      6'b101111 : begin
        _zz_194 = img_reg_array_0_47_real;
        _zz_195 = img_reg_array_0_47_imag;
        _zz_196 = img_reg_array_1_47_real;
        _zz_197 = img_reg_array_1_47_imag;
        _zz_198 = img_reg_array_2_47_real;
        _zz_199 = img_reg_array_2_47_imag;
        _zz_200 = img_reg_array_3_47_real;
        _zz_201 = img_reg_array_3_47_imag;
        _zz_202 = img_reg_array_4_47_real;
        _zz_203 = img_reg_array_4_47_imag;
        _zz_204 = img_reg_array_5_47_real;
        _zz_205 = img_reg_array_5_47_imag;
        _zz_206 = img_reg_array_6_47_real;
        _zz_207 = img_reg_array_6_47_imag;
        _zz_208 = img_reg_array_7_47_real;
        _zz_209 = img_reg_array_7_47_imag;
        _zz_210 = img_reg_array_8_47_real;
        _zz_211 = img_reg_array_8_47_imag;
        _zz_212 = img_reg_array_9_47_real;
        _zz_213 = img_reg_array_9_47_imag;
        _zz_214 = img_reg_array_10_47_real;
        _zz_215 = img_reg_array_10_47_imag;
        _zz_216 = img_reg_array_11_47_real;
        _zz_217 = img_reg_array_11_47_imag;
        _zz_218 = img_reg_array_12_47_real;
        _zz_219 = img_reg_array_12_47_imag;
        _zz_220 = img_reg_array_13_47_real;
        _zz_221 = img_reg_array_13_47_imag;
        _zz_222 = img_reg_array_14_47_real;
        _zz_223 = img_reg_array_14_47_imag;
        _zz_224 = img_reg_array_15_47_real;
        _zz_225 = img_reg_array_15_47_imag;
        _zz_226 = img_reg_array_16_47_real;
        _zz_227 = img_reg_array_16_47_imag;
        _zz_228 = img_reg_array_17_47_real;
        _zz_229 = img_reg_array_17_47_imag;
        _zz_230 = img_reg_array_18_47_real;
        _zz_231 = img_reg_array_18_47_imag;
        _zz_232 = img_reg_array_19_47_real;
        _zz_233 = img_reg_array_19_47_imag;
        _zz_234 = img_reg_array_20_47_real;
        _zz_235 = img_reg_array_20_47_imag;
        _zz_236 = img_reg_array_21_47_real;
        _zz_237 = img_reg_array_21_47_imag;
        _zz_238 = img_reg_array_22_47_real;
        _zz_239 = img_reg_array_22_47_imag;
        _zz_240 = img_reg_array_23_47_real;
        _zz_241 = img_reg_array_23_47_imag;
        _zz_242 = img_reg_array_24_47_real;
        _zz_243 = img_reg_array_24_47_imag;
        _zz_244 = img_reg_array_25_47_real;
        _zz_245 = img_reg_array_25_47_imag;
        _zz_246 = img_reg_array_26_47_real;
        _zz_247 = img_reg_array_26_47_imag;
        _zz_248 = img_reg_array_27_47_real;
        _zz_249 = img_reg_array_27_47_imag;
        _zz_250 = img_reg_array_28_47_real;
        _zz_251 = img_reg_array_28_47_imag;
        _zz_252 = img_reg_array_29_47_real;
        _zz_253 = img_reg_array_29_47_imag;
        _zz_254 = img_reg_array_30_47_real;
        _zz_255 = img_reg_array_30_47_imag;
        _zz_256 = img_reg_array_31_47_real;
        _zz_257 = img_reg_array_31_47_imag;
        _zz_258 = img_reg_array_32_47_real;
        _zz_259 = img_reg_array_32_47_imag;
        _zz_260 = img_reg_array_33_47_real;
        _zz_261 = img_reg_array_33_47_imag;
        _zz_262 = img_reg_array_34_47_real;
        _zz_263 = img_reg_array_34_47_imag;
        _zz_264 = img_reg_array_35_47_real;
        _zz_265 = img_reg_array_35_47_imag;
        _zz_266 = img_reg_array_36_47_real;
        _zz_267 = img_reg_array_36_47_imag;
        _zz_268 = img_reg_array_37_47_real;
        _zz_269 = img_reg_array_37_47_imag;
        _zz_270 = img_reg_array_38_47_real;
        _zz_271 = img_reg_array_38_47_imag;
        _zz_272 = img_reg_array_39_47_real;
        _zz_273 = img_reg_array_39_47_imag;
        _zz_274 = img_reg_array_40_47_real;
        _zz_275 = img_reg_array_40_47_imag;
        _zz_276 = img_reg_array_41_47_real;
        _zz_277 = img_reg_array_41_47_imag;
        _zz_278 = img_reg_array_42_47_real;
        _zz_279 = img_reg_array_42_47_imag;
        _zz_280 = img_reg_array_43_47_real;
        _zz_281 = img_reg_array_43_47_imag;
        _zz_282 = img_reg_array_44_47_real;
        _zz_283 = img_reg_array_44_47_imag;
        _zz_284 = img_reg_array_45_47_real;
        _zz_285 = img_reg_array_45_47_imag;
        _zz_286 = img_reg_array_46_47_real;
        _zz_287 = img_reg_array_46_47_imag;
        _zz_288 = img_reg_array_47_47_real;
        _zz_289 = img_reg_array_47_47_imag;
        _zz_290 = img_reg_array_48_47_real;
        _zz_291 = img_reg_array_48_47_imag;
        _zz_292 = img_reg_array_49_47_real;
        _zz_293 = img_reg_array_49_47_imag;
        _zz_294 = img_reg_array_50_47_real;
        _zz_295 = img_reg_array_50_47_imag;
        _zz_296 = img_reg_array_51_47_real;
        _zz_297 = img_reg_array_51_47_imag;
        _zz_298 = img_reg_array_52_47_real;
        _zz_299 = img_reg_array_52_47_imag;
        _zz_300 = img_reg_array_53_47_real;
        _zz_301 = img_reg_array_53_47_imag;
        _zz_302 = img_reg_array_54_47_real;
        _zz_303 = img_reg_array_54_47_imag;
        _zz_304 = img_reg_array_55_47_real;
        _zz_305 = img_reg_array_55_47_imag;
        _zz_306 = img_reg_array_56_47_real;
        _zz_307 = img_reg_array_56_47_imag;
        _zz_308 = img_reg_array_57_47_real;
        _zz_309 = img_reg_array_57_47_imag;
        _zz_310 = img_reg_array_58_47_real;
        _zz_311 = img_reg_array_58_47_imag;
        _zz_312 = img_reg_array_59_47_real;
        _zz_313 = img_reg_array_59_47_imag;
        _zz_314 = img_reg_array_60_47_real;
        _zz_315 = img_reg_array_60_47_imag;
        _zz_316 = img_reg_array_61_47_real;
        _zz_317 = img_reg_array_61_47_imag;
        _zz_318 = img_reg_array_62_47_real;
        _zz_319 = img_reg_array_62_47_imag;
        _zz_320 = img_reg_array_63_47_real;
        _zz_321 = img_reg_array_63_47_imag;
      end
      6'b110000 : begin
        _zz_194 = img_reg_array_0_48_real;
        _zz_195 = img_reg_array_0_48_imag;
        _zz_196 = img_reg_array_1_48_real;
        _zz_197 = img_reg_array_1_48_imag;
        _zz_198 = img_reg_array_2_48_real;
        _zz_199 = img_reg_array_2_48_imag;
        _zz_200 = img_reg_array_3_48_real;
        _zz_201 = img_reg_array_3_48_imag;
        _zz_202 = img_reg_array_4_48_real;
        _zz_203 = img_reg_array_4_48_imag;
        _zz_204 = img_reg_array_5_48_real;
        _zz_205 = img_reg_array_5_48_imag;
        _zz_206 = img_reg_array_6_48_real;
        _zz_207 = img_reg_array_6_48_imag;
        _zz_208 = img_reg_array_7_48_real;
        _zz_209 = img_reg_array_7_48_imag;
        _zz_210 = img_reg_array_8_48_real;
        _zz_211 = img_reg_array_8_48_imag;
        _zz_212 = img_reg_array_9_48_real;
        _zz_213 = img_reg_array_9_48_imag;
        _zz_214 = img_reg_array_10_48_real;
        _zz_215 = img_reg_array_10_48_imag;
        _zz_216 = img_reg_array_11_48_real;
        _zz_217 = img_reg_array_11_48_imag;
        _zz_218 = img_reg_array_12_48_real;
        _zz_219 = img_reg_array_12_48_imag;
        _zz_220 = img_reg_array_13_48_real;
        _zz_221 = img_reg_array_13_48_imag;
        _zz_222 = img_reg_array_14_48_real;
        _zz_223 = img_reg_array_14_48_imag;
        _zz_224 = img_reg_array_15_48_real;
        _zz_225 = img_reg_array_15_48_imag;
        _zz_226 = img_reg_array_16_48_real;
        _zz_227 = img_reg_array_16_48_imag;
        _zz_228 = img_reg_array_17_48_real;
        _zz_229 = img_reg_array_17_48_imag;
        _zz_230 = img_reg_array_18_48_real;
        _zz_231 = img_reg_array_18_48_imag;
        _zz_232 = img_reg_array_19_48_real;
        _zz_233 = img_reg_array_19_48_imag;
        _zz_234 = img_reg_array_20_48_real;
        _zz_235 = img_reg_array_20_48_imag;
        _zz_236 = img_reg_array_21_48_real;
        _zz_237 = img_reg_array_21_48_imag;
        _zz_238 = img_reg_array_22_48_real;
        _zz_239 = img_reg_array_22_48_imag;
        _zz_240 = img_reg_array_23_48_real;
        _zz_241 = img_reg_array_23_48_imag;
        _zz_242 = img_reg_array_24_48_real;
        _zz_243 = img_reg_array_24_48_imag;
        _zz_244 = img_reg_array_25_48_real;
        _zz_245 = img_reg_array_25_48_imag;
        _zz_246 = img_reg_array_26_48_real;
        _zz_247 = img_reg_array_26_48_imag;
        _zz_248 = img_reg_array_27_48_real;
        _zz_249 = img_reg_array_27_48_imag;
        _zz_250 = img_reg_array_28_48_real;
        _zz_251 = img_reg_array_28_48_imag;
        _zz_252 = img_reg_array_29_48_real;
        _zz_253 = img_reg_array_29_48_imag;
        _zz_254 = img_reg_array_30_48_real;
        _zz_255 = img_reg_array_30_48_imag;
        _zz_256 = img_reg_array_31_48_real;
        _zz_257 = img_reg_array_31_48_imag;
        _zz_258 = img_reg_array_32_48_real;
        _zz_259 = img_reg_array_32_48_imag;
        _zz_260 = img_reg_array_33_48_real;
        _zz_261 = img_reg_array_33_48_imag;
        _zz_262 = img_reg_array_34_48_real;
        _zz_263 = img_reg_array_34_48_imag;
        _zz_264 = img_reg_array_35_48_real;
        _zz_265 = img_reg_array_35_48_imag;
        _zz_266 = img_reg_array_36_48_real;
        _zz_267 = img_reg_array_36_48_imag;
        _zz_268 = img_reg_array_37_48_real;
        _zz_269 = img_reg_array_37_48_imag;
        _zz_270 = img_reg_array_38_48_real;
        _zz_271 = img_reg_array_38_48_imag;
        _zz_272 = img_reg_array_39_48_real;
        _zz_273 = img_reg_array_39_48_imag;
        _zz_274 = img_reg_array_40_48_real;
        _zz_275 = img_reg_array_40_48_imag;
        _zz_276 = img_reg_array_41_48_real;
        _zz_277 = img_reg_array_41_48_imag;
        _zz_278 = img_reg_array_42_48_real;
        _zz_279 = img_reg_array_42_48_imag;
        _zz_280 = img_reg_array_43_48_real;
        _zz_281 = img_reg_array_43_48_imag;
        _zz_282 = img_reg_array_44_48_real;
        _zz_283 = img_reg_array_44_48_imag;
        _zz_284 = img_reg_array_45_48_real;
        _zz_285 = img_reg_array_45_48_imag;
        _zz_286 = img_reg_array_46_48_real;
        _zz_287 = img_reg_array_46_48_imag;
        _zz_288 = img_reg_array_47_48_real;
        _zz_289 = img_reg_array_47_48_imag;
        _zz_290 = img_reg_array_48_48_real;
        _zz_291 = img_reg_array_48_48_imag;
        _zz_292 = img_reg_array_49_48_real;
        _zz_293 = img_reg_array_49_48_imag;
        _zz_294 = img_reg_array_50_48_real;
        _zz_295 = img_reg_array_50_48_imag;
        _zz_296 = img_reg_array_51_48_real;
        _zz_297 = img_reg_array_51_48_imag;
        _zz_298 = img_reg_array_52_48_real;
        _zz_299 = img_reg_array_52_48_imag;
        _zz_300 = img_reg_array_53_48_real;
        _zz_301 = img_reg_array_53_48_imag;
        _zz_302 = img_reg_array_54_48_real;
        _zz_303 = img_reg_array_54_48_imag;
        _zz_304 = img_reg_array_55_48_real;
        _zz_305 = img_reg_array_55_48_imag;
        _zz_306 = img_reg_array_56_48_real;
        _zz_307 = img_reg_array_56_48_imag;
        _zz_308 = img_reg_array_57_48_real;
        _zz_309 = img_reg_array_57_48_imag;
        _zz_310 = img_reg_array_58_48_real;
        _zz_311 = img_reg_array_58_48_imag;
        _zz_312 = img_reg_array_59_48_real;
        _zz_313 = img_reg_array_59_48_imag;
        _zz_314 = img_reg_array_60_48_real;
        _zz_315 = img_reg_array_60_48_imag;
        _zz_316 = img_reg_array_61_48_real;
        _zz_317 = img_reg_array_61_48_imag;
        _zz_318 = img_reg_array_62_48_real;
        _zz_319 = img_reg_array_62_48_imag;
        _zz_320 = img_reg_array_63_48_real;
        _zz_321 = img_reg_array_63_48_imag;
      end
      6'b110001 : begin
        _zz_194 = img_reg_array_0_49_real;
        _zz_195 = img_reg_array_0_49_imag;
        _zz_196 = img_reg_array_1_49_real;
        _zz_197 = img_reg_array_1_49_imag;
        _zz_198 = img_reg_array_2_49_real;
        _zz_199 = img_reg_array_2_49_imag;
        _zz_200 = img_reg_array_3_49_real;
        _zz_201 = img_reg_array_3_49_imag;
        _zz_202 = img_reg_array_4_49_real;
        _zz_203 = img_reg_array_4_49_imag;
        _zz_204 = img_reg_array_5_49_real;
        _zz_205 = img_reg_array_5_49_imag;
        _zz_206 = img_reg_array_6_49_real;
        _zz_207 = img_reg_array_6_49_imag;
        _zz_208 = img_reg_array_7_49_real;
        _zz_209 = img_reg_array_7_49_imag;
        _zz_210 = img_reg_array_8_49_real;
        _zz_211 = img_reg_array_8_49_imag;
        _zz_212 = img_reg_array_9_49_real;
        _zz_213 = img_reg_array_9_49_imag;
        _zz_214 = img_reg_array_10_49_real;
        _zz_215 = img_reg_array_10_49_imag;
        _zz_216 = img_reg_array_11_49_real;
        _zz_217 = img_reg_array_11_49_imag;
        _zz_218 = img_reg_array_12_49_real;
        _zz_219 = img_reg_array_12_49_imag;
        _zz_220 = img_reg_array_13_49_real;
        _zz_221 = img_reg_array_13_49_imag;
        _zz_222 = img_reg_array_14_49_real;
        _zz_223 = img_reg_array_14_49_imag;
        _zz_224 = img_reg_array_15_49_real;
        _zz_225 = img_reg_array_15_49_imag;
        _zz_226 = img_reg_array_16_49_real;
        _zz_227 = img_reg_array_16_49_imag;
        _zz_228 = img_reg_array_17_49_real;
        _zz_229 = img_reg_array_17_49_imag;
        _zz_230 = img_reg_array_18_49_real;
        _zz_231 = img_reg_array_18_49_imag;
        _zz_232 = img_reg_array_19_49_real;
        _zz_233 = img_reg_array_19_49_imag;
        _zz_234 = img_reg_array_20_49_real;
        _zz_235 = img_reg_array_20_49_imag;
        _zz_236 = img_reg_array_21_49_real;
        _zz_237 = img_reg_array_21_49_imag;
        _zz_238 = img_reg_array_22_49_real;
        _zz_239 = img_reg_array_22_49_imag;
        _zz_240 = img_reg_array_23_49_real;
        _zz_241 = img_reg_array_23_49_imag;
        _zz_242 = img_reg_array_24_49_real;
        _zz_243 = img_reg_array_24_49_imag;
        _zz_244 = img_reg_array_25_49_real;
        _zz_245 = img_reg_array_25_49_imag;
        _zz_246 = img_reg_array_26_49_real;
        _zz_247 = img_reg_array_26_49_imag;
        _zz_248 = img_reg_array_27_49_real;
        _zz_249 = img_reg_array_27_49_imag;
        _zz_250 = img_reg_array_28_49_real;
        _zz_251 = img_reg_array_28_49_imag;
        _zz_252 = img_reg_array_29_49_real;
        _zz_253 = img_reg_array_29_49_imag;
        _zz_254 = img_reg_array_30_49_real;
        _zz_255 = img_reg_array_30_49_imag;
        _zz_256 = img_reg_array_31_49_real;
        _zz_257 = img_reg_array_31_49_imag;
        _zz_258 = img_reg_array_32_49_real;
        _zz_259 = img_reg_array_32_49_imag;
        _zz_260 = img_reg_array_33_49_real;
        _zz_261 = img_reg_array_33_49_imag;
        _zz_262 = img_reg_array_34_49_real;
        _zz_263 = img_reg_array_34_49_imag;
        _zz_264 = img_reg_array_35_49_real;
        _zz_265 = img_reg_array_35_49_imag;
        _zz_266 = img_reg_array_36_49_real;
        _zz_267 = img_reg_array_36_49_imag;
        _zz_268 = img_reg_array_37_49_real;
        _zz_269 = img_reg_array_37_49_imag;
        _zz_270 = img_reg_array_38_49_real;
        _zz_271 = img_reg_array_38_49_imag;
        _zz_272 = img_reg_array_39_49_real;
        _zz_273 = img_reg_array_39_49_imag;
        _zz_274 = img_reg_array_40_49_real;
        _zz_275 = img_reg_array_40_49_imag;
        _zz_276 = img_reg_array_41_49_real;
        _zz_277 = img_reg_array_41_49_imag;
        _zz_278 = img_reg_array_42_49_real;
        _zz_279 = img_reg_array_42_49_imag;
        _zz_280 = img_reg_array_43_49_real;
        _zz_281 = img_reg_array_43_49_imag;
        _zz_282 = img_reg_array_44_49_real;
        _zz_283 = img_reg_array_44_49_imag;
        _zz_284 = img_reg_array_45_49_real;
        _zz_285 = img_reg_array_45_49_imag;
        _zz_286 = img_reg_array_46_49_real;
        _zz_287 = img_reg_array_46_49_imag;
        _zz_288 = img_reg_array_47_49_real;
        _zz_289 = img_reg_array_47_49_imag;
        _zz_290 = img_reg_array_48_49_real;
        _zz_291 = img_reg_array_48_49_imag;
        _zz_292 = img_reg_array_49_49_real;
        _zz_293 = img_reg_array_49_49_imag;
        _zz_294 = img_reg_array_50_49_real;
        _zz_295 = img_reg_array_50_49_imag;
        _zz_296 = img_reg_array_51_49_real;
        _zz_297 = img_reg_array_51_49_imag;
        _zz_298 = img_reg_array_52_49_real;
        _zz_299 = img_reg_array_52_49_imag;
        _zz_300 = img_reg_array_53_49_real;
        _zz_301 = img_reg_array_53_49_imag;
        _zz_302 = img_reg_array_54_49_real;
        _zz_303 = img_reg_array_54_49_imag;
        _zz_304 = img_reg_array_55_49_real;
        _zz_305 = img_reg_array_55_49_imag;
        _zz_306 = img_reg_array_56_49_real;
        _zz_307 = img_reg_array_56_49_imag;
        _zz_308 = img_reg_array_57_49_real;
        _zz_309 = img_reg_array_57_49_imag;
        _zz_310 = img_reg_array_58_49_real;
        _zz_311 = img_reg_array_58_49_imag;
        _zz_312 = img_reg_array_59_49_real;
        _zz_313 = img_reg_array_59_49_imag;
        _zz_314 = img_reg_array_60_49_real;
        _zz_315 = img_reg_array_60_49_imag;
        _zz_316 = img_reg_array_61_49_real;
        _zz_317 = img_reg_array_61_49_imag;
        _zz_318 = img_reg_array_62_49_real;
        _zz_319 = img_reg_array_62_49_imag;
        _zz_320 = img_reg_array_63_49_real;
        _zz_321 = img_reg_array_63_49_imag;
      end
      6'b110010 : begin
        _zz_194 = img_reg_array_0_50_real;
        _zz_195 = img_reg_array_0_50_imag;
        _zz_196 = img_reg_array_1_50_real;
        _zz_197 = img_reg_array_1_50_imag;
        _zz_198 = img_reg_array_2_50_real;
        _zz_199 = img_reg_array_2_50_imag;
        _zz_200 = img_reg_array_3_50_real;
        _zz_201 = img_reg_array_3_50_imag;
        _zz_202 = img_reg_array_4_50_real;
        _zz_203 = img_reg_array_4_50_imag;
        _zz_204 = img_reg_array_5_50_real;
        _zz_205 = img_reg_array_5_50_imag;
        _zz_206 = img_reg_array_6_50_real;
        _zz_207 = img_reg_array_6_50_imag;
        _zz_208 = img_reg_array_7_50_real;
        _zz_209 = img_reg_array_7_50_imag;
        _zz_210 = img_reg_array_8_50_real;
        _zz_211 = img_reg_array_8_50_imag;
        _zz_212 = img_reg_array_9_50_real;
        _zz_213 = img_reg_array_9_50_imag;
        _zz_214 = img_reg_array_10_50_real;
        _zz_215 = img_reg_array_10_50_imag;
        _zz_216 = img_reg_array_11_50_real;
        _zz_217 = img_reg_array_11_50_imag;
        _zz_218 = img_reg_array_12_50_real;
        _zz_219 = img_reg_array_12_50_imag;
        _zz_220 = img_reg_array_13_50_real;
        _zz_221 = img_reg_array_13_50_imag;
        _zz_222 = img_reg_array_14_50_real;
        _zz_223 = img_reg_array_14_50_imag;
        _zz_224 = img_reg_array_15_50_real;
        _zz_225 = img_reg_array_15_50_imag;
        _zz_226 = img_reg_array_16_50_real;
        _zz_227 = img_reg_array_16_50_imag;
        _zz_228 = img_reg_array_17_50_real;
        _zz_229 = img_reg_array_17_50_imag;
        _zz_230 = img_reg_array_18_50_real;
        _zz_231 = img_reg_array_18_50_imag;
        _zz_232 = img_reg_array_19_50_real;
        _zz_233 = img_reg_array_19_50_imag;
        _zz_234 = img_reg_array_20_50_real;
        _zz_235 = img_reg_array_20_50_imag;
        _zz_236 = img_reg_array_21_50_real;
        _zz_237 = img_reg_array_21_50_imag;
        _zz_238 = img_reg_array_22_50_real;
        _zz_239 = img_reg_array_22_50_imag;
        _zz_240 = img_reg_array_23_50_real;
        _zz_241 = img_reg_array_23_50_imag;
        _zz_242 = img_reg_array_24_50_real;
        _zz_243 = img_reg_array_24_50_imag;
        _zz_244 = img_reg_array_25_50_real;
        _zz_245 = img_reg_array_25_50_imag;
        _zz_246 = img_reg_array_26_50_real;
        _zz_247 = img_reg_array_26_50_imag;
        _zz_248 = img_reg_array_27_50_real;
        _zz_249 = img_reg_array_27_50_imag;
        _zz_250 = img_reg_array_28_50_real;
        _zz_251 = img_reg_array_28_50_imag;
        _zz_252 = img_reg_array_29_50_real;
        _zz_253 = img_reg_array_29_50_imag;
        _zz_254 = img_reg_array_30_50_real;
        _zz_255 = img_reg_array_30_50_imag;
        _zz_256 = img_reg_array_31_50_real;
        _zz_257 = img_reg_array_31_50_imag;
        _zz_258 = img_reg_array_32_50_real;
        _zz_259 = img_reg_array_32_50_imag;
        _zz_260 = img_reg_array_33_50_real;
        _zz_261 = img_reg_array_33_50_imag;
        _zz_262 = img_reg_array_34_50_real;
        _zz_263 = img_reg_array_34_50_imag;
        _zz_264 = img_reg_array_35_50_real;
        _zz_265 = img_reg_array_35_50_imag;
        _zz_266 = img_reg_array_36_50_real;
        _zz_267 = img_reg_array_36_50_imag;
        _zz_268 = img_reg_array_37_50_real;
        _zz_269 = img_reg_array_37_50_imag;
        _zz_270 = img_reg_array_38_50_real;
        _zz_271 = img_reg_array_38_50_imag;
        _zz_272 = img_reg_array_39_50_real;
        _zz_273 = img_reg_array_39_50_imag;
        _zz_274 = img_reg_array_40_50_real;
        _zz_275 = img_reg_array_40_50_imag;
        _zz_276 = img_reg_array_41_50_real;
        _zz_277 = img_reg_array_41_50_imag;
        _zz_278 = img_reg_array_42_50_real;
        _zz_279 = img_reg_array_42_50_imag;
        _zz_280 = img_reg_array_43_50_real;
        _zz_281 = img_reg_array_43_50_imag;
        _zz_282 = img_reg_array_44_50_real;
        _zz_283 = img_reg_array_44_50_imag;
        _zz_284 = img_reg_array_45_50_real;
        _zz_285 = img_reg_array_45_50_imag;
        _zz_286 = img_reg_array_46_50_real;
        _zz_287 = img_reg_array_46_50_imag;
        _zz_288 = img_reg_array_47_50_real;
        _zz_289 = img_reg_array_47_50_imag;
        _zz_290 = img_reg_array_48_50_real;
        _zz_291 = img_reg_array_48_50_imag;
        _zz_292 = img_reg_array_49_50_real;
        _zz_293 = img_reg_array_49_50_imag;
        _zz_294 = img_reg_array_50_50_real;
        _zz_295 = img_reg_array_50_50_imag;
        _zz_296 = img_reg_array_51_50_real;
        _zz_297 = img_reg_array_51_50_imag;
        _zz_298 = img_reg_array_52_50_real;
        _zz_299 = img_reg_array_52_50_imag;
        _zz_300 = img_reg_array_53_50_real;
        _zz_301 = img_reg_array_53_50_imag;
        _zz_302 = img_reg_array_54_50_real;
        _zz_303 = img_reg_array_54_50_imag;
        _zz_304 = img_reg_array_55_50_real;
        _zz_305 = img_reg_array_55_50_imag;
        _zz_306 = img_reg_array_56_50_real;
        _zz_307 = img_reg_array_56_50_imag;
        _zz_308 = img_reg_array_57_50_real;
        _zz_309 = img_reg_array_57_50_imag;
        _zz_310 = img_reg_array_58_50_real;
        _zz_311 = img_reg_array_58_50_imag;
        _zz_312 = img_reg_array_59_50_real;
        _zz_313 = img_reg_array_59_50_imag;
        _zz_314 = img_reg_array_60_50_real;
        _zz_315 = img_reg_array_60_50_imag;
        _zz_316 = img_reg_array_61_50_real;
        _zz_317 = img_reg_array_61_50_imag;
        _zz_318 = img_reg_array_62_50_real;
        _zz_319 = img_reg_array_62_50_imag;
        _zz_320 = img_reg_array_63_50_real;
        _zz_321 = img_reg_array_63_50_imag;
      end
      6'b110011 : begin
        _zz_194 = img_reg_array_0_51_real;
        _zz_195 = img_reg_array_0_51_imag;
        _zz_196 = img_reg_array_1_51_real;
        _zz_197 = img_reg_array_1_51_imag;
        _zz_198 = img_reg_array_2_51_real;
        _zz_199 = img_reg_array_2_51_imag;
        _zz_200 = img_reg_array_3_51_real;
        _zz_201 = img_reg_array_3_51_imag;
        _zz_202 = img_reg_array_4_51_real;
        _zz_203 = img_reg_array_4_51_imag;
        _zz_204 = img_reg_array_5_51_real;
        _zz_205 = img_reg_array_5_51_imag;
        _zz_206 = img_reg_array_6_51_real;
        _zz_207 = img_reg_array_6_51_imag;
        _zz_208 = img_reg_array_7_51_real;
        _zz_209 = img_reg_array_7_51_imag;
        _zz_210 = img_reg_array_8_51_real;
        _zz_211 = img_reg_array_8_51_imag;
        _zz_212 = img_reg_array_9_51_real;
        _zz_213 = img_reg_array_9_51_imag;
        _zz_214 = img_reg_array_10_51_real;
        _zz_215 = img_reg_array_10_51_imag;
        _zz_216 = img_reg_array_11_51_real;
        _zz_217 = img_reg_array_11_51_imag;
        _zz_218 = img_reg_array_12_51_real;
        _zz_219 = img_reg_array_12_51_imag;
        _zz_220 = img_reg_array_13_51_real;
        _zz_221 = img_reg_array_13_51_imag;
        _zz_222 = img_reg_array_14_51_real;
        _zz_223 = img_reg_array_14_51_imag;
        _zz_224 = img_reg_array_15_51_real;
        _zz_225 = img_reg_array_15_51_imag;
        _zz_226 = img_reg_array_16_51_real;
        _zz_227 = img_reg_array_16_51_imag;
        _zz_228 = img_reg_array_17_51_real;
        _zz_229 = img_reg_array_17_51_imag;
        _zz_230 = img_reg_array_18_51_real;
        _zz_231 = img_reg_array_18_51_imag;
        _zz_232 = img_reg_array_19_51_real;
        _zz_233 = img_reg_array_19_51_imag;
        _zz_234 = img_reg_array_20_51_real;
        _zz_235 = img_reg_array_20_51_imag;
        _zz_236 = img_reg_array_21_51_real;
        _zz_237 = img_reg_array_21_51_imag;
        _zz_238 = img_reg_array_22_51_real;
        _zz_239 = img_reg_array_22_51_imag;
        _zz_240 = img_reg_array_23_51_real;
        _zz_241 = img_reg_array_23_51_imag;
        _zz_242 = img_reg_array_24_51_real;
        _zz_243 = img_reg_array_24_51_imag;
        _zz_244 = img_reg_array_25_51_real;
        _zz_245 = img_reg_array_25_51_imag;
        _zz_246 = img_reg_array_26_51_real;
        _zz_247 = img_reg_array_26_51_imag;
        _zz_248 = img_reg_array_27_51_real;
        _zz_249 = img_reg_array_27_51_imag;
        _zz_250 = img_reg_array_28_51_real;
        _zz_251 = img_reg_array_28_51_imag;
        _zz_252 = img_reg_array_29_51_real;
        _zz_253 = img_reg_array_29_51_imag;
        _zz_254 = img_reg_array_30_51_real;
        _zz_255 = img_reg_array_30_51_imag;
        _zz_256 = img_reg_array_31_51_real;
        _zz_257 = img_reg_array_31_51_imag;
        _zz_258 = img_reg_array_32_51_real;
        _zz_259 = img_reg_array_32_51_imag;
        _zz_260 = img_reg_array_33_51_real;
        _zz_261 = img_reg_array_33_51_imag;
        _zz_262 = img_reg_array_34_51_real;
        _zz_263 = img_reg_array_34_51_imag;
        _zz_264 = img_reg_array_35_51_real;
        _zz_265 = img_reg_array_35_51_imag;
        _zz_266 = img_reg_array_36_51_real;
        _zz_267 = img_reg_array_36_51_imag;
        _zz_268 = img_reg_array_37_51_real;
        _zz_269 = img_reg_array_37_51_imag;
        _zz_270 = img_reg_array_38_51_real;
        _zz_271 = img_reg_array_38_51_imag;
        _zz_272 = img_reg_array_39_51_real;
        _zz_273 = img_reg_array_39_51_imag;
        _zz_274 = img_reg_array_40_51_real;
        _zz_275 = img_reg_array_40_51_imag;
        _zz_276 = img_reg_array_41_51_real;
        _zz_277 = img_reg_array_41_51_imag;
        _zz_278 = img_reg_array_42_51_real;
        _zz_279 = img_reg_array_42_51_imag;
        _zz_280 = img_reg_array_43_51_real;
        _zz_281 = img_reg_array_43_51_imag;
        _zz_282 = img_reg_array_44_51_real;
        _zz_283 = img_reg_array_44_51_imag;
        _zz_284 = img_reg_array_45_51_real;
        _zz_285 = img_reg_array_45_51_imag;
        _zz_286 = img_reg_array_46_51_real;
        _zz_287 = img_reg_array_46_51_imag;
        _zz_288 = img_reg_array_47_51_real;
        _zz_289 = img_reg_array_47_51_imag;
        _zz_290 = img_reg_array_48_51_real;
        _zz_291 = img_reg_array_48_51_imag;
        _zz_292 = img_reg_array_49_51_real;
        _zz_293 = img_reg_array_49_51_imag;
        _zz_294 = img_reg_array_50_51_real;
        _zz_295 = img_reg_array_50_51_imag;
        _zz_296 = img_reg_array_51_51_real;
        _zz_297 = img_reg_array_51_51_imag;
        _zz_298 = img_reg_array_52_51_real;
        _zz_299 = img_reg_array_52_51_imag;
        _zz_300 = img_reg_array_53_51_real;
        _zz_301 = img_reg_array_53_51_imag;
        _zz_302 = img_reg_array_54_51_real;
        _zz_303 = img_reg_array_54_51_imag;
        _zz_304 = img_reg_array_55_51_real;
        _zz_305 = img_reg_array_55_51_imag;
        _zz_306 = img_reg_array_56_51_real;
        _zz_307 = img_reg_array_56_51_imag;
        _zz_308 = img_reg_array_57_51_real;
        _zz_309 = img_reg_array_57_51_imag;
        _zz_310 = img_reg_array_58_51_real;
        _zz_311 = img_reg_array_58_51_imag;
        _zz_312 = img_reg_array_59_51_real;
        _zz_313 = img_reg_array_59_51_imag;
        _zz_314 = img_reg_array_60_51_real;
        _zz_315 = img_reg_array_60_51_imag;
        _zz_316 = img_reg_array_61_51_real;
        _zz_317 = img_reg_array_61_51_imag;
        _zz_318 = img_reg_array_62_51_real;
        _zz_319 = img_reg_array_62_51_imag;
        _zz_320 = img_reg_array_63_51_real;
        _zz_321 = img_reg_array_63_51_imag;
      end
      6'b110100 : begin
        _zz_194 = img_reg_array_0_52_real;
        _zz_195 = img_reg_array_0_52_imag;
        _zz_196 = img_reg_array_1_52_real;
        _zz_197 = img_reg_array_1_52_imag;
        _zz_198 = img_reg_array_2_52_real;
        _zz_199 = img_reg_array_2_52_imag;
        _zz_200 = img_reg_array_3_52_real;
        _zz_201 = img_reg_array_3_52_imag;
        _zz_202 = img_reg_array_4_52_real;
        _zz_203 = img_reg_array_4_52_imag;
        _zz_204 = img_reg_array_5_52_real;
        _zz_205 = img_reg_array_5_52_imag;
        _zz_206 = img_reg_array_6_52_real;
        _zz_207 = img_reg_array_6_52_imag;
        _zz_208 = img_reg_array_7_52_real;
        _zz_209 = img_reg_array_7_52_imag;
        _zz_210 = img_reg_array_8_52_real;
        _zz_211 = img_reg_array_8_52_imag;
        _zz_212 = img_reg_array_9_52_real;
        _zz_213 = img_reg_array_9_52_imag;
        _zz_214 = img_reg_array_10_52_real;
        _zz_215 = img_reg_array_10_52_imag;
        _zz_216 = img_reg_array_11_52_real;
        _zz_217 = img_reg_array_11_52_imag;
        _zz_218 = img_reg_array_12_52_real;
        _zz_219 = img_reg_array_12_52_imag;
        _zz_220 = img_reg_array_13_52_real;
        _zz_221 = img_reg_array_13_52_imag;
        _zz_222 = img_reg_array_14_52_real;
        _zz_223 = img_reg_array_14_52_imag;
        _zz_224 = img_reg_array_15_52_real;
        _zz_225 = img_reg_array_15_52_imag;
        _zz_226 = img_reg_array_16_52_real;
        _zz_227 = img_reg_array_16_52_imag;
        _zz_228 = img_reg_array_17_52_real;
        _zz_229 = img_reg_array_17_52_imag;
        _zz_230 = img_reg_array_18_52_real;
        _zz_231 = img_reg_array_18_52_imag;
        _zz_232 = img_reg_array_19_52_real;
        _zz_233 = img_reg_array_19_52_imag;
        _zz_234 = img_reg_array_20_52_real;
        _zz_235 = img_reg_array_20_52_imag;
        _zz_236 = img_reg_array_21_52_real;
        _zz_237 = img_reg_array_21_52_imag;
        _zz_238 = img_reg_array_22_52_real;
        _zz_239 = img_reg_array_22_52_imag;
        _zz_240 = img_reg_array_23_52_real;
        _zz_241 = img_reg_array_23_52_imag;
        _zz_242 = img_reg_array_24_52_real;
        _zz_243 = img_reg_array_24_52_imag;
        _zz_244 = img_reg_array_25_52_real;
        _zz_245 = img_reg_array_25_52_imag;
        _zz_246 = img_reg_array_26_52_real;
        _zz_247 = img_reg_array_26_52_imag;
        _zz_248 = img_reg_array_27_52_real;
        _zz_249 = img_reg_array_27_52_imag;
        _zz_250 = img_reg_array_28_52_real;
        _zz_251 = img_reg_array_28_52_imag;
        _zz_252 = img_reg_array_29_52_real;
        _zz_253 = img_reg_array_29_52_imag;
        _zz_254 = img_reg_array_30_52_real;
        _zz_255 = img_reg_array_30_52_imag;
        _zz_256 = img_reg_array_31_52_real;
        _zz_257 = img_reg_array_31_52_imag;
        _zz_258 = img_reg_array_32_52_real;
        _zz_259 = img_reg_array_32_52_imag;
        _zz_260 = img_reg_array_33_52_real;
        _zz_261 = img_reg_array_33_52_imag;
        _zz_262 = img_reg_array_34_52_real;
        _zz_263 = img_reg_array_34_52_imag;
        _zz_264 = img_reg_array_35_52_real;
        _zz_265 = img_reg_array_35_52_imag;
        _zz_266 = img_reg_array_36_52_real;
        _zz_267 = img_reg_array_36_52_imag;
        _zz_268 = img_reg_array_37_52_real;
        _zz_269 = img_reg_array_37_52_imag;
        _zz_270 = img_reg_array_38_52_real;
        _zz_271 = img_reg_array_38_52_imag;
        _zz_272 = img_reg_array_39_52_real;
        _zz_273 = img_reg_array_39_52_imag;
        _zz_274 = img_reg_array_40_52_real;
        _zz_275 = img_reg_array_40_52_imag;
        _zz_276 = img_reg_array_41_52_real;
        _zz_277 = img_reg_array_41_52_imag;
        _zz_278 = img_reg_array_42_52_real;
        _zz_279 = img_reg_array_42_52_imag;
        _zz_280 = img_reg_array_43_52_real;
        _zz_281 = img_reg_array_43_52_imag;
        _zz_282 = img_reg_array_44_52_real;
        _zz_283 = img_reg_array_44_52_imag;
        _zz_284 = img_reg_array_45_52_real;
        _zz_285 = img_reg_array_45_52_imag;
        _zz_286 = img_reg_array_46_52_real;
        _zz_287 = img_reg_array_46_52_imag;
        _zz_288 = img_reg_array_47_52_real;
        _zz_289 = img_reg_array_47_52_imag;
        _zz_290 = img_reg_array_48_52_real;
        _zz_291 = img_reg_array_48_52_imag;
        _zz_292 = img_reg_array_49_52_real;
        _zz_293 = img_reg_array_49_52_imag;
        _zz_294 = img_reg_array_50_52_real;
        _zz_295 = img_reg_array_50_52_imag;
        _zz_296 = img_reg_array_51_52_real;
        _zz_297 = img_reg_array_51_52_imag;
        _zz_298 = img_reg_array_52_52_real;
        _zz_299 = img_reg_array_52_52_imag;
        _zz_300 = img_reg_array_53_52_real;
        _zz_301 = img_reg_array_53_52_imag;
        _zz_302 = img_reg_array_54_52_real;
        _zz_303 = img_reg_array_54_52_imag;
        _zz_304 = img_reg_array_55_52_real;
        _zz_305 = img_reg_array_55_52_imag;
        _zz_306 = img_reg_array_56_52_real;
        _zz_307 = img_reg_array_56_52_imag;
        _zz_308 = img_reg_array_57_52_real;
        _zz_309 = img_reg_array_57_52_imag;
        _zz_310 = img_reg_array_58_52_real;
        _zz_311 = img_reg_array_58_52_imag;
        _zz_312 = img_reg_array_59_52_real;
        _zz_313 = img_reg_array_59_52_imag;
        _zz_314 = img_reg_array_60_52_real;
        _zz_315 = img_reg_array_60_52_imag;
        _zz_316 = img_reg_array_61_52_real;
        _zz_317 = img_reg_array_61_52_imag;
        _zz_318 = img_reg_array_62_52_real;
        _zz_319 = img_reg_array_62_52_imag;
        _zz_320 = img_reg_array_63_52_real;
        _zz_321 = img_reg_array_63_52_imag;
      end
      6'b110101 : begin
        _zz_194 = img_reg_array_0_53_real;
        _zz_195 = img_reg_array_0_53_imag;
        _zz_196 = img_reg_array_1_53_real;
        _zz_197 = img_reg_array_1_53_imag;
        _zz_198 = img_reg_array_2_53_real;
        _zz_199 = img_reg_array_2_53_imag;
        _zz_200 = img_reg_array_3_53_real;
        _zz_201 = img_reg_array_3_53_imag;
        _zz_202 = img_reg_array_4_53_real;
        _zz_203 = img_reg_array_4_53_imag;
        _zz_204 = img_reg_array_5_53_real;
        _zz_205 = img_reg_array_5_53_imag;
        _zz_206 = img_reg_array_6_53_real;
        _zz_207 = img_reg_array_6_53_imag;
        _zz_208 = img_reg_array_7_53_real;
        _zz_209 = img_reg_array_7_53_imag;
        _zz_210 = img_reg_array_8_53_real;
        _zz_211 = img_reg_array_8_53_imag;
        _zz_212 = img_reg_array_9_53_real;
        _zz_213 = img_reg_array_9_53_imag;
        _zz_214 = img_reg_array_10_53_real;
        _zz_215 = img_reg_array_10_53_imag;
        _zz_216 = img_reg_array_11_53_real;
        _zz_217 = img_reg_array_11_53_imag;
        _zz_218 = img_reg_array_12_53_real;
        _zz_219 = img_reg_array_12_53_imag;
        _zz_220 = img_reg_array_13_53_real;
        _zz_221 = img_reg_array_13_53_imag;
        _zz_222 = img_reg_array_14_53_real;
        _zz_223 = img_reg_array_14_53_imag;
        _zz_224 = img_reg_array_15_53_real;
        _zz_225 = img_reg_array_15_53_imag;
        _zz_226 = img_reg_array_16_53_real;
        _zz_227 = img_reg_array_16_53_imag;
        _zz_228 = img_reg_array_17_53_real;
        _zz_229 = img_reg_array_17_53_imag;
        _zz_230 = img_reg_array_18_53_real;
        _zz_231 = img_reg_array_18_53_imag;
        _zz_232 = img_reg_array_19_53_real;
        _zz_233 = img_reg_array_19_53_imag;
        _zz_234 = img_reg_array_20_53_real;
        _zz_235 = img_reg_array_20_53_imag;
        _zz_236 = img_reg_array_21_53_real;
        _zz_237 = img_reg_array_21_53_imag;
        _zz_238 = img_reg_array_22_53_real;
        _zz_239 = img_reg_array_22_53_imag;
        _zz_240 = img_reg_array_23_53_real;
        _zz_241 = img_reg_array_23_53_imag;
        _zz_242 = img_reg_array_24_53_real;
        _zz_243 = img_reg_array_24_53_imag;
        _zz_244 = img_reg_array_25_53_real;
        _zz_245 = img_reg_array_25_53_imag;
        _zz_246 = img_reg_array_26_53_real;
        _zz_247 = img_reg_array_26_53_imag;
        _zz_248 = img_reg_array_27_53_real;
        _zz_249 = img_reg_array_27_53_imag;
        _zz_250 = img_reg_array_28_53_real;
        _zz_251 = img_reg_array_28_53_imag;
        _zz_252 = img_reg_array_29_53_real;
        _zz_253 = img_reg_array_29_53_imag;
        _zz_254 = img_reg_array_30_53_real;
        _zz_255 = img_reg_array_30_53_imag;
        _zz_256 = img_reg_array_31_53_real;
        _zz_257 = img_reg_array_31_53_imag;
        _zz_258 = img_reg_array_32_53_real;
        _zz_259 = img_reg_array_32_53_imag;
        _zz_260 = img_reg_array_33_53_real;
        _zz_261 = img_reg_array_33_53_imag;
        _zz_262 = img_reg_array_34_53_real;
        _zz_263 = img_reg_array_34_53_imag;
        _zz_264 = img_reg_array_35_53_real;
        _zz_265 = img_reg_array_35_53_imag;
        _zz_266 = img_reg_array_36_53_real;
        _zz_267 = img_reg_array_36_53_imag;
        _zz_268 = img_reg_array_37_53_real;
        _zz_269 = img_reg_array_37_53_imag;
        _zz_270 = img_reg_array_38_53_real;
        _zz_271 = img_reg_array_38_53_imag;
        _zz_272 = img_reg_array_39_53_real;
        _zz_273 = img_reg_array_39_53_imag;
        _zz_274 = img_reg_array_40_53_real;
        _zz_275 = img_reg_array_40_53_imag;
        _zz_276 = img_reg_array_41_53_real;
        _zz_277 = img_reg_array_41_53_imag;
        _zz_278 = img_reg_array_42_53_real;
        _zz_279 = img_reg_array_42_53_imag;
        _zz_280 = img_reg_array_43_53_real;
        _zz_281 = img_reg_array_43_53_imag;
        _zz_282 = img_reg_array_44_53_real;
        _zz_283 = img_reg_array_44_53_imag;
        _zz_284 = img_reg_array_45_53_real;
        _zz_285 = img_reg_array_45_53_imag;
        _zz_286 = img_reg_array_46_53_real;
        _zz_287 = img_reg_array_46_53_imag;
        _zz_288 = img_reg_array_47_53_real;
        _zz_289 = img_reg_array_47_53_imag;
        _zz_290 = img_reg_array_48_53_real;
        _zz_291 = img_reg_array_48_53_imag;
        _zz_292 = img_reg_array_49_53_real;
        _zz_293 = img_reg_array_49_53_imag;
        _zz_294 = img_reg_array_50_53_real;
        _zz_295 = img_reg_array_50_53_imag;
        _zz_296 = img_reg_array_51_53_real;
        _zz_297 = img_reg_array_51_53_imag;
        _zz_298 = img_reg_array_52_53_real;
        _zz_299 = img_reg_array_52_53_imag;
        _zz_300 = img_reg_array_53_53_real;
        _zz_301 = img_reg_array_53_53_imag;
        _zz_302 = img_reg_array_54_53_real;
        _zz_303 = img_reg_array_54_53_imag;
        _zz_304 = img_reg_array_55_53_real;
        _zz_305 = img_reg_array_55_53_imag;
        _zz_306 = img_reg_array_56_53_real;
        _zz_307 = img_reg_array_56_53_imag;
        _zz_308 = img_reg_array_57_53_real;
        _zz_309 = img_reg_array_57_53_imag;
        _zz_310 = img_reg_array_58_53_real;
        _zz_311 = img_reg_array_58_53_imag;
        _zz_312 = img_reg_array_59_53_real;
        _zz_313 = img_reg_array_59_53_imag;
        _zz_314 = img_reg_array_60_53_real;
        _zz_315 = img_reg_array_60_53_imag;
        _zz_316 = img_reg_array_61_53_real;
        _zz_317 = img_reg_array_61_53_imag;
        _zz_318 = img_reg_array_62_53_real;
        _zz_319 = img_reg_array_62_53_imag;
        _zz_320 = img_reg_array_63_53_real;
        _zz_321 = img_reg_array_63_53_imag;
      end
      6'b110110 : begin
        _zz_194 = img_reg_array_0_54_real;
        _zz_195 = img_reg_array_0_54_imag;
        _zz_196 = img_reg_array_1_54_real;
        _zz_197 = img_reg_array_1_54_imag;
        _zz_198 = img_reg_array_2_54_real;
        _zz_199 = img_reg_array_2_54_imag;
        _zz_200 = img_reg_array_3_54_real;
        _zz_201 = img_reg_array_3_54_imag;
        _zz_202 = img_reg_array_4_54_real;
        _zz_203 = img_reg_array_4_54_imag;
        _zz_204 = img_reg_array_5_54_real;
        _zz_205 = img_reg_array_5_54_imag;
        _zz_206 = img_reg_array_6_54_real;
        _zz_207 = img_reg_array_6_54_imag;
        _zz_208 = img_reg_array_7_54_real;
        _zz_209 = img_reg_array_7_54_imag;
        _zz_210 = img_reg_array_8_54_real;
        _zz_211 = img_reg_array_8_54_imag;
        _zz_212 = img_reg_array_9_54_real;
        _zz_213 = img_reg_array_9_54_imag;
        _zz_214 = img_reg_array_10_54_real;
        _zz_215 = img_reg_array_10_54_imag;
        _zz_216 = img_reg_array_11_54_real;
        _zz_217 = img_reg_array_11_54_imag;
        _zz_218 = img_reg_array_12_54_real;
        _zz_219 = img_reg_array_12_54_imag;
        _zz_220 = img_reg_array_13_54_real;
        _zz_221 = img_reg_array_13_54_imag;
        _zz_222 = img_reg_array_14_54_real;
        _zz_223 = img_reg_array_14_54_imag;
        _zz_224 = img_reg_array_15_54_real;
        _zz_225 = img_reg_array_15_54_imag;
        _zz_226 = img_reg_array_16_54_real;
        _zz_227 = img_reg_array_16_54_imag;
        _zz_228 = img_reg_array_17_54_real;
        _zz_229 = img_reg_array_17_54_imag;
        _zz_230 = img_reg_array_18_54_real;
        _zz_231 = img_reg_array_18_54_imag;
        _zz_232 = img_reg_array_19_54_real;
        _zz_233 = img_reg_array_19_54_imag;
        _zz_234 = img_reg_array_20_54_real;
        _zz_235 = img_reg_array_20_54_imag;
        _zz_236 = img_reg_array_21_54_real;
        _zz_237 = img_reg_array_21_54_imag;
        _zz_238 = img_reg_array_22_54_real;
        _zz_239 = img_reg_array_22_54_imag;
        _zz_240 = img_reg_array_23_54_real;
        _zz_241 = img_reg_array_23_54_imag;
        _zz_242 = img_reg_array_24_54_real;
        _zz_243 = img_reg_array_24_54_imag;
        _zz_244 = img_reg_array_25_54_real;
        _zz_245 = img_reg_array_25_54_imag;
        _zz_246 = img_reg_array_26_54_real;
        _zz_247 = img_reg_array_26_54_imag;
        _zz_248 = img_reg_array_27_54_real;
        _zz_249 = img_reg_array_27_54_imag;
        _zz_250 = img_reg_array_28_54_real;
        _zz_251 = img_reg_array_28_54_imag;
        _zz_252 = img_reg_array_29_54_real;
        _zz_253 = img_reg_array_29_54_imag;
        _zz_254 = img_reg_array_30_54_real;
        _zz_255 = img_reg_array_30_54_imag;
        _zz_256 = img_reg_array_31_54_real;
        _zz_257 = img_reg_array_31_54_imag;
        _zz_258 = img_reg_array_32_54_real;
        _zz_259 = img_reg_array_32_54_imag;
        _zz_260 = img_reg_array_33_54_real;
        _zz_261 = img_reg_array_33_54_imag;
        _zz_262 = img_reg_array_34_54_real;
        _zz_263 = img_reg_array_34_54_imag;
        _zz_264 = img_reg_array_35_54_real;
        _zz_265 = img_reg_array_35_54_imag;
        _zz_266 = img_reg_array_36_54_real;
        _zz_267 = img_reg_array_36_54_imag;
        _zz_268 = img_reg_array_37_54_real;
        _zz_269 = img_reg_array_37_54_imag;
        _zz_270 = img_reg_array_38_54_real;
        _zz_271 = img_reg_array_38_54_imag;
        _zz_272 = img_reg_array_39_54_real;
        _zz_273 = img_reg_array_39_54_imag;
        _zz_274 = img_reg_array_40_54_real;
        _zz_275 = img_reg_array_40_54_imag;
        _zz_276 = img_reg_array_41_54_real;
        _zz_277 = img_reg_array_41_54_imag;
        _zz_278 = img_reg_array_42_54_real;
        _zz_279 = img_reg_array_42_54_imag;
        _zz_280 = img_reg_array_43_54_real;
        _zz_281 = img_reg_array_43_54_imag;
        _zz_282 = img_reg_array_44_54_real;
        _zz_283 = img_reg_array_44_54_imag;
        _zz_284 = img_reg_array_45_54_real;
        _zz_285 = img_reg_array_45_54_imag;
        _zz_286 = img_reg_array_46_54_real;
        _zz_287 = img_reg_array_46_54_imag;
        _zz_288 = img_reg_array_47_54_real;
        _zz_289 = img_reg_array_47_54_imag;
        _zz_290 = img_reg_array_48_54_real;
        _zz_291 = img_reg_array_48_54_imag;
        _zz_292 = img_reg_array_49_54_real;
        _zz_293 = img_reg_array_49_54_imag;
        _zz_294 = img_reg_array_50_54_real;
        _zz_295 = img_reg_array_50_54_imag;
        _zz_296 = img_reg_array_51_54_real;
        _zz_297 = img_reg_array_51_54_imag;
        _zz_298 = img_reg_array_52_54_real;
        _zz_299 = img_reg_array_52_54_imag;
        _zz_300 = img_reg_array_53_54_real;
        _zz_301 = img_reg_array_53_54_imag;
        _zz_302 = img_reg_array_54_54_real;
        _zz_303 = img_reg_array_54_54_imag;
        _zz_304 = img_reg_array_55_54_real;
        _zz_305 = img_reg_array_55_54_imag;
        _zz_306 = img_reg_array_56_54_real;
        _zz_307 = img_reg_array_56_54_imag;
        _zz_308 = img_reg_array_57_54_real;
        _zz_309 = img_reg_array_57_54_imag;
        _zz_310 = img_reg_array_58_54_real;
        _zz_311 = img_reg_array_58_54_imag;
        _zz_312 = img_reg_array_59_54_real;
        _zz_313 = img_reg_array_59_54_imag;
        _zz_314 = img_reg_array_60_54_real;
        _zz_315 = img_reg_array_60_54_imag;
        _zz_316 = img_reg_array_61_54_real;
        _zz_317 = img_reg_array_61_54_imag;
        _zz_318 = img_reg_array_62_54_real;
        _zz_319 = img_reg_array_62_54_imag;
        _zz_320 = img_reg_array_63_54_real;
        _zz_321 = img_reg_array_63_54_imag;
      end
      6'b110111 : begin
        _zz_194 = img_reg_array_0_55_real;
        _zz_195 = img_reg_array_0_55_imag;
        _zz_196 = img_reg_array_1_55_real;
        _zz_197 = img_reg_array_1_55_imag;
        _zz_198 = img_reg_array_2_55_real;
        _zz_199 = img_reg_array_2_55_imag;
        _zz_200 = img_reg_array_3_55_real;
        _zz_201 = img_reg_array_3_55_imag;
        _zz_202 = img_reg_array_4_55_real;
        _zz_203 = img_reg_array_4_55_imag;
        _zz_204 = img_reg_array_5_55_real;
        _zz_205 = img_reg_array_5_55_imag;
        _zz_206 = img_reg_array_6_55_real;
        _zz_207 = img_reg_array_6_55_imag;
        _zz_208 = img_reg_array_7_55_real;
        _zz_209 = img_reg_array_7_55_imag;
        _zz_210 = img_reg_array_8_55_real;
        _zz_211 = img_reg_array_8_55_imag;
        _zz_212 = img_reg_array_9_55_real;
        _zz_213 = img_reg_array_9_55_imag;
        _zz_214 = img_reg_array_10_55_real;
        _zz_215 = img_reg_array_10_55_imag;
        _zz_216 = img_reg_array_11_55_real;
        _zz_217 = img_reg_array_11_55_imag;
        _zz_218 = img_reg_array_12_55_real;
        _zz_219 = img_reg_array_12_55_imag;
        _zz_220 = img_reg_array_13_55_real;
        _zz_221 = img_reg_array_13_55_imag;
        _zz_222 = img_reg_array_14_55_real;
        _zz_223 = img_reg_array_14_55_imag;
        _zz_224 = img_reg_array_15_55_real;
        _zz_225 = img_reg_array_15_55_imag;
        _zz_226 = img_reg_array_16_55_real;
        _zz_227 = img_reg_array_16_55_imag;
        _zz_228 = img_reg_array_17_55_real;
        _zz_229 = img_reg_array_17_55_imag;
        _zz_230 = img_reg_array_18_55_real;
        _zz_231 = img_reg_array_18_55_imag;
        _zz_232 = img_reg_array_19_55_real;
        _zz_233 = img_reg_array_19_55_imag;
        _zz_234 = img_reg_array_20_55_real;
        _zz_235 = img_reg_array_20_55_imag;
        _zz_236 = img_reg_array_21_55_real;
        _zz_237 = img_reg_array_21_55_imag;
        _zz_238 = img_reg_array_22_55_real;
        _zz_239 = img_reg_array_22_55_imag;
        _zz_240 = img_reg_array_23_55_real;
        _zz_241 = img_reg_array_23_55_imag;
        _zz_242 = img_reg_array_24_55_real;
        _zz_243 = img_reg_array_24_55_imag;
        _zz_244 = img_reg_array_25_55_real;
        _zz_245 = img_reg_array_25_55_imag;
        _zz_246 = img_reg_array_26_55_real;
        _zz_247 = img_reg_array_26_55_imag;
        _zz_248 = img_reg_array_27_55_real;
        _zz_249 = img_reg_array_27_55_imag;
        _zz_250 = img_reg_array_28_55_real;
        _zz_251 = img_reg_array_28_55_imag;
        _zz_252 = img_reg_array_29_55_real;
        _zz_253 = img_reg_array_29_55_imag;
        _zz_254 = img_reg_array_30_55_real;
        _zz_255 = img_reg_array_30_55_imag;
        _zz_256 = img_reg_array_31_55_real;
        _zz_257 = img_reg_array_31_55_imag;
        _zz_258 = img_reg_array_32_55_real;
        _zz_259 = img_reg_array_32_55_imag;
        _zz_260 = img_reg_array_33_55_real;
        _zz_261 = img_reg_array_33_55_imag;
        _zz_262 = img_reg_array_34_55_real;
        _zz_263 = img_reg_array_34_55_imag;
        _zz_264 = img_reg_array_35_55_real;
        _zz_265 = img_reg_array_35_55_imag;
        _zz_266 = img_reg_array_36_55_real;
        _zz_267 = img_reg_array_36_55_imag;
        _zz_268 = img_reg_array_37_55_real;
        _zz_269 = img_reg_array_37_55_imag;
        _zz_270 = img_reg_array_38_55_real;
        _zz_271 = img_reg_array_38_55_imag;
        _zz_272 = img_reg_array_39_55_real;
        _zz_273 = img_reg_array_39_55_imag;
        _zz_274 = img_reg_array_40_55_real;
        _zz_275 = img_reg_array_40_55_imag;
        _zz_276 = img_reg_array_41_55_real;
        _zz_277 = img_reg_array_41_55_imag;
        _zz_278 = img_reg_array_42_55_real;
        _zz_279 = img_reg_array_42_55_imag;
        _zz_280 = img_reg_array_43_55_real;
        _zz_281 = img_reg_array_43_55_imag;
        _zz_282 = img_reg_array_44_55_real;
        _zz_283 = img_reg_array_44_55_imag;
        _zz_284 = img_reg_array_45_55_real;
        _zz_285 = img_reg_array_45_55_imag;
        _zz_286 = img_reg_array_46_55_real;
        _zz_287 = img_reg_array_46_55_imag;
        _zz_288 = img_reg_array_47_55_real;
        _zz_289 = img_reg_array_47_55_imag;
        _zz_290 = img_reg_array_48_55_real;
        _zz_291 = img_reg_array_48_55_imag;
        _zz_292 = img_reg_array_49_55_real;
        _zz_293 = img_reg_array_49_55_imag;
        _zz_294 = img_reg_array_50_55_real;
        _zz_295 = img_reg_array_50_55_imag;
        _zz_296 = img_reg_array_51_55_real;
        _zz_297 = img_reg_array_51_55_imag;
        _zz_298 = img_reg_array_52_55_real;
        _zz_299 = img_reg_array_52_55_imag;
        _zz_300 = img_reg_array_53_55_real;
        _zz_301 = img_reg_array_53_55_imag;
        _zz_302 = img_reg_array_54_55_real;
        _zz_303 = img_reg_array_54_55_imag;
        _zz_304 = img_reg_array_55_55_real;
        _zz_305 = img_reg_array_55_55_imag;
        _zz_306 = img_reg_array_56_55_real;
        _zz_307 = img_reg_array_56_55_imag;
        _zz_308 = img_reg_array_57_55_real;
        _zz_309 = img_reg_array_57_55_imag;
        _zz_310 = img_reg_array_58_55_real;
        _zz_311 = img_reg_array_58_55_imag;
        _zz_312 = img_reg_array_59_55_real;
        _zz_313 = img_reg_array_59_55_imag;
        _zz_314 = img_reg_array_60_55_real;
        _zz_315 = img_reg_array_60_55_imag;
        _zz_316 = img_reg_array_61_55_real;
        _zz_317 = img_reg_array_61_55_imag;
        _zz_318 = img_reg_array_62_55_real;
        _zz_319 = img_reg_array_62_55_imag;
        _zz_320 = img_reg_array_63_55_real;
        _zz_321 = img_reg_array_63_55_imag;
      end
      6'b111000 : begin
        _zz_194 = img_reg_array_0_56_real;
        _zz_195 = img_reg_array_0_56_imag;
        _zz_196 = img_reg_array_1_56_real;
        _zz_197 = img_reg_array_1_56_imag;
        _zz_198 = img_reg_array_2_56_real;
        _zz_199 = img_reg_array_2_56_imag;
        _zz_200 = img_reg_array_3_56_real;
        _zz_201 = img_reg_array_3_56_imag;
        _zz_202 = img_reg_array_4_56_real;
        _zz_203 = img_reg_array_4_56_imag;
        _zz_204 = img_reg_array_5_56_real;
        _zz_205 = img_reg_array_5_56_imag;
        _zz_206 = img_reg_array_6_56_real;
        _zz_207 = img_reg_array_6_56_imag;
        _zz_208 = img_reg_array_7_56_real;
        _zz_209 = img_reg_array_7_56_imag;
        _zz_210 = img_reg_array_8_56_real;
        _zz_211 = img_reg_array_8_56_imag;
        _zz_212 = img_reg_array_9_56_real;
        _zz_213 = img_reg_array_9_56_imag;
        _zz_214 = img_reg_array_10_56_real;
        _zz_215 = img_reg_array_10_56_imag;
        _zz_216 = img_reg_array_11_56_real;
        _zz_217 = img_reg_array_11_56_imag;
        _zz_218 = img_reg_array_12_56_real;
        _zz_219 = img_reg_array_12_56_imag;
        _zz_220 = img_reg_array_13_56_real;
        _zz_221 = img_reg_array_13_56_imag;
        _zz_222 = img_reg_array_14_56_real;
        _zz_223 = img_reg_array_14_56_imag;
        _zz_224 = img_reg_array_15_56_real;
        _zz_225 = img_reg_array_15_56_imag;
        _zz_226 = img_reg_array_16_56_real;
        _zz_227 = img_reg_array_16_56_imag;
        _zz_228 = img_reg_array_17_56_real;
        _zz_229 = img_reg_array_17_56_imag;
        _zz_230 = img_reg_array_18_56_real;
        _zz_231 = img_reg_array_18_56_imag;
        _zz_232 = img_reg_array_19_56_real;
        _zz_233 = img_reg_array_19_56_imag;
        _zz_234 = img_reg_array_20_56_real;
        _zz_235 = img_reg_array_20_56_imag;
        _zz_236 = img_reg_array_21_56_real;
        _zz_237 = img_reg_array_21_56_imag;
        _zz_238 = img_reg_array_22_56_real;
        _zz_239 = img_reg_array_22_56_imag;
        _zz_240 = img_reg_array_23_56_real;
        _zz_241 = img_reg_array_23_56_imag;
        _zz_242 = img_reg_array_24_56_real;
        _zz_243 = img_reg_array_24_56_imag;
        _zz_244 = img_reg_array_25_56_real;
        _zz_245 = img_reg_array_25_56_imag;
        _zz_246 = img_reg_array_26_56_real;
        _zz_247 = img_reg_array_26_56_imag;
        _zz_248 = img_reg_array_27_56_real;
        _zz_249 = img_reg_array_27_56_imag;
        _zz_250 = img_reg_array_28_56_real;
        _zz_251 = img_reg_array_28_56_imag;
        _zz_252 = img_reg_array_29_56_real;
        _zz_253 = img_reg_array_29_56_imag;
        _zz_254 = img_reg_array_30_56_real;
        _zz_255 = img_reg_array_30_56_imag;
        _zz_256 = img_reg_array_31_56_real;
        _zz_257 = img_reg_array_31_56_imag;
        _zz_258 = img_reg_array_32_56_real;
        _zz_259 = img_reg_array_32_56_imag;
        _zz_260 = img_reg_array_33_56_real;
        _zz_261 = img_reg_array_33_56_imag;
        _zz_262 = img_reg_array_34_56_real;
        _zz_263 = img_reg_array_34_56_imag;
        _zz_264 = img_reg_array_35_56_real;
        _zz_265 = img_reg_array_35_56_imag;
        _zz_266 = img_reg_array_36_56_real;
        _zz_267 = img_reg_array_36_56_imag;
        _zz_268 = img_reg_array_37_56_real;
        _zz_269 = img_reg_array_37_56_imag;
        _zz_270 = img_reg_array_38_56_real;
        _zz_271 = img_reg_array_38_56_imag;
        _zz_272 = img_reg_array_39_56_real;
        _zz_273 = img_reg_array_39_56_imag;
        _zz_274 = img_reg_array_40_56_real;
        _zz_275 = img_reg_array_40_56_imag;
        _zz_276 = img_reg_array_41_56_real;
        _zz_277 = img_reg_array_41_56_imag;
        _zz_278 = img_reg_array_42_56_real;
        _zz_279 = img_reg_array_42_56_imag;
        _zz_280 = img_reg_array_43_56_real;
        _zz_281 = img_reg_array_43_56_imag;
        _zz_282 = img_reg_array_44_56_real;
        _zz_283 = img_reg_array_44_56_imag;
        _zz_284 = img_reg_array_45_56_real;
        _zz_285 = img_reg_array_45_56_imag;
        _zz_286 = img_reg_array_46_56_real;
        _zz_287 = img_reg_array_46_56_imag;
        _zz_288 = img_reg_array_47_56_real;
        _zz_289 = img_reg_array_47_56_imag;
        _zz_290 = img_reg_array_48_56_real;
        _zz_291 = img_reg_array_48_56_imag;
        _zz_292 = img_reg_array_49_56_real;
        _zz_293 = img_reg_array_49_56_imag;
        _zz_294 = img_reg_array_50_56_real;
        _zz_295 = img_reg_array_50_56_imag;
        _zz_296 = img_reg_array_51_56_real;
        _zz_297 = img_reg_array_51_56_imag;
        _zz_298 = img_reg_array_52_56_real;
        _zz_299 = img_reg_array_52_56_imag;
        _zz_300 = img_reg_array_53_56_real;
        _zz_301 = img_reg_array_53_56_imag;
        _zz_302 = img_reg_array_54_56_real;
        _zz_303 = img_reg_array_54_56_imag;
        _zz_304 = img_reg_array_55_56_real;
        _zz_305 = img_reg_array_55_56_imag;
        _zz_306 = img_reg_array_56_56_real;
        _zz_307 = img_reg_array_56_56_imag;
        _zz_308 = img_reg_array_57_56_real;
        _zz_309 = img_reg_array_57_56_imag;
        _zz_310 = img_reg_array_58_56_real;
        _zz_311 = img_reg_array_58_56_imag;
        _zz_312 = img_reg_array_59_56_real;
        _zz_313 = img_reg_array_59_56_imag;
        _zz_314 = img_reg_array_60_56_real;
        _zz_315 = img_reg_array_60_56_imag;
        _zz_316 = img_reg_array_61_56_real;
        _zz_317 = img_reg_array_61_56_imag;
        _zz_318 = img_reg_array_62_56_real;
        _zz_319 = img_reg_array_62_56_imag;
        _zz_320 = img_reg_array_63_56_real;
        _zz_321 = img_reg_array_63_56_imag;
      end
      6'b111001 : begin
        _zz_194 = img_reg_array_0_57_real;
        _zz_195 = img_reg_array_0_57_imag;
        _zz_196 = img_reg_array_1_57_real;
        _zz_197 = img_reg_array_1_57_imag;
        _zz_198 = img_reg_array_2_57_real;
        _zz_199 = img_reg_array_2_57_imag;
        _zz_200 = img_reg_array_3_57_real;
        _zz_201 = img_reg_array_3_57_imag;
        _zz_202 = img_reg_array_4_57_real;
        _zz_203 = img_reg_array_4_57_imag;
        _zz_204 = img_reg_array_5_57_real;
        _zz_205 = img_reg_array_5_57_imag;
        _zz_206 = img_reg_array_6_57_real;
        _zz_207 = img_reg_array_6_57_imag;
        _zz_208 = img_reg_array_7_57_real;
        _zz_209 = img_reg_array_7_57_imag;
        _zz_210 = img_reg_array_8_57_real;
        _zz_211 = img_reg_array_8_57_imag;
        _zz_212 = img_reg_array_9_57_real;
        _zz_213 = img_reg_array_9_57_imag;
        _zz_214 = img_reg_array_10_57_real;
        _zz_215 = img_reg_array_10_57_imag;
        _zz_216 = img_reg_array_11_57_real;
        _zz_217 = img_reg_array_11_57_imag;
        _zz_218 = img_reg_array_12_57_real;
        _zz_219 = img_reg_array_12_57_imag;
        _zz_220 = img_reg_array_13_57_real;
        _zz_221 = img_reg_array_13_57_imag;
        _zz_222 = img_reg_array_14_57_real;
        _zz_223 = img_reg_array_14_57_imag;
        _zz_224 = img_reg_array_15_57_real;
        _zz_225 = img_reg_array_15_57_imag;
        _zz_226 = img_reg_array_16_57_real;
        _zz_227 = img_reg_array_16_57_imag;
        _zz_228 = img_reg_array_17_57_real;
        _zz_229 = img_reg_array_17_57_imag;
        _zz_230 = img_reg_array_18_57_real;
        _zz_231 = img_reg_array_18_57_imag;
        _zz_232 = img_reg_array_19_57_real;
        _zz_233 = img_reg_array_19_57_imag;
        _zz_234 = img_reg_array_20_57_real;
        _zz_235 = img_reg_array_20_57_imag;
        _zz_236 = img_reg_array_21_57_real;
        _zz_237 = img_reg_array_21_57_imag;
        _zz_238 = img_reg_array_22_57_real;
        _zz_239 = img_reg_array_22_57_imag;
        _zz_240 = img_reg_array_23_57_real;
        _zz_241 = img_reg_array_23_57_imag;
        _zz_242 = img_reg_array_24_57_real;
        _zz_243 = img_reg_array_24_57_imag;
        _zz_244 = img_reg_array_25_57_real;
        _zz_245 = img_reg_array_25_57_imag;
        _zz_246 = img_reg_array_26_57_real;
        _zz_247 = img_reg_array_26_57_imag;
        _zz_248 = img_reg_array_27_57_real;
        _zz_249 = img_reg_array_27_57_imag;
        _zz_250 = img_reg_array_28_57_real;
        _zz_251 = img_reg_array_28_57_imag;
        _zz_252 = img_reg_array_29_57_real;
        _zz_253 = img_reg_array_29_57_imag;
        _zz_254 = img_reg_array_30_57_real;
        _zz_255 = img_reg_array_30_57_imag;
        _zz_256 = img_reg_array_31_57_real;
        _zz_257 = img_reg_array_31_57_imag;
        _zz_258 = img_reg_array_32_57_real;
        _zz_259 = img_reg_array_32_57_imag;
        _zz_260 = img_reg_array_33_57_real;
        _zz_261 = img_reg_array_33_57_imag;
        _zz_262 = img_reg_array_34_57_real;
        _zz_263 = img_reg_array_34_57_imag;
        _zz_264 = img_reg_array_35_57_real;
        _zz_265 = img_reg_array_35_57_imag;
        _zz_266 = img_reg_array_36_57_real;
        _zz_267 = img_reg_array_36_57_imag;
        _zz_268 = img_reg_array_37_57_real;
        _zz_269 = img_reg_array_37_57_imag;
        _zz_270 = img_reg_array_38_57_real;
        _zz_271 = img_reg_array_38_57_imag;
        _zz_272 = img_reg_array_39_57_real;
        _zz_273 = img_reg_array_39_57_imag;
        _zz_274 = img_reg_array_40_57_real;
        _zz_275 = img_reg_array_40_57_imag;
        _zz_276 = img_reg_array_41_57_real;
        _zz_277 = img_reg_array_41_57_imag;
        _zz_278 = img_reg_array_42_57_real;
        _zz_279 = img_reg_array_42_57_imag;
        _zz_280 = img_reg_array_43_57_real;
        _zz_281 = img_reg_array_43_57_imag;
        _zz_282 = img_reg_array_44_57_real;
        _zz_283 = img_reg_array_44_57_imag;
        _zz_284 = img_reg_array_45_57_real;
        _zz_285 = img_reg_array_45_57_imag;
        _zz_286 = img_reg_array_46_57_real;
        _zz_287 = img_reg_array_46_57_imag;
        _zz_288 = img_reg_array_47_57_real;
        _zz_289 = img_reg_array_47_57_imag;
        _zz_290 = img_reg_array_48_57_real;
        _zz_291 = img_reg_array_48_57_imag;
        _zz_292 = img_reg_array_49_57_real;
        _zz_293 = img_reg_array_49_57_imag;
        _zz_294 = img_reg_array_50_57_real;
        _zz_295 = img_reg_array_50_57_imag;
        _zz_296 = img_reg_array_51_57_real;
        _zz_297 = img_reg_array_51_57_imag;
        _zz_298 = img_reg_array_52_57_real;
        _zz_299 = img_reg_array_52_57_imag;
        _zz_300 = img_reg_array_53_57_real;
        _zz_301 = img_reg_array_53_57_imag;
        _zz_302 = img_reg_array_54_57_real;
        _zz_303 = img_reg_array_54_57_imag;
        _zz_304 = img_reg_array_55_57_real;
        _zz_305 = img_reg_array_55_57_imag;
        _zz_306 = img_reg_array_56_57_real;
        _zz_307 = img_reg_array_56_57_imag;
        _zz_308 = img_reg_array_57_57_real;
        _zz_309 = img_reg_array_57_57_imag;
        _zz_310 = img_reg_array_58_57_real;
        _zz_311 = img_reg_array_58_57_imag;
        _zz_312 = img_reg_array_59_57_real;
        _zz_313 = img_reg_array_59_57_imag;
        _zz_314 = img_reg_array_60_57_real;
        _zz_315 = img_reg_array_60_57_imag;
        _zz_316 = img_reg_array_61_57_real;
        _zz_317 = img_reg_array_61_57_imag;
        _zz_318 = img_reg_array_62_57_real;
        _zz_319 = img_reg_array_62_57_imag;
        _zz_320 = img_reg_array_63_57_real;
        _zz_321 = img_reg_array_63_57_imag;
      end
      6'b111010 : begin
        _zz_194 = img_reg_array_0_58_real;
        _zz_195 = img_reg_array_0_58_imag;
        _zz_196 = img_reg_array_1_58_real;
        _zz_197 = img_reg_array_1_58_imag;
        _zz_198 = img_reg_array_2_58_real;
        _zz_199 = img_reg_array_2_58_imag;
        _zz_200 = img_reg_array_3_58_real;
        _zz_201 = img_reg_array_3_58_imag;
        _zz_202 = img_reg_array_4_58_real;
        _zz_203 = img_reg_array_4_58_imag;
        _zz_204 = img_reg_array_5_58_real;
        _zz_205 = img_reg_array_5_58_imag;
        _zz_206 = img_reg_array_6_58_real;
        _zz_207 = img_reg_array_6_58_imag;
        _zz_208 = img_reg_array_7_58_real;
        _zz_209 = img_reg_array_7_58_imag;
        _zz_210 = img_reg_array_8_58_real;
        _zz_211 = img_reg_array_8_58_imag;
        _zz_212 = img_reg_array_9_58_real;
        _zz_213 = img_reg_array_9_58_imag;
        _zz_214 = img_reg_array_10_58_real;
        _zz_215 = img_reg_array_10_58_imag;
        _zz_216 = img_reg_array_11_58_real;
        _zz_217 = img_reg_array_11_58_imag;
        _zz_218 = img_reg_array_12_58_real;
        _zz_219 = img_reg_array_12_58_imag;
        _zz_220 = img_reg_array_13_58_real;
        _zz_221 = img_reg_array_13_58_imag;
        _zz_222 = img_reg_array_14_58_real;
        _zz_223 = img_reg_array_14_58_imag;
        _zz_224 = img_reg_array_15_58_real;
        _zz_225 = img_reg_array_15_58_imag;
        _zz_226 = img_reg_array_16_58_real;
        _zz_227 = img_reg_array_16_58_imag;
        _zz_228 = img_reg_array_17_58_real;
        _zz_229 = img_reg_array_17_58_imag;
        _zz_230 = img_reg_array_18_58_real;
        _zz_231 = img_reg_array_18_58_imag;
        _zz_232 = img_reg_array_19_58_real;
        _zz_233 = img_reg_array_19_58_imag;
        _zz_234 = img_reg_array_20_58_real;
        _zz_235 = img_reg_array_20_58_imag;
        _zz_236 = img_reg_array_21_58_real;
        _zz_237 = img_reg_array_21_58_imag;
        _zz_238 = img_reg_array_22_58_real;
        _zz_239 = img_reg_array_22_58_imag;
        _zz_240 = img_reg_array_23_58_real;
        _zz_241 = img_reg_array_23_58_imag;
        _zz_242 = img_reg_array_24_58_real;
        _zz_243 = img_reg_array_24_58_imag;
        _zz_244 = img_reg_array_25_58_real;
        _zz_245 = img_reg_array_25_58_imag;
        _zz_246 = img_reg_array_26_58_real;
        _zz_247 = img_reg_array_26_58_imag;
        _zz_248 = img_reg_array_27_58_real;
        _zz_249 = img_reg_array_27_58_imag;
        _zz_250 = img_reg_array_28_58_real;
        _zz_251 = img_reg_array_28_58_imag;
        _zz_252 = img_reg_array_29_58_real;
        _zz_253 = img_reg_array_29_58_imag;
        _zz_254 = img_reg_array_30_58_real;
        _zz_255 = img_reg_array_30_58_imag;
        _zz_256 = img_reg_array_31_58_real;
        _zz_257 = img_reg_array_31_58_imag;
        _zz_258 = img_reg_array_32_58_real;
        _zz_259 = img_reg_array_32_58_imag;
        _zz_260 = img_reg_array_33_58_real;
        _zz_261 = img_reg_array_33_58_imag;
        _zz_262 = img_reg_array_34_58_real;
        _zz_263 = img_reg_array_34_58_imag;
        _zz_264 = img_reg_array_35_58_real;
        _zz_265 = img_reg_array_35_58_imag;
        _zz_266 = img_reg_array_36_58_real;
        _zz_267 = img_reg_array_36_58_imag;
        _zz_268 = img_reg_array_37_58_real;
        _zz_269 = img_reg_array_37_58_imag;
        _zz_270 = img_reg_array_38_58_real;
        _zz_271 = img_reg_array_38_58_imag;
        _zz_272 = img_reg_array_39_58_real;
        _zz_273 = img_reg_array_39_58_imag;
        _zz_274 = img_reg_array_40_58_real;
        _zz_275 = img_reg_array_40_58_imag;
        _zz_276 = img_reg_array_41_58_real;
        _zz_277 = img_reg_array_41_58_imag;
        _zz_278 = img_reg_array_42_58_real;
        _zz_279 = img_reg_array_42_58_imag;
        _zz_280 = img_reg_array_43_58_real;
        _zz_281 = img_reg_array_43_58_imag;
        _zz_282 = img_reg_array_44_58_real;
        _zz_283 = img_reg_array_44_58_imag;
        _zz_284 = img_reg_array_45_58_real;
        _zz_285 = img_reg_array_45_58_imag;
        _zz_286 = img_reg_array_46_58_real;
        _zz_287 = img_reg_array_46_58_imag;
        _zz_288 = img_reg_array_47_58_real;
        _zz_289 = img_reg_array_47_58_imag;
        _zz_290 = img_reg_array_48_58_real;
        _zz_291 = img_reg_array_48_58_imag;
        _zz_292 = img_reg_array_49_58_real;
        _zz_293 = img_reg_array_49_58_imag;
        _zz_294 = img_reg_array_50_58_real;
        _zz_295 = img_reg_array_50_58_imag;
        _zz_296 = img_reg_array_51_58_real;
        _zz_297 = img_reg_array_51_58_imag;
        _zz_298 = img_reg_array_52_58_real;
        _zz_299 = img_reg_array_52_58_imag;
        _zz_300 = img_reg_array_53_58_real;
        _zz_301 = img_reg_array_53_58_imag;
        _zz_302 = img_reg_array_54_58_real;
        _zz_303 = img_reg_array_54_58_imag;
        _zz_304 = img_reg_array_55_58_real;
        _zz_305 = img_reg_array_55_58_imag;
        _zz_306 = img_reg_array_56_58_real;
        _zz_307 = img_reg_array_56_58_imag;
        _zz_308 = img_reg_array_57_58_real;
        _zz_309 = img_reg_array_57_58_imag;
        _zz_310 = img_reg_array_58_58_real;
        _zz_311 = img_reg_array_58_58_imag;
        _zz_312 = img_reg_array_59_58_real;
        _zz_313 = img_reg_array_59_58_imag;
        _zz_314 = img_reg_array_60_58_real;
        _zz_315 = img_reg_array_60_58_imag;
        _zz_316 = img_reg_array_61_58_real;
        _zz_317 = img_reg_array_61_58_imag;
        _zz_318 = img_reg_array_62_58_real;
        _zz_319 = img_reg_array_62_58_imag;
        _zz_320 = img_reg_array_63_58_real;
        _zz_321 = img_reg_array_63_58_imag;
      end
      6'b111011 : begin
        _zz_194 = img_reg_array_0_59_real;
        _zz_195 = img_reg_array_0_59_imag;
        _zz_196 = img_reg_array_1_59_real;
        _zz_197 = img_reg_array_1_59_imag;
        _zz_198 = img_reg_array_2_59_real;
        _zz_199 = img_reg_array_2_59_imag;
        _zz_200 = img_reg_array_3_59_real;
        _zz_201 = img_reg_array_3_59_imag;
        _zz_202 = img_reg_array_4_59_real;
        _zz_203 = img_reg_array_4_59_imag;
        _zz_204 = img_reg_array_5_59_real;
        _zz_205 = img_reg_array_5_59_imag;
        _zz_206 = img_reg_array_6_59_real;
        _zz_207 = img_reg_array_6_59_imag;
        _zz_208 = img_reg_array_7_59_real;
        _zz_209 = img_reg_array_7_59_imag;
        _zz_210 = img_reg_array_8_59_real;
        _zz_211 = img_reg_array_8_59_imag;
        _zz_212 = img_reg_array_9_59_real;
        _zz_213 = img_reg_array_9_59_imag;
        _zz_214 = img_reg_array_10_59_real;
        _zz_215 = img_reg_array_10_59_imag;
        _zz_216 = img_reg_array_11_59_real;
        _zz_217 = img_reg_array_11_59_imag;
        _zz_218 = img_reg_array_12_59_real;
        _zz_219 = img_reg_array_12_59_imag;
        _zz_220 = img_reg_array_13_59_real;
        _zz_221 = img_reg_array_13_59_imag;
        _zz_222 = img_reg_array_14_59_real;
        _zz_223 = img_reg_array_14_59_imag;
        _zz_224 = img_reg_array_15_59_real;
        _zz_225 = img_reg_array_15_59_imag;
        _zz_226 = img_reg_array_16_59_real;
        _zz_227 = img_reg_array_16_59_imag;
        _zz_228 = img_reg_array_17_59_real;
        _zz_229 = img_reg_array_17_59_imag;
        _zz_230 = img_reg_array_18_59_real;
        _zz_231 = img_reg_array_18_59_imag;
        _zz_232 = img_reg_array_19_59_real;
        _zz_233 = img_reg_array_19_59_imag;
        _zz_234 = img_reg_array_20_59_real;
        _zz_235 = img_reg_array_20_59_imag;
        _zz_236 = img_reg_array_21_59_real;
        _zz_237 = img_reg_array_21_59_imag;
        _zz_238 = img_reg_array_22_59_real;
        _zz_239 = img_reg_array_22_59_imag;
        _zz_240 = img_reg_array_23_59_real;
        _zz_241 = img_reg_array_23_59_imag;
        _zz_242 = img_reg_array_24_59_real;
        _zz_243 = img_reg_array_24_59_imag;
        _zz_244 = img_reg_array_25_59_real;
        _zz_245 = img_reg_array_25_59_imag;
        _zz_246 = img_reg_array_26_59_real;
        _zz_247 = img_reg_array_26_59_imag;
        _zz_248 = img_reg_array_27_59_real;
        _zz_249 = img_reg_array_27_59_imag;
        _zz_250 = img_reg_array_28_59_real;
        _zz_251 = img_reg_array_28_59_imag;
        _zz_252 = img_reg_array_29_59_real;
        _zz_253 = img_reg_array_29_59_imag;
        _zz_254 = img_reg_array_30_59_real;
        _zz_255 = img_reg_array_30_59_imag;
        _zz_256 = img_reg_array_31_59_real;
        _zz_257 = img_reg_array_31_59_imag;
        _zz_258 = img_reg_array_32_59_real;
        _zz_259 = img_reg_array_32_59_imag;
        _zz_260 = img_reg_array_33_59_real;
        _zz_261 = img_reg_array_33_59_imag;
        _zz_262 = img_reg_array_34_59_real;
        _zz_263 = img_reg_array_34_59_imag;
        _zz_264 = img_reg_array_35_59_real;
        _zz_265 = img_reg_array_35_59_imag;
        _zz_266 = img_reg_array_36_59_real;
        _zz_267 = img_reg_array_36_59_imag;
        _zz_268 = img_reg_array_37_59_real;
        _zz_269 = img_reg_array_37_59_imag;
        _zz_270 = img_reg_array_38_59_real;
        _zz_271 = img_reg_array_38_59_imag;
        _zz_272 = img_reg_array_39_59_real;
        _zz_273 = img_reg_array_39_59_imag;
        _zz_274 = img_reg_array_40_59_real;
        _zz_275 = img_reg_array_40_59_imag;
        _zz_276 = img_reg_array_41_59_real;
        _zz_277 = img_reg_array_41_59_imag;
        _zz_278 = img_reg_array_42_59_real;
        _zz_279 = img_reg_array_42_59_imag;
        _zz_280 = img_reg_array_43_59_real;
        _zz_281 = img_reg_array_43_59_imag;
        _zz_282 = img_reg_array_44_59_real;
        _zz_283 = img_reg_array_44_59_imag;
        _zz_284 = img_reg_array_45_59_real;
        _zz_285 = img_reg_array_45_59_imag;
        _zz_286 = img_reg_array_46_59_real;
        _zz_287 = img_reg_array_46_59_imag;
        _zz_288 = img_reg_array_47_59_real;
        _zz_289 = img_reg_array_47_59_imag;
        _zz_290 = img_reg_array_48_59_real;
        _zz_291 = img_reg_array_48_59_imag;
        _zz_292 = img_reg_array_49_59_real;
        _zz_293 = img_reg_array_49_59_imag;
        _zz_294 = img_reg_array_50_59_real;
        _zz_295 = img_reg_array_50_59_imag;
        _zz_296 = img_reg_array_51_59_real;
        _zz_297 = img_reg_array_51_59_imag;
        _zz_298 = img_reg_array_52_59_real;
        _zz_299 = img_reg_array_52_59_imag;
        _zz_300 = img_reg_array_53_59_real;
        _zz_301 = img_reg_array_53_59_imag;
        _zz_302 = img_reg_array_54_59_real;
        _zz_303 = img_reg_array_54_59_imag;
        _zz_304 = img_reg_array_55_59_real;
        _zz_305 = img_reg_array_55_59_imag;
        _zz_306 = img_reg_array_56_59_real;
        _zz_307 = img_reg_array_56_59_imag;
        _zz_308 = img_reg_array_57_59_real;
        _zz_309 = img_reg_array_57_59_imag;
        _zz_310 = img_reg_array_58_59_real;
        _zz_311 = img_reg_array_58_59_imag;
        _zz_312 = img_reg_array_59_59_real;
        _zz_313 = img_reg_array_59_59_imag;
        _zz_314 = img_reg_array_60_59_real;
        _zz_315 = img_reg_array_60_59_imag;
        _zz_316 = img_reg_array_61_59_real;
        _zz_317 = img_reg_array_61_59_imag;
        _zz_318 = img_reg_array_62_59_real;
        _zz_319 = img_reg_array_62_59_imag;
        _zz_320 = img_reg_array_63_59_real;
        _zz_321 = img_reg_array_63_59_imag;
      end
      6'b111100 : begin
        _zz_194 = img_reg_array_0_60_real;
        _zz_195 = img_reg_array_0_60_imag;
        _zz_196 = img_reg_array_1_60_real;
        _zz_197 = img_reg_array_1_60_imag;
        _zz_198 = img_reg_array_2_60_real;
        _zz_199 = img_reg_array_2_60_imag;
        _zz_200 = img_reg_array_3_60_real;
        _zz_201 = img_reg_array_3_60_imag;
        _zz_202 = img_reg_array_4_60_real;
        _zz_203 = img_reg_array_4_60_imag;
        _zz_204 = img_reg_array_5_60_real;
        _zz_205 = img_reg_array_5_60_imag;
        _zz_206 = img_reg_array_6_60_real;
        _zz_207 = img_reg_array_6_60_imag;
        _zz_208 = img_reg_array_7_60_real;
        _zz_209 = img_reg_array_7_60_imag;
        _zz_210 = img_reg_array_8_60_real;
        _zz_211 = img_reg_array_8_60_imag;
        _zz_212 = img_reg_array_9_60_real;
        _zz_213 = img_reg_array_9_60_imag;
        _zz_214 = img_reg_array_10_60_real;
        _zz_215 = img_reg_array_10_60_imag;
        _zz_216 = img_reg_array_11_60_real;
        _zz_217 = img_reg_array_11_60_imag;
        _zz_218 = img_reg_array_12_60_real;
        _zz_219 = img_reg_array_12_60_imag;
        _zz_220 = img_reg_array_13_60_real;
        _zz_221 = img_reg_array_13_60_imag;
        _zz_222 = img_reg_array_14_60_real;
        _zz_223 = img_reg_array_14_60_imag;
        _zz_224 = img_reg_array_15_60_real;
        _zz_225 = img_reg_array_15_60_imag;
        _zz_226 = img_reg_array_16_60_real;
        _zz_227 = img_reg_array_16_60_imag;
        _zz_228 = img_reg_array_17_60_real;
        _zz_229 = img_reg_array_17_60_imag;
        _zz_230 = img_reg_array_18_60_real;
        _zz_231 = img_reg_array_18_60_imag;
        _zz_232 = img_reg_array_19_60_real;
        _zz_233 = img_reg_array_19_60_imag;
        _zz_234 = img_reg_array_20_60_real;
        _zz_235 = img_reg_array_20_60_imag;
        _zz_236 = img_reg_array_21_60_real;
        _zz_237 = img_reg_array_21_60_imag;
        _zz_238 = img_reg_array_22_60_real;
        _zz_239 = img_reg_array_22_60_imag;
        _zz_240 = img_reg_array_23_60_real;
        _zz_241 = img_reg_array_23_60_imag;
        _zz_242 = img_reg_array_24_60_real;
        _zz_243 = img_reg_array_24_60_imag;
        _zz_244 = img_reg_array_25_60_real;
        _zz_245 = img_reg_array_25_60_imag;
        _zz_246 = img_reg_array_26_60_real;
        _zz_247 = img_reg_array_26_60_imag;
        _zz_248 = img_reg_array_27_60_real;
        _zz_249 = img_reg_array_27_60_imag;
        _zz_250 = img_reg_array_28_60_real;
        _zz_251 = img_reg_array_28_60_imag;
        _zz_252 = img_reg_array_29_60_real;
        _zz_253 = img_reg_array_29_60_imag;
        _zz_254 = img_reg_array_30_60_real;
        _zz_255 = img_reg_array_30_60_imag;
        _zz_256 = img_reg_array_31_60_real;
        _zz_257 = img_reg_array_31_60_imag;
        _zz_258 = img_reg_array_32_60_real;
        _zz_259 = img_reg_array_32_60_imag;
        _zz_260 = img_reg_array_33_60_real;
        _zz_261 = img_reg_array_33_60_imag;
        _zz_262 = img_reg_array_34_60_real;
        _zz_263 = img_reg_array_34_60_imag;
        _zz_264 = img_reg_array_35_60_real;
        _zz_265 = img_reg_array_35_60_imag;
        _zz_266 = img_reg_array_36_60_real;
        _zz_267 = img_reg_array_36_60_imag;
        _zz_268 = img_reg_array_37_60_real;
        _zz_269 = img_reg_array_37_60_imag;
        _zz_270 = img_reg_array_38_60_real;
        _zz_271 = img_reg_array_38_60_imag;
        _zz_272 = img_reg_array_39_60_real;
        _zz_273 = img_reg_array_39_60_imag;
        _zz_274 = img_reg_array_40_60_real;
        _zz_275 = img_reg_array_40_60_imag;
        _zz_276 = img_reg_array_41_60_real;
        _zz_277 = img_reg_array_41_60_imag;
        _zz_278 = img_reg_array_42_60_real;
        _zz_279 = img_reg_array_42_60_imag;
        _zz_280 = img_reg_array_43_60_real;
        _zz_281 = img_reg_array_43_60_imag;
        _zz_282 = img_reg_array_44_60_real;
        _zz_283 = img_reg_array_44_60_imag;
        _zz_284 = img_reg_array_45_60_real;
        _zz_285 = img_reg_array_45_60_imag;
        _zz_286 = img_reg_array_46_60_real;
        _zz_287 = img_reg_array_46_60_imag;
        _zz_288 = img_reg_array_47_60_real;
        _zz_289 = img_reg_array_47_60_imag;
        _zz_290 = img_reg_array_48_60_real;
        _zz_291 = img_reg_array_48_60_imag;
        _zz_292 = img_reg_array_49_60_real;
        _zz_293 = img_reg_array_49_60_imag;
        _zz_294 = img_reg_array_50_60_real;
        _zz_295 = img_reg_array_50_60_imag;
        _zz_296 = img_reg_array_51_60_real;
        _zz_297 = img_reg_array_51_60_imag;
        _zz_298 = img_reg_array_52_60_real;
        _zz_299 = img_reg_array_52_60_imag;
        _zz_300 = img_reg_array_53_60_real;
        _zz_301 = img_reg_array_53_60_imag;
        _zz_302 = img_reg_array_54_60_real;
        _zz_303 = img_reg_array_54_60_imag;
        _zz_304 = img_reg_array_55_60_real;
        _zz_305 = img_reg_array_55_60_imag;
        _zz_306 = img_reg_array_56_60_real;
        _zz_307 = img_reg_array_56_60_imag;
        _zz_308 = img_reg_array_57_60_real;
        _zz_309 = img_reg_array_57_60_imag;
        _zz_310 = img_reg_array_58_60_real;
        _zz_311 = img_reg_array_58_60_imag;
        _zz_312 = img_reg_array_59_60_real;
        _zz_313 = img_reg_array_59_60_imag;
        _zz_314 = img_reg_array_60_60_real;
        _zz_315 = img_reg_array_60_60_imag;
        _zz_316 = img_reg_array_61_60_real;
        _zz_317 = img_reg_array_61_60_imag;
        _zz_318 = img_reg_array_62_60_real;
        _zz_319 = img_reg_array_62_60_imag;
        _zz_320 = img_reg_array_63_60_real;
        _zz_321 = img_reg_array_63_60_imag;
      end
      6'b111101 : begin
        _zz_194 = img_reg_array_0_61_real;
        _zz_195 = img_reg_array_0_61_imag;
        _zz_196 = img_reg_array_1_61_real;
        _zz_197 = img_reg_array_1_61_imag;
        _zz_198 = img_reg_array_2_61_real;
        _zz_199 = img_reg_array_2_61_imag;
        _zz_200 = img_reg_array_3_61_real;
        _zz_201 = img_reg_array_3_61_imag;
        _zz_202 = img_reg_array_4_61_real;
        _zz_203 = img_reg_array_4_61_imag;
        _zz_204 = img_reg_array_5_61_real;
        _zz_205 = img_reg_array_5_61_imag;
        _zz_206 = img_reg_array_6_61_real;
        _zz_207 = img_reg_array_6_61_imag;
        _zz_208 = img_reg_array_7_61_real;
        _zz_209 = img_reg_array_7_61_imag;
        _zz_210 = img_reg_array_8_61_real;
        _zz_211 = img_reg_array_8_61_imag;
        _zz_212 = img_reg_array_9_61_real;
        _zz_213 = img_reg_array_9_61_imag;
        _zz_214 = img_reg_array_10_61_real;
        _zz_215 = img_reg_array_10_61_imag;
        _zz_216 = img_reg_array_11_61_real;
        _zz_217 = img_reg_array_11_61_imag;
        _zz_218 = img_reg_array_12_61_real;
        _zz_219 = img_reg_array_12_61_imag;
        _zz_220 = img_reg_array_13_61_real;
        _zz_221 = img_reg_array_13_61_imag;
        _zz_222 = img_reg_array_14_61_real;
        _zz_223 = img_reg_array_14_61_imag;
        _zz_224 = img_reg_array_15_61_real;
        _zz_225 = img_reg_array_15_61_imag;
        _zz_226 = img_reg_array_16_61_real;
        _zz_227 = img_reg_array_16_61_imag;
        _zz_228 = img_reg_array_17_61_real;
        _zz_229 = img_reg_array_17_61_imag;
        _zz_230 = img_reg_array_18_61_real;
        _zz_231 = img_reg_array_18_61_imag;
        _zz_232 = img_reg_array_19_61_real;
        _zz_233 = img_reg_array_19_61_imag;
        _zz_234 = img_reg_array_20_61_real;
        _zz_235 = img_reg_array_20_61_imag;
        _zz_236 = img_reg_array_21_61_real;
        _zz_237 = img_reg_array_21_61_imag;
        _zz_238 = img_reg_array_22_61_real;
        _zz_239 = img_reg_array_22_61_imag;
        _zz_240 = img_reg_array_23_61_real;
        _zz_241 = img_reg_array_23_61_imag;
        _zz_242 = img_reg_array_24_61_real;
        _zz_243 = img_reg_array_24_61_imag;
        _zz_244 = img_reg_array_25_61_real;
        _zz_245 = img_reg_array_25_61_imag;
        _zz_246 = img_reg_array_26_61_real;
        _zz_247 = img_reg_array_26_61_imag;
        _zz_248 = img_reg_array_27_61_real;
        _zz_249 = img_reg_array_27_61_imag;
        _zz_250 = img_reg_array_28_61_real;
        _zz_251 = img_reg_array_28_61_imag;
        _zz_252 = img_reg_array_29_61_real;
        _zz_253 = img_reg_array_29_61_imag;
        _zz_254 = img_reg_array_30_61_real;
        _zz_255 = img_reg_array_30_61_imag;
        _zz_256 = img_reg_array_31_61_real;
        _zz_257 = img_reg_array_31_61_imag;
        _zz_258 = img_reg_array_32_61_real;
        _zz_259 = img_reg_array_32_61_imag;
        _zz_260 = img_reg_array_33_61_real;
        _zz_261 = img_reg_array_33_61_imag;
        _zz_262 = img_reg_array_34_61_real;
        _zz_263 = img_reg_array_34_61_imag;
        _zz_264 = img_reg_array_35_61_real;
        _zz_265 = img_reg_array_35_61_imag;
        _zz_266 = img_reg_array_36_61_real;
        _zz_267 = img_reg_array_36_61_imag;
        _zz_268 = img_reg_array_37_61_real;
        _zz_269 = img_reg_array_37_61_imag;
        _zz_270 = img_reg_array_38_61_real;
        _zz_271 = img_reg_array_38_61_imag;
        _zz_272 = img_reg_array_39_61_real;
        _zz_273 = img_reg_array_39_61_imag;
        _zz_274 = img_reg_array_40_61_real;
        _zz_275 = img_reg_array_40_61_imag;
        _zz_276 = img_reg_array_41_61_real;
        _zz_277 = img_reg_array_41_61_imag;
        _zz_278 = img_reg_array_42_61_real;
        _zz_279 = img_reg_array_42_61_imag;
        _zz_280 = img_reg_array_43_61_real;
        _zz_281 = img_reg_array_43_61_imag;
        _zz_282 = img_reg_array_44_61_real;
        _zz_283 = img_reg_array_44_61_imag;
        _zz_284 = img_reg_array_45_61_real;
        _zz_285 = img_reg_array_45_61_imag;
        _zz_286 = img_reg_array_46_61_real;
        _zz_287 = img_reg_array_46_61_imag;
        _zz_288 = img_reg_array_47_61_real;
        _zz_289 = img_reg_array_47_61_imag;
        _zz_290 = img_reg_array_48_61_real;
        _zz_291 = img_reg_array_48_61_imag;
        _zz_292 = img_reg_array_49_61_real;
        _zz_293 = img_reg_array_49_61_imag;
        _zz_294 = img_reg_array_50_61_real;
        _zz_295 = img_reg_array_50_61_imag;
        _zz_296 = img_reg_array_51_61_real;
        _zz_297 = img_reg_array_51_61_imag;
        _zz_298 = img_reg_array_52_61_real;
        _zz_299 = img_reg_array_52_61_imag;
        _zz_300 = img_reg_array_53_61_real;
        _zz_301 = img_reg_array_53_61_imag;
        _zz_302 = img_reg_array_54_61_real;
        _zz_303 = img_reg_array_54_61_imag;
        _zz_304 = img_reg_array_55_61_real;
        _zz_305 = img_reg_array_55_61_imag;
        _zz_306 = img_reg_array_56_61_real;
        _zz_307 = img_reg_array_56_61_imag;
        _zz_308 = img_reg_array_57_61_real;
        _zz_309 = img_reg_array_57_61_imag;
        _zz_310 = img_reg_array_58_61_real;
        _zz_311 = img_reg_array_58_61_imag;
        _zz_312 = img_reg_array_59_61_real;
        _zz_313 = img_reg_array_59_61_imag;
        _zz_314 = img_reg_array_60_61_real;
        _zz_315 = img_reg_array_60_61_imag;
        _zz_316 = img_reg_array_61_61_real;
        _zz_317 = img_reg_array_61_61_imag;
        _zz_318 = img_reg_array_62_61_real;
        _zz_319 = img_reg_array_62_61_imag;
        _zz_320 = img_reg_array_63_61_real;
        _zz_321 = img_reg_array_63_61_imag;
      end
      6'b111110 : begin
        _zz_194 = img_reg_array_0_62_real;
        _zz_195 = img_reg_array_0_62_imag;
        _zz_196 = img_reg_array_1_62_real;
        _zz_197 = img_reg_array_1_62_imag;
        _zz_198 = img_reg_array_2_62_real;
        _zz_199 = img_reg_array_2_62_imag;
        _zz_200 = img_reg_array_3_62_real;
        _zz_201 = img_reg_array_3_62_imag;
        _zz_202 = img_reg_array_4_62_real;
        _zz_203 = img_reg_array_4_62_imag;
        _zz_204 = img_reg_array_5_62_real;
        _zz_205 = img_reg_array_5_62_imag;
        _zz_206 = img_reg_array_6_62_real;
        _zz_207 = img_reg_array_6_62_imag;
        _zz_208 = img_reg_array_7_62_real;
        _zz_209 = img_reg_array_7_62_imag;
        _zz_210 = img_reg_array_8_62_real;
        _zz_211 = img_reg_array_8_62_imag;
        _zz_212 = img_reg_array_9_62_real;
        _zz_213 = img_reg_array_9_62_imag;
        _zz_214 = img_reg_array_10_62_real;
        _zz_215 = img_reg_array_10_62_imag;
        _zz_216 = img_reg_array_11_62_real;
        _zz_217 = img_reg_array_11_62_imag;
        _zz_218 = img_reg_array_12_62_real;
        _zz_219 = img_reg_array_12_62_imag;
        _zz_220 = img_reg_array_13_62_real;
        _zz_221 = img_reg_array_13_62_imag;
        _zz_222 = img_reg_array_14_62_real;
        _zz_223 = img_reg_array_14_62_imag;
        _zz_224 = img_reg_array_15_62_real;
        _zz_225 = img_reg_array_15_62_imag;
        _zz_226 = img_reg_array_16_62_real;
        _zz_227 = img_reg_array_16_62_imag;
        _zz_228 = img_reg_array_17_62_real;
        _zz_229 = img_reg_array_17_62_imag;
        _zz_230 = img_reg_array_18_62_real;
        _zz_231 = img_reg_array_18_62_imag;
        _zz_232 = img_reg_array_19_62_real;
        _zz_233 = img_reg_array_19_62_imag;
        _zz_234 = img_reg_array_20_62_real;
        _zz_235 = img_reg_array_20_62_imag;
        _zz_236 = img_reg_array_21_62_real;
        _zz_237 = img_reg_array_21_62_imag;
        _zz_238 = img_reg_array_22_62_real;
        _zz_239 = img_reg_array_22_62_imag;
        _zz_240 = img_reg_array_23_62_real;
        _zz_241 = img_reg_array_23_62_imag;
        _zz_242 = img_reg_array_24_62_real;
        _zz_243 = img_reg_array_24_62_imag;
        _zz_244 = img_reg_array_25_62_real;
        _zz_245 = img_reg_array_25_62_imag;
        _zz_246 = img_reg_array_26_62_real;
        _zz_247 = img_reg_array_26_62_imag;
        _zz_248 = img_reg_array_27_62_real;
        _zz_249 = img_reg_array_27_62_imag;
        _zz_250 = img_reg_array_28_62_real;
        _zz_251 = img_reg_array_28_62_imag;
        _zz_252 = img_reg_array_29_62_real;
        _zz_253 = img_reg_array_29_62_imag;
        _zz_254 = img_reg_array_30_62_real;
        _zz_255 = img_reg_array_30_62_imag;
        _zz_256 = img_reg_array_31_62_real;
        _zz_257 = img_reg_array_31_62_imag;
        _zz_258 = img_reg_array_32_62_real;
        _zz_259 = img_reg_array_32_62_imag;
        _zz_260 = img_reg_array_33_62_real;
        _zz_261 = img_reg_array_33_62_imag;
        _zz_262 = img_reg_array_34_62_real;
        _zz_263 = img_reg_array_34_62_imag;
        _zz_264 = img_reg_array_35_62_real;
        _zz_265 = img_reg_array_35_62_imag;
        _zz_266 = img_reg_array_36_62_real;
        _zz_267 = img_reg_array_36_62_imag;
        _zz_268 = img_reg_array_37_62_real;
        _zz_269 = img_reg_array_37_62_imag;
        _zz_270 = img_reg_array_38_62_real;
        _zz_271 = img_reg_array_38_62_imag;
        _zz_272 = img_reg_array_39_62_real;
        _zz_273 = img_reg_array_39_62_imag;
        _zz_274 = img_reg_array_40_62_real;
        _zz_275 = img_reg_array_40_62_imag;
        _zz_276 = img_reg_array_41_62_real;
        _zz_277 = img_reg_array_41_62_imag;
        _zz_278 = img_reg_array_42_62_real;
        _zz_279 = img_reg_array_42_62_imag;
        _zz_280 = img_reg_array_43_62_real;
        _zz_281 = img_reg_array_43_62_imag;
        _zz_282 = img_reg_array_44_62_real;
        _zz_283 = img_reg_array_44_62_imag;
        _zz_284 = img_reg_array_45_62_real;
        _zz_285 = img_reg_array_45_62_imag;
        _zz_286 = img_reg_array_46_62_real;
        _zz_287 = img_reg_array_46_62_imag;
        _zz_288 = img_reg_array_47_62_real;
        _zz_289 = img_reg_array_47_62_imag;
        _zz_290 = img_reg_array_48_62_real;
        _zz_291 = img_reg_array_48_62_imag;
        _zz_292 = img_reg_array_49_62_real;
        _zz_293 = img_reg_array_49_62_imag;
        _zz_294 = img_reg_array_50_62_real;
        _zz_295 = img_reg_array_50_62_imag;
        _zz_296 = img_reg_array_51_62_real;
        _zz_297 = img_reg_array_51_62_imag;
        _zz_298 = img_reg_array_52_62_real;
        _zz_299 = img_reg_array_52_62_imag;
        _zz_300 = img_reg_array_53_62_real;
        _zz_301 = img_reg_array_53_62_imag;
        _zz_302 = img_reg_array_54_62_real;
        _zz_303 = img_reg_array_54_62_imag;
        _zz_304 = img_reg_array_55_62_real;
        _zz_305 = img_reg_array_55_62_imag;
        _zz_306 = img_reg_array_56_62_real;
        _zz_307 = img_reg_array_56_62_imag;
        _zz_308 = img_reg_array_57_62_real;
        _zz_309 = img_reg_array_57_62_imag;
        _zz_310 = img_reg_array_58_62_real;
        _zz_311 = img_reg_array_58_62_imag;
        _zz_312 = img_reg_array_59_62_real;
        _zz_313 = img_reg_array_59_62_imag;
        _zz_314 = img_reg_array_60_62_real;
        _zz_315 = img_reg_array_60_62_imag;
        _zz_316 = img_reg_array_61_62_real;
        _zz_317 = img_reg_array_61_62_imag;
        _zz_318 = img_reg_array_62_62_real;
        _zz_319 = img_reg_array_62_62_imag;
        _zz_320 = img_reg_array_63_62_real;
        _zz_321 = img_reg_array_63_62_imag;
      end
      default : begin
        _zz_194 = img_reg_array_0_63_real;
        _zz_195 = img_reg_array_0_63_imag;
        _zz_196 = img_reg_array_1_63_real;
        _zz_197 = img_reg_array_1_63_imag;
        _zz_198 = img_reg_array_2_63_real;
        _zz_199 = img_reg_array_2_63_imag;
        _zz_200 = img_reg_array_3_63_real;
        _zz_201 = img_reg_array_3_63_imag;
        _zz_202 = img_reg_array_4_63_real;
        _zz_203 = img_reg_array_4_63_imag;
        _zz_204 = img_reg_array_5_63_real;
        _zz_205 = img_reg_array_5_63_imag;
        _zz_206 = img_reg_array_6_63_real;
        _zz_207 = img_reg_array_6_63_imag;
        _zz_208 = img_reg_array_7_63_real;
        _zz_209 = img_reg_array_7_63_imag;
        _zz_210 = img_reg_array_8_63_real;
        _zz_211 = img_reg_array_8_63_imag;
        _zz_212 = img_reg_array_9_63_real;
        _zz_213 = img_reg_array_9_63_imag;
        _zz_214 = img_reg_array_10_63_real;
        _zz_215 = img_reg_array_10_63_imag;
        _zz_216 = img_reg_array_11_63_real;
        _zz_217 = img_reg_array_11_63_imag;
        _zz_218 = img_reg_array_12_63_real;
        _zz_219 = img_reg_array_12_63_imag;
        _zz_220 = img_reg_array_13_63_real;
        _zz_221 = img_reg_array_13_63_imag;
        _zz_222 = img_reg_array_14_63_real;
        _zz_223 = img_reg_array_14_63_imag;
        _zz_224 = img_reg_array_15_63_real;
        _zz_225 = img_reg_array_15_63_imag;
        _zz_226 = img_reg_array_16_63_real;
        _zz_227 = img_reg_array_16_63_imag;
        _zz_228 = img_reg_array_17_63_real;
        _zz_229 = img_reg_array_17_63_imag;
        _zz_230 = img_reg_array_18_63_real;
        _zz_231 = img_reg_array_18_63_imag;
        _zz_232 = img_reg_array_19_63_real;
        _zz_233 = img_reg_array_19_63_imag;
        _zz_234 = img_reg_array_20_63_real;
        _zz_235 = img_reg_array_20_63_imag;
        _zz_236 = img_reg_array_21_63_real;
        _zz_237 = img_reg_array_21_63_imag;
        _zz_238 = img_reg_array_22_63_real;
        _zz_239 = img_reg_array_22_63_imag;
        _zz_240 = img_reg_array_23_63_real;
        _zz_241 = img_reg_array_23_63_imag;
        _zz_242 = img_reg_array_24_63_real;
        _zz_243 = img_reg_array_24_63_imag;
        _zz_244 = img_reg_array_25_63_real;
        _zz_245 = img_reg_array_25_63_imag;
        _zz_246 = img_reg_array_26_63_real;
        _zz_247 = img_reg_array_26_63_imag;
        _zz_248 = img_reg_array_27_63_real;
        _zz_249 = img_reg_array_27_63_imag;
        _zz_250 = img_reg_array_28_63_real;
        _zz_251 = img_reg_array_28_63_imag;
        _zz_252 = img_reg_array_29_63_real;
        _zz_253 = img_reg_array_29_63_imag;
        _zz_254 = img_reg_array_30_63_real;
        _zz_255 = img_reg_array_30_63_imag;
        _zz_256 = img_reg_array_31_63_real;
        _zz_257 = img_reg_array_31_63_imag;
        _zz_258 = img_reg_array_32_63_real;
        _zz_259 = img_reg_array_32_63_imag;
        _zz_260 = img_reg_array_33_63_real;
        _zz_261 = img_reg_array_33_63_imag;
        _zz_262 = img_reg_array_34_63_real;
        _zz_263 = img_reg_array_34_63_imag;
        _zz_264 = img_reg_array_35_63_real;
        _zz_265 = img_reg_array_35_63_imag;
        _zz_266 = img_reg_array_36_63_real;
        _zz_267 = img_reg_array_36_63_imag;
        _zz_268 = img_reg_array_37_63_real;
        _zz_269 = img_reg_array_37_63_imag;
        _zz_270 = img_reg_array_38_63_real;
        _zz_271 = img_reg_array_38_63_imag;
        _zz_272 = img_reg_array_39_63_real;
        _zz_273 = img_reg_array_39_63_imag;
        _zz_274 = img_reg_array_40_63_real;
        _zz_275 = img_reg_array_40_63_imag;
        _zz_276 = img_reg_array_41_63_real;
        _zz_277 = img_reg_array_41_63_imag;
        _zz_278 = img_reg_array_42_63_real;
        _zz_279 = img_reg_array_42_63_imag;
        _zz_280 = img_reg_array_43_63_real;
        _zz_281 = img_reg_array_43_63_imag;
        _zz_282 = img_reg_array_44_63_real;
        _zz_283 = img_reg_array_44_63_imag;
        _zz_284 = img_reg_array_45_63_real;
        _zz_285 = img_reg_array_45_63_imag;
        _zz_286 = img_reg_array_46_63_real;
        _zz_287 = img_reg_array_46_63_imag;
        _zz_288 = img_reg_array_47_63_real;
        _zz_289 = img_reg_array_47_63_imag;
        _zz_290 = img_reg_array_48_63_real;
        _zz_291 = img_reg_array_48_63_imag;
        _zz_292 = img_reg_array_49_63_real;
        _zz_293 = img_reg_array_49_63_imag;
        _zz_294 = img_reg_array_50_63_real;
        _zz_295 = img_reg_array_50_63_imag;
        _zz_296 = img_reg_array_51_63_real;
        _zz_297 = img_reg_array_51_63_imag;
        _zz_298 = img_reg_array_52_63_real;
        _zz_299 = img_reg_array_52_63_imag;
        _zz_300 = img_reg_array_53_63_real;
        _zz_301 = img_reg_array_53_63_imag;
        _zz_302 = img_reg_array_54_63_real;
        _zz_303 = img_reg_array_54_63_imag;
        _zz_304 = img_reg_array_55_63_real;
        _zz_305 = img_reg_array_55_63_imag;
        _zz_306 = img_reg_array_56_63_real;
        _zz_307 = img_reg_array_56_63_imag;
        _zz_308 = img_reg_array_57_63_real;
        _zz_309 = img_reg_array_57_63_imag;
        _zz_310 = img_reg_array_58_63_real;
        _zz_311 = img_reg_array_58_63_imag;
        _zz_312 = img_reg_array_59_63_real;
        _zz_313 = img_reg_array_59_63_imag;
        _zz_314 = img_reg_array_60_63_real;
        _zz_315 = img_reg_array_60_63_imag;
        _zz_316 = img_reg_array_61_63_real;
        _zz_317 = img_reg_array_61_63_imag;
        _zz_318 = img_reg_array_62_63_real;
        _zz_319 = img_reg_array_62_63_imag;
        _zz_320 = img_reg_array_63_63_real;
        _zz_321 = img_reg_array_63_63_imag;
      end
    endcase
  end

  always @ (*) begin
    row_addr_willIncrement = 1'b0;
    if(myFFT_2_fft_row_valid)begin
      row_addr_willIncrement = 1'b1;
    end
  end

  assign row_addr_willClear = 1'b0;
  assign row_addr_willOverflowIfInc = (row_addr_value == 6'h3f);
  assign row_addr_willOverflow = (row_addr_willOverflowIfInc && row_addr_willIncrement);
  always @ (*) begin
    row_addr_valueNext = (row_addr_value + _zz_323);
    if(row_addr_willClear)begin
      row_addr_valueNext = 6'h0;
    end
  end

  assign _zz_1 = ({63'd0,1'b1} <<< row_addr_value);
  assign _zz_2 = _zz_1[0];
  assign _zz_3 = _zz_1[1];
  assign _zz_4 = _zz_1[2];
  assign _zz_5 = _zz_1[3];
  assign _zz_6 = _zz_1[4];
  assign _zz_7 = _zz_1[5];
  assign _zz_8 = _zz_1[6];
  assign _zz_9 = _zz_1[7];
  assign _zz_10 = _zz_1[8];
  assign _zz_11 = _zz_1[9];
  assign _zz_12 = _zz_1[10];
  assign _zz_13 = _zz_1[11];
  assign _zz_14 = _zz_1[12];
  assign _zz_15 = _zz_1[13];
  assign _zz_16 = _zz_1[14];
  assign _zz_17 = _zz_1[15];
  assign _zz_18 = _zz_1[16];
  assign _zz_19 = _zz_1[17];
  assign _zz_20 = _zz_1[18];
  assign _zz_21 = _zz_1[19];
  assign _zz_22 = _zz_1[20];
  assign _zz_23 = _zz_1[21];
  assign _zz_24 = _zz_1[22];
  assign _zz_25 = _zz_1[23];
  assign _zz_26 = _zz_1[24];
  assign _zz_27 = _zz_1[25];
  assign _zz_28 = _zz_1[26];
  assign _zz_29 = _zz_1[27];
  assign _zz_30 = _zz_1[28];
  assign _zz_31 = _zz_1[29];
  assign _zz_32 = _zz_1[30];
  assign _zz_33 = _zz_1[31];
  assign _zz_34 = _zz_1[32];
  assign _zz_35 = _zz_1[33];
  assign _zz_36 = _zz_1[34];
  assign _zz_37 = _zz_1[35];
  assign _zz_38 = _zz_1[36];
  assign _zz_39 = _zz_1[37];
  assign _zz_40 = _zz_1[38];
  assign _zz_41 = _zz_1[39];
  assign _zz_42 = _zz_1[40];
  assign _zz_43 = _zz_1[41];
  assign _zz_44 = _zz_1[42];
  assign _zz_45 = _zz_1[43];
  assign _zz_46 = _zz_1[44];
  assign _zz_47 = _zz_1[45];
  assign _zz_48 = _zz_1[46];
  assign _zz_49 = _zz_1[47];
  assign _zz_50 = _zz_1[48];
  assign _zz_51 = _zz_1[49];
  assign _zz_52 = _zz_1[50];
  assign _zz_53 = _zz_1[51];
  assign _zz_54 = _zz_1[52];
  assign _zz_55 = _zz_1[53];
  assign _zz_56 = _zz_1[54];
  assign _zz_57 = _zz_1[55];
  assign _zz_58 = _zz_1[56];
  assign _zz_59 = _zz_1[57];
  assign _zz_60 = _zz_1[58];
  assign _zz_61 = _zz_1[59];
  assign _zz_62 = _zz_1[60];
  assign _zz_63 = _zz_1[61];
  assign _zz_64 = _zz_1[62];
  assign _zz_65 = _zz_1[63];
  assign _zz_66 = myFFT_2_fft_row_payload_0_real;
  assign _zz_67 = myFFT_2_fft_row_payload_0_imag;
  assign _zz_68 = myFFT_2_fft_row_payload_1_real;
  assign _zz_69 = myFFT_2_fft_row_payload_1_imag;
  assign _zz_70 = myFFT_2_fft_row_payload_2_real;
  assign _zz_71 = myFFT_2_fft_row_payload_2_imag;
  assign _zz_72 = myFFT_2_fft_row_payload_3_real;
  assign _zz_73 = myFFT_2_fft_row_payload_3_imag;
  assign _zz_74 = myFFT_2_fft_row_payload_4_real;
  assign _zz_75 = myFFT_2_fft_row_payload_4_imag;
  assign _zz_76 = myFFT_2_fft_row_payload_5_real;
  assign _zz_77 = myFFT_2_fft_row_payload_5_imag;
  assign _zz_78 = myFFT_2_fft_row_payload_6_real;
  assign _zz_79 = myFFT_2_fft_row_payload_6_imag;
  assign _zz_80 = myFFT_2_fft_row_payload_7_real;
  assign _zz_81 = myFFT_2_fft_row_payload_7_imag;
  assign _zz_82 = myFFT_2_fft_row_payload_8_real;
  assign _zz_83 = myFFT_2_fft_row_payload_8_imag;
  assign _zz_84 = myFFT_2_fft_row_payload_9_real;
  assign _zz_85 = myFFT_2_fft_row_payload_9_imag;
  assign _zz_86 = myFFT_2_fft_row_payload_10_real;
  assign _zz_87 = myFFT_2_fft_row_payload_10_imag;
  assign _zz_88 = myFFT_2_fft_row_payload_11_real;
  assign _zz_89 = myFFT_2_fft_row_payload_11_imag;
  assign _zz_90 = myFFT_2_fft_row_payload_12_real;
  assign _zz_91 = myFFT_2_fft_row_payload_12_imag;
  assign _zz_92 = myFFT_2_fft_row_payload_13_real;
  assign _zz_93 = myFFT_2_fft_row_payload_13_imag;
  assign _zz_94 = myFFT_2_fft_row_payload_14_real;
  assign _zz_95 = myFFT_2_fft_row_payload_14_imag;
  assign _zz_96 = myFFT_2_fft_row_payload_15_real;
  assign _zz_97 = myFFT_2_fft_row_payload_15_imag;
  assign _zz_98 = myFFT_2_fft_row_payload_16_real;
  assign _zz_99 = myFFT_2_fft_row_payload_16_imag;
  assign _zz_100 = myFFT_2_fft_row_payload_17_real;
  assign _zz_101 = myFFT_2_fft_row_payload_17_imag;
  assign _zz_102 = myFFT_2_fft_row_payload_18_real;
  assign _zz_103 = myFFT_2_fft_row_payload_18_imag;
  assign _zz_104 = myFFT_2_fft_row_payload_19_real;
  assign _zz_105 = myFFT_2_fft_row_payload_19_imag;
  assign _zz_106 = myFFT_2_fft_row_payload_20_real;
  assign _zz_107 = myFFT_2_fft_row_payload_20_imag;
  assign _zz_108 = myFFT_2_fft_row_payload_21_real;
  assign _zz_109 = myFFT_2_fft_row_payload_21_imag;
  assign _zz_110 = myFFT_2_fft_row_payload_22_real;
  assign _zz_111 = myFFT_2_fft_row_payload_22_imag;
  assign _zz_112 = myFFT_2_fft_row_payload_23_real;
  assign _zz_113 = myFFT_2_fft_row_payload_23_imag;
  assign _zz_114 = myFFT_2_fft_row_payload_24_real;
  assign _zz_115 = myFFT_2_fft_row_payload_24_imag;
  assign _zz_116 = myFFT_2_fft_row_payload_25_real;
  assign _zz_117 = myFFT_2_fft_row_payload_25_imag;
  assign _zz_118 = myFFT_2_fft_row_payload_26_real;
  assign _zz_119 = myFFT_2_fft_row_payload_26_imag;
  assign _zz_120 = myFFT_2_fft_row_payload_27_real;
  assign _zz_121 = myFFT_2_fft_row_payload_27_imag;
  assign _zz_122 = myFFT_2_fft_row_payload_28_real;
  assign _zz_123 = myFFT_2_fft_row_payload_28_imag;
  assign _zz_124 = myFFT_2_fft_row_payload_29_real;
  assign _zz_125 = myFFT_2_fft_row_payload_29_imag;
  assign _zz_126 = myFFT_2_fft_row_payload_30_real;
  assign _zz_127 = myFFT_2_fft_row_payload_30_imag;
  assign _zz_128 = myFFT_2_fft_row_payload_31_real;
  assign _zz_129 = myFFT_2_fft_row_payload_31_imag;
  assign _zz_130 = myFFT_2_fft_row_payload_32_real;
  assign _zz_131 = myFFT_2_fft_row_payload_32_imag;
  assign _zz_132 = myFFT_2_fft_row_payload_33_real;
  assign _zz_133 = myFFT_2_fft_row_payload_33_imag;
  assign _zz_134 = myFFT_2_fft_row_payload_34_real;
  assign _zz_135 = myFFT_2_fft_row_payload_34_imag;
  assign _zz_136 = myFFT_2_fft_row_payload_35_real;
  assign _zz_137 = myFFT_2_fft_row_payload_35_imag;
  assign _zz_138 = myFFT_2_fft_row_payload_36_real;
  assign _zz_139 = myFFT_2_fft_row_payload_36_imag;
  assign _zz_140 = myFFT_2_fft_row_payload_37_real;
  assign _zz_141 = myFFT_2_fft_row_payload_37_imag;
  assign _zz_142 = myFFT_2_fft_row_payload_38_real;
  assign _zz_143 = myFFT_2_fft_row_payload_38_imag;
  assign _zz_144 = myFFT_2_fft_row_payload_39_real;
  assign _zz_145 = myFFT_2_fft_row_payload_39_imag;
  assign _zz_146 = myFFT_2_fft_row_payload_40_real;
  assign _zz_147 = myFFT_2_fft_row_payload_40_imag;
  assign _zz_148 = myFFT_2_fft_row_payload_41_real;
  assign _zz_149 = myFFT_2_fft_row_payload_41_imag;
  assign _zz_150 = myFFT_2_fft_row_payload_42_real;
  assign _zz_151 = myFFT_2_fft_row_payload_42_imag;
  assign _zz_152 = myFFT_2_fft_row_payload_43_real;
  assign _zz_153 = myFFT_2_fft_row_payload_43_imag;
  assign _zz_154 = myFFT_2_fft_row_payload_44_real;
  assign _zz_155 = myFFT_2_fft_row_payload_44_imag;
  assign _zz_156 = myFFT_2_fft_row_payload_45_real;
  assign _zz_157 = myFFT_2_fft_row_payload_45_imag;
  assign _zz_158 = myFFT_2_fft_row_payload_46_real;
  assign _zz_159 = myFFT_2_fft_row_payload_46_imag;
  assign _zz_160 = myFFT_2_fft_row_payload_47_real;
  assign _zz_161 = myFFT_2_fft_row_payload_47_imag;
  assign _zz_162 = myFFT_2_fft_row_payload_48_real;
  assign _zz_163 = myFFT_2_fft_row_payload_48_imag;
  assign _zz_164 = myFFT_2_fft_row_payload_49_real;
  assign _zz_165 = myFFT_2_fft_row_payload_49_imag;
  assign _zz_166 = myFFT_2_fft_row_payload_50_real;
  assign _zz_167 = myFFT_2_fft_row_payload_50_imag;
  assign _zz_168 = myFFT_2_fft_row_payload_51_real;
  assign _zz_169 = myFFT_2_fft_row_payload_51_imag;
  assign _zz_170 = myFFT_2_fft_row_payload_52_real;
  assign _zz_171 = myFFT_2_fft_row_payload_52_imag;
  assign _zz_172 = myFFT_2_fft_row_payload_53_real;
  assign _zz_173 = myFFT_2_fft_row_payload_53_imag;
  assign _zz_174 = myFFT_2_fft_row_payload_54_real;
  assign _zz_175 = myFFT_2_fft_row_payload_54_imag;
  assign _zz_176 = myFFT_2_fft_row_payload_55_real;
  assign _zz_177 = myFFT_2_fft_row_payload_55_imag;
  assign _zz_178 = myFFT_2_fft_row_payload_56_real;
  assign _zz_179 = myFFT_2_fft_row_payload_56_imag;
  assign _zz_180 = myFFT_2_fft_row_payload_57_real;
  assign _zz_181 = myFFT_2_fft_row_payload_57_imag;
  assign _zz_182 = myFFT_2_fft_row_payload_58_real;
  assign _zz_183 = myFFT_2_fft_row_payload_58_imag;
  assign _zz_184 = myFFT_2_fft_row_payload_59_real;
  assign _zz_185 = myFFT_2_fft_row_payload_59_imag;
  assign _zz_186 = myFFT_2_fft_row_payload_60_real;
  assign _zz_187 = myFFT_2_fft_row_payload_60_imag;
  assign _zz_188 = myFFT_2_fft_row_payload_61_real;
  assign _zz_189 = myFFT_2_fft_row_payload_61_imag;
  assign _zz_190 = myFFT_2_fft_row_payload_62_real;
  assign _zz_191 = myFFT_2_fft_row_payload_62_imag;
  assign _zz_192 = myFFT_2_fft_row_payload_63_real;
  assign _zz_193 = myFFT_2_fft_row_payload_63_imag;
  always @ (*) begin
    null_cnt_willIncrement = 1'b0;
    if(null_cond_period)begin
      null_cnt_willIncrement = 1'b1;
    end
  end

  assign null_cnt_willClear = 1'b0;
  assign null_cnt_willOverflowIfInc = (null_cnt_value == 6'h3f);
  assign null_cnt_willOverflow = (null_cnt_willOverflowIfInc && null_cnt_willIncrement);
  always @ (*) begin
    null_cnt_valueNext = (null_cnt_value + _zz_325);
    if(null_cnt_willClear)begin
      null_cnt_valueNext = 6'h0;
    end
  end

  assign null_cond_period = (row_addr_willOverflow || null_cond_period_minus_1);
  assign fft_col_in_payload_0_real = _zz_194;
  assign fft_col_in_payload_0_imag = _zz_195;
  assign fft_col_in_payload_1_real = _zz_196;
  assign fft_col_in_payload_1_imag = _zz_197;
  assign fft_col_in_payload_2_real = _zz_198;
  assign fft_col_in_payload_2_imag = _zz_199;
  assign fft_col_in_payload_3_real = _zz_200;
  assign fft_col_in_payload_3_imag = _zz_201;
  assign fft_col_in_payload_4_real = _zz_202;
  assign fft_col_in_payload_4_imag = _zz_203;
  assign fft_col_in_payload_5_real = _zz_204;
  assign fft_col_in_payload_5_imag = _zz_205;
  assign fft_col_in_payload_6_real = _zz_206;
  assign fft_col_in_payload_6_imag = _zz_207;
  assign fft_col_in_payload_7_real = _zz_208;
  assign fft_col_in_payload_7_imag = _zz_209;
  assign fft_col_in_payload_8_real = _zz_210;
  assign fft_col_in_payload_8_imag = _zz_211;
  assign fft_col_in_payload_9_real = _zz_212;
  assign fft_col_in_payload_9_imag = _zz_213;
  assign fft_col_in_payload_10_real = _zz_214;
  assign fft_col_in_payload_10_imag = _zz_215;
  assign fft_col_in_payload_11_real = _zz_216;
  assign fft_col_in_payload_11_imag = _zz_217;
  assign fft_col_in_payload_12_real = _zz_218;
  assign fft_col_in_payload_12_imag = _zz_219;
  assign fft_col_in_payload_13_real = _zz_220;
  assign fft_col_in_payload_13_imag = _zz_221;
  assign fft_col_in_payload_14_real = _zz_222;
  assign fft_col_in_payload_14_imag = _zz_223;
  assign fft_col_in_payload_15_real = _zz_224;
  assign fft_col_in_payload_15_imag = _zz_225;
  assign fft_col_in_payload_16_real = _zz_226;
  assign fft_col_in_payload_16_imag = _zz_227;
  assign fft_col_in_payload_17_real = _zz_228;
  assign fft_col_in_payload_17_imag = _zz_229;
  assign fft_col_in_payload_18_real = _zz_230;
  assign fft_col_in_payload_18_imag = _zz_231;
  assign fft_col_in_payload_19_real = _zz_232;
  assign fft_col_in_payload_19_imag = _zz_233;
  assign fft_col_in_payload_20_real = _zz_234;
  assign fft_col_in_payload_20_imag = _zz_235;
  assign fft_col_in_payload_21_real = _zz_236;
  assign fft_col_in_payload_21_imag = _zz_237;
  assign fft_col_in_payload_22_real = _zz_238;
  assign fft_col_in_payload_22_imag = _zz_239;
  assign fft_col_in_payload_23_real = _zz_240;
  assign fft_col_in_payload_23_imag = _zz_241;
  assign fft_col_in_payload_24_real = _zz_242;
  assign fft_col_in_payload_24_imag = _zz_243;
  assign fft_col_in_payload_25_real = _zz_244;
  assign fft_col_in_payload_25_imag = _zz_245;
  assign fft_col_in_payload_26_real = _zz_246;
  assign fft_col_in_payload_26_imag = _zz_247;
  assign fft_col_in_payload_27_real = _zz_248;
  assign fft_col_in_payload_27_imag = _zz_249;
  assign fft_col_in_payload_28_real = _zz_250;
  assign fft_col_in_payload_28_imag = _zz_251;
  assign fft_col_in_payload_29_real = _zz_252;
  assign fft_col_in_payload_29_imag = _zz_253;
  assign fft_col_in_payload_30_real = _zz_254;
  assign fft_col_in_payload_30_imag = _zz_255;
  assign fft_col_in_payload_31_real = _zz_256;
  assign fft_col_in_payload_31_imag = _zz_257;
  assign fft_col_in_payload_32_real = _zz_258;
  assign fft_col_in_payload_32_imag = _zz_259;
  assign fft_col_in_payload_33_real = _zz_260;
  assign fft_col_in_payload_33_imag = _zz_261;
  assign fft_col_in_payload_34_real = _zz_262;
  assign fft_col_in_payload_34_imag = _zz_263;
  assign fft_col_in_payload_35_real = _zz_264;
  assign fft_col_in_payload_35_imag = _zz_265;
  assign fft_col_in_payload_36_real = _zz_266;
  assign fft_col_in_payload_36_imag = _zz_267;
  assign fft_col_in_payload_37_real = _zz_268;
  assign fft_col_in_payload_37_imag = _zz_269;
  assign fft_col_in_payload_38_real = _zz_270;
  assign fft_col_in_payload_38_imag = _zz_271;
  assign fft_col_in_payload_39_real = _zz_272;
  assign fft_col_in_payload_39_imag = _zz_273;
  assign fft_col_in_payload_40_real = _zz_274;
  assign fft_col_in_payload_40_imag = _zz_275;
  assign fft_col_in_payload_41_real = _zz_276;
  assign fft_col_in_payload_41_imag = _zz_277;
  assign fft_col_in_payload_42_real = _zz_278;
  assign fft_col_in_payload_42_imag = _zz_279;
  assign fft_col_in_payload_43_real = _zz_280;
  assign fft_col_in_payload_43_imag = _zz_281;
  assign fft_col_in_payload_44_real = _zz_282;
  assign fft_col_in_payload_44_imag = _zz_283;
  assign fft_col_in_payload_45_real = _zz_284;
  assign fft_col_in_payload_45_imag = _zz_285;
  assign fft_col_in_payload_46_real = _zz_286;
  assign fft_col_in_payload_46_imag = _zz_287;
  assign fft_col_in_payload_47_real = _zz_288;
  assign fft_col_in_payload_47_imag = _zz_289;
  assign fft_col_in_payload_48_real = _zz_290;
  assign fft_col_in_payload_48_imag = _zz_291;
  assign fft_col_in_payload_49_real = _zz_292;
  assign fft_col_in_payload_49_imag = _zz_293;
  assign fft_col_in_payload_50_real = _zz_294;
  assign fft_col_in_payload_50_imag = _zz_295;
  assign fft_col_in_payload_51_real = _zz_296;
  assign fft_col_in_payload_51_imag = _zz_297;
  assign fft_col_in_payload_52_real = _zz_298;
  assign fft_col_in_payload_52_imag = _zz_299;
  assign fft_col_in_payload_53_real = _zz_300;
  assign fft_col_in_payload_53_imag = _zz_301;
  assign fft_col_in_payload_54_real = _zz_302;
  assign fft_col_in_payload_54_imag = _zz_303;
  assign fft_col_in_payload_55_real = _zz_304;
  assign fft_col_in_payload_55_imag = _zz_305;
  assign fft_col_in_payload_56_real = _zz_306;
  assign fft_col_in_payload_56_imag = _zz_307;
  assign fft_col_in_payload_57_real = _zz_308;
  assign fft_col_in_payload_57_imag = _zz_309;
  assign fft_col_in_payload_58_real = _zz_310;
  assign fft_col_in_payload_58_imag = _zz_311;
  assign fft_col_in_payload_59_real = _zz_312;
  assign fft_col_in_payload_59_imag = _zz_313;
  assign fft_col_in_payload_60_real = _zz_314;
  assign fft_col_in_payload_60_imag = _zz_315;
  assign fft_col_in_payload_61_real = _zz_316;
  assign fft_col_in_payload_61_imag = _zz_317;
  assign fft_col_in_payload_62_real = _zz_318;
  assign fft_col_in_payload_62_imag = _zz_319;
  assign fft_col_in_payload_63_real = _zz_320;
  assign fft_col_in_payload_63_imag = _zz_321;
  assign fft_col_in_valid = null_cond_period_regNext;
  assign io_line_out_valid = myFFT_3_fft_col_out_regNext_valid;
  assign io_line_out_payload_0_real = myFFT_3_fft_col_out_regNext_payload_0_real;
  assign io_line_out_payload_0_imag = myFFT_3_fft_col_out_regNext_payload_0_imag;
  assign io_line_out_payload_1_real = myFFT_3_fft_col_out_regNext_payload_1_real;
  assign io_line_out_payload_1_imag = myFFT_3_fft_col_out_regNext_payload_1_imag;
  assign io_line_out_payload_2_real = myFFT_3_fft_col_out_regNext_payload_2_real;
  assign io_line_out_payload_2_imag = myFFT_3_fft_col_out_regNext_payload_2_imag;
  assign io_line_out_payload_3_real = myFFT_3_fft_col_out_regNext_payload_3_real;
  assign io_line_out_payload_3_imag = myFFT_3_fft_col_out_regNext_payload_3_imag;
  assign io_line_out_payload_4_real = myFFT_3_fft_col_out_regNext_payload_4_real;
  assign io_line_out_payload_4_imag = myFFT_3_fft_col_out_regNext_payload_4_imag;
  assign io_line_out_payload_5_real = myFFT_3_fft_col_out_regNext_payload_5_real;
  assign io_line_out_payload_5_imag = myFFT_3_fft_col_out_regNext_payload_5_imag;
  assign io_line_out_payload_6_real = myFFT_3_fft_col_out_regNext_payload_6_real;
  assign io_line_out_payload_6_imag = myFFT_3_fft_col_out_regNext_payload_6_imag;
  assign io_line_out_payload_7_real = myFFT_3_fft_col_out_regNext_payload_7_real;
  assign io_line_out_payload_7_imag = myFFT_3_fft_col_out_regNext_payload_7_imag;
  assign io_line_out_payload_8_real = myFFT_3_fft_col_out_regNext_payload_8_real;
  assign io_line_out_payload_8_imag = myFFT_3_fft_col_out_regNext_payload_8_imag;
  assign io_line_out_payload_9_real = myFFT_3_fft_col_out_regNext_payload_9_real;
  assign io_line_out_payload_9_imag = myFFT_3_fft_col_out_regNext_payload_9_imag;
  assign io_line_out_payload_10_real = myFFT_3_fft_col_out_regNext_payload_10_real;
  assign io_line_out_payload_10_imag = myFFT_3_fft_col_out_regNext_payload_10_imag;
  assign io_line_out_payload_11_real = myFFT_3_fft_col_out_regNext_payload_11_real;
  assign io_line_out_payload_11_imag = myFFT_3_fft_col_out_regNext_payload_11_imag;
  assign io_line_out_payload_12_real = myFFT_3_fft_col_out_regNext_payload_12_real;
  assign io_line_out_payload_12_imag = myFFT_3_fft_col_out_regNext_payload_12_imag;
  assign io_line_out_payload_13_real = myFFT_3_fft_col_out_regNext_payload_13_real;
  assign io_line_out_payload_13_imag = myFFT_3_fft_col_out_regNext_payload_13_imag;
  assign io_line_out_payload_14_real = myFFT_3_fft_col_out_regNext_payload_14_real;
  assign io_line_out_payload_14_imag = myFFT_3_fft_col_out_regNext_payload_14_imag;
  assign io_line_out_payload_15_real = myFFT_3_fft_col_out_regNext_payload_15_real;
  assign io_line_out_payload_15_imag = myFFT_3_fft_col_out_regNext_payload_15_imag;
  assign io_line_out_payload_16_real = myFFT_3_fft_col_out_regNext_payload_16_real;
  assign io_line_out_payload_16_imag = myFFT_3_fft_col_out_regNext_payload_16_imag;
  assign io_line_out_payload_17_real = myFFT_3_fft_col_out_regNext_payload_17_real;
  assign io_line_out_payload_17_imag = myFFT_3_fft_col_out_regNext_payload_17_imag;
  assign io_line_out_payload_18_real = myFFT_3_fft_col_out_regNext_payload_18_real;
  assign io_line_out_payload_18_imag = myFFT_3_fft_col_out_regNext_payload_18_imag;
  assign io_line_out_payload_19_real = myFFT_3_fft_col_out_regNext_payload_19_real;
  assign io_line_out_payload_19_imag = myFFT_3_fft_col_out_regNext_payload_19_imag;
  assign io_line_out_payload_20_real = myFFT_3_fft_col_out_regNext_payload_20_real;
  assign io_line_out_payload_20_imag = myFFT_3_fft_col_out_regNext_payload_20_imag;
  assign io_line_out_payload_21_real = myFFT_3_fft_col_out_regNext_payload_21_real;
  assign io_line_out_payload_21_imag = myFFT_3_fft_col_out_regNext_payload_21_imag;
  assign io_line_out_payload_22_real = myFFT_3_fft_col_out_regNext_payload_22_real;
  assign io_line_out_payload_22_imag = myFFT_3_fft_col_out_regNext_payload_22_imag;
  assign io_line_out_payload_23_real = myFFT_3_fft_col_out_regNext_payload_23_real;
  assign io_line_out_payload_23_imag = myFFT_3_fft_col_out_regNext_payload_23_imag;
  assign io_line_out_payload_24_real = myFFT_3_fft_col_out_regNext_payload_24_real;
  assign io_line_out_payload_24_imag = myFFT_3_fft_col_out_regNext_payload_24_imag;
  assign io_line_out_payload_25_real = myFFT_3_fft_col_out_regNext_payload_25_real;
  assign io_line_out_payload_25_imag = myFFT_3_fft_col_out_regNext_payload_25_imag;
  assign io_line_out_payload_26_real = myFFT_3_fft_col_out_regNext_payload_26_real;
  assign io_line_out_payload_26_imag = myFFT_3_fft_col_out_regNext_payload_26_imag;
  assign io_line_out_payload_27_real = myFFT_3_fft_col_out_regNext_payload_27_real;
  assign io_line_out_payload_27_imag = myFFT_3_fft_col_out_regNext_payload_27_imag;
  assign io_line_out_payload_28_real = myFFT_3_fft_col_out_regNext_payload_28_real;
  assign io_line_out_payload_28_imag = myFFT_3_fft_col_out_regNext_payload_28_imag;
  assign io_line_out_payload_29_real = myFFT_3_fft_col_out_regNext_payload_29_real;
  assign io_line_out_payload_29_imag = myFFT_3_fft_col_out_regNext_payload_29_imag;
  assign io_line_out_payload_30_real = myFFT_3_fft_col_out_regNext_payload_30_real;
  assign io_line_out_payload_30_imag = myFFT_3_fft_col_out_regNext_payload_30_imag;
  assign io_line_out_payload_31_real = myFFT_3_fft_col_out_regNext_payload_31_real;
  assign io_line_out_payload_31_imag = myFFT_3_fft_col_out_regNext_payload_31_imag;
  assign io_line_out_payload_32_real = myFFT_3_fft_col_out_regNext_payload_32_real;
  assign io_line_out_payload_32_imag = myFFT_3_fft_col_out_regNext_payload_32_imag;
  assign io_line_out_payload_33_real = myFFT_3_fft_col_out_regNext_payload_33_real;
  assign io_line_out_payload_33_imag = myFFT_3_fft_col_out_regNext_payload_33_imag;
  assign io_line_out_payload_34_real = myFFT_3_fft_col_out_regNext_payload_34_real;
  assign io_line_out_payload_34_imag = myFFT_3_fft_col_out_regNext_payload_34_imag;
  assign io_line_out_payload_35_real = myFFT_3_fft_col_out_regNext_payload_35_real;
  assign io_line_out_payload_35_imag = myFFT_3_fft_col_out_regNext_payload_35_imag;
  assign io_line_out_payload_36_real = myFFT_3_fft_col_out_regNext_payload_36_real;
  assign io_line_out_payload_36_imag = myFFT_3_fft_col_out_regNext_payload_36_imag;
  assign io_line_out_payload_37_real = myFFT_3_fft_col_out_regNext_payload_37_real;
  assign io_line_out_payload_37_imag = myFFT_3_fft_col_out_regNext_payload_37_imag;
  assign io_line_out_payload_38_real = myFFT_3_fft_col_out_regNext_payload_38_real;
  assign io_line_out_payload_38_imag = myFFT_3_fft_col_out_regNext_payload_38_imag;
  assign io_line_out_payload_39_real = myFFT_3_fft_col_out_regNext_payload_39_real;
  assign io_line_out_payload_39_imag = myFFT_3_fft_col_out_regNext_payload_39_imag;
  assign io_line_out_payload_40_real = myFFT_3_fft_col_out_regNext_payload_40_real;
  assign io_line_out_payload_40_imag = myFFT_3_fft_col_out_regNext_payload_40_imag;
  assign io_line_out_payload_41_real = myFFT_3_fft_col_out_regNext_payload_41_real;
  assign io_line_out_payload_41_imag = myFFT_3_fft_col_out_regNext_payload_41_imag;
  assign io_line_out_payload_42_real = myFFT_3_fft_col_out_regNext_payload_42_real;
  assign io_line_out_payload_42_imag = myFFT_3_fft_col_out_regNext_payload_42_imag;
  assign io_line_out_payload_43_real = myFFT_3_fft_col_out_regNext_payload_43_real;
  assign io_line_out_payload_43_imag = myFFT_3_fft_col_out_regNext_payload_43_imag;
  assign io_line_out_payload_44_real = myFFT_3_fft_col_out_regNext_payload_44_real;
  assign io_line_out_payload_44_imag = myFFT_3_fft_col_out_regNext_payload_44_imag;
  assign io_line_out_payload_45_real = myFFT_3_fft_col_out_regNext_payload_45_real;
  assign io_line_out_payload_45_imag = myFFT_3_fft_col_out_regNext_payload_45_imag;
  assign io_line_out_payload_46_real = myFFT_3_fft_col_out_regNext_payload_46_real;
  assign io_line_out_payload_46_imag = myFFT_3_fft_col_out_regNext_payload_46_imag;
  assign io_line_out_payload_47_real = myFFT_3_fft_col_out_regNext_payload_47_real;
  assign io_line_out_payload_47_imag = myFFT_3_fft_col_out_regNext_payload_47_imag;
  assign io_line_out_payload_48_real = myFFT_3_fft_col_out_regNext_payload_48_real;
  assign io_line_out_payload_48_imag = myFFT_3_fft_col_out_regNext_payload_48_imag;
  assign io_line_out_payload_49_real = myFFT_3_fft_col_out_regNext_payload_49_real;
  assign io_line_out_payload_49_imag = myFFT_3_fft_col_out_regNext_payload_49_imag;
  assign io_line_out_payload_50_real = myFFT_3_fft_col_out_regNext_payload_50_real;
  assign io_line_out_payload_50_imag = myFFT_3_fft_col_out_regNext_payload_50_imag;
  assign io_line_out_payload_51_real = myFFT_3_fft_col_out_regNext_payload_51_real;
  assign io_line_out_payload_51_imag = myFFT_3_fft_col_out_regNext_payload_51_imag;
  assign io_line_out_payload_52_real = myFFT_3_fft_col_out_regNext_payload_52_real;
  assign io_line_out_payload_52_imag = myFFT_3_fft_col_out_regNext_payload_52_imag;
  assign io_line_out_payload_53_real = myFFT_3_fft_col_out_regNext_payload_53_real;
  assign io_line_out_payload_53_imag = myFFT_3_fft_col_out_regNext_payload_53_imag;
  assign io_line_out_payload_54_real = myFFT_3_fft_col_out_regNext_payload_54_real;
  assign io_line_out_payload_54_imag = myFFT_3_fft_col_out_regNext_payload_54_imag;
  assign io_line_out_payload_55_real = myFFT_3_fft_col_out_regNext_payload_55_real;
  assign io_line_out_payload_55_imag = myFFT_3_fft_col_out_regNext_payload_55_imag;
  assign io_line_out_payload_56_real = myFFT_3_fft_col_out_regNext_payload_56_real;
  assign io_line_out_payload_56_imag = myFFT_3_fft_col_out_regNext_payload_56_imag;
  assign io_line_out_payload_57_real = myFFT_3_fft_col_out_regNext_payload_57_real;
  assign io_line_out_payload_57_imag = myFFT_3_fft_col_out_regNext_payload_57_imag;
  assign io_line_out_payload_58_real = myFFT_3_fft_col_out_regNext_payload_58_real;
  assign io_line_out_payload_58_imag = myFFT_3_fft_col_out_regNext_payload_58_imag;
  assign io_line_out_payload_59_real = myFFT_3_fft_col_out_regNext_payload_59_real;
  assign io_line_out_payload_59_imag = myFFT_3_fft_col_out_regNext_payload_59_imag;
  assign io_line_out_payload_60_real = myFFT_3_fft_col_out_regNext_payload_60_real;
  assign io_line_out_payload_60_imag = myFFT_3_fft_col_out_regNext_payload_60_imag;
  assign io_line_out_payload_61_real = myFFT_3_fft_col_out_regNext_payload_61_real;
  assign io_line_out_payload_61_imag = myFFT_3_fft_col_out_regNext_payload_61_imag;
  assign io_line_out_payload_62_real = myFFT_3_fft_col_out_regNext_payload_62_real;
  assign io_line_out_payload_62_imag = myFFT_3_fft_col_out_regNext_payload_62_imag;
  assign io_line_out_payload_63_real = myFFT_3_fft_col_out_regNext_payload_63_real;
  assign io_line_out_payload_63_imag = myFFT_3_fft_col_out_regNext_payload_63_imag;
  always @ (posedge clk or posedge reset) begin
    if (reset) begin
      row_addr_value <= 6'h0;
      null_cnt_value <= 6'h0;
      null_cond_period_minus_1 <= 1'b0;
      null_cond_period_regNext <= 1'b0;
      myFFT_3_fft_col_out_regNext_valid <= 1'b0;
    end else begin
      row_addr_value <= row_addr_valueNext;
      null_cnt_value <= null_cnt_valueNext;
      if(row_addr_willOverflow)begin
        null_cond_period_minus_1 <= 1'b1;
      end else begin
        if(null_cnt_willOverflow)begin
          null_cond_period_minus_1 <= 1'b0;
        end
      end
      null_cond_period_regNext <= null_cond_period;
      myFFT_3_fft_col_out_regNext_valid <= myFFT_3_fft_col_out_valid;
    end
  end

  always @ (posedge clk) begin
    if(myFFT_2_fft_row_valid)begin
      if(_zz_2)begin
        img_reg_array_0_0_real <= _zz_66;
      end
      if(_zz_3)begin
        img_reg_array_1_0_real <= _zz_66;
      end
      if(_zz_4)begin
        img_reg_array_2_0_real <= _zz_66;
      end
      if(_zz_5)begin
        img_reg_array_3_0_real <= _zz_66;
      end
      if(_zz_6)begin
        img_reg_array_4_0_real <= _zz_66;
      end
      if(_zz_7)begin
        img_reg_array_5_0_real <= _zz_66;
      end
      if(_zz_8)begin
        img_reg_array_6_0_real <= _zz_66;
      end
      if(_zz_9)begin
        img_reg_array_7_0_real <= _zz_66;
      end
      if(_zz_10)begin
        img_reg_array_8_0_real <= _zz_66;
      end
      if(_zz_11)begin
        img_reg_array_9_0_real <= _zz_66;
      end
      if(_zz_12)begin
        img_reg_array_10_0_real <= _zz_66;
      end
      if(_zz_13)begin
        img_reg_array_11_0_real <= _zz_66;
      end
      if(_zz_14)begin
        img_reg_array_12_0_real <= _zz_66;
      end
      if(_zz_15)begin
        img_reg_array_13_0_real <= _zz_66;
      end
      if(_zz_16)begin
        img_reg_array_14_0_real <= _zz_66;
      end
      if(_zz_17)begin
        img_reg_array_15_0_real <= _zz_66;
      end
      if(_zz_18)begin
        img_reg_array_16_0_real <= _zz_66;
      end
      if(_zz_19)begin
        img_reg_array_17_0_real <= _zz_66;
      end
      if(_zz_20)begin
        img_reg_array_18_0_real <= _zz_66;
      end
      if(_zz_21)begin
        img_reg_array_19_0_real <= _zz_66;
      end
      if(_zz_22)begin
        img_reg_array_20_0_real <= _zz_66;
      end
      if(_zz_23)begin
        img_reg_array_21_0_real <= _zz_66;
      end
      if(_zz_24)begin
        img_reg_array_22_0_real <= _zz_66;
      end
      if(_zz_25)begin
        img_reg_array_23_0_real <= _zz_66;
      end
      if(_zz_26)begin
        img_reg_array_24_0_real <= _zz_66;
      end
      if(_zz_27)begin
        img_reg_array_25_0_real <= _zz_66;
      end
      if(_zz_28)begin
        img_reg_array_26_0_real <= _zz_66;
      end
      if(_zz_29)begin
        img_reg_array_27_0_real <= _zz_66;
      end
      if(_zz_30)begin
        img_reg_array_28_0_real <= _zz_66;
      end
      if(_zz_31)begin
        img_reg_array_29_0_real <= _zz_66;
      end
      if(_zz_32)begin
        img_reg_array_30_0_real <= _zz_66;
      end
      if(_zz_33)begin
        img_reg_array_31_0_real <= _zz_66;
      end
      if(_zz_34)begin
        img_reg_array_32_0_real <= _zz_66;
      end
      if(_zz_35)begin
        img_reg_array_33_0_real <= _zz_66;
      end
      if(_zz_36)begin
        img_reg_array_34_0_real <= _zz_66;
      end
      if(_zz_37)begin
        img_reg_array_35_0_real <= _zz_66;
      end
      if(_zz_38)begin
        img_reg_array_36_0_real <= _zz_66;
      end
      if(_zz_39)begin
        img_reg_array_37_0_real <= _zz_66;
      end
      if(_zz_40)begin
        img_reg_array_38_0_real <= _zz_66;
      end
      if(_zz_41)begin
        img_reg_array_39_0_real <= _zz_66;
      end
      if(_zz_42)begin
        img_reg_array_40_0_real <= _zz_66;
      end
      if(_zz_43)begin
        img_reg_array_41_0_real <= _zz_66;
      end
      if(_zz_44)begin
        img_reg_array_42_0_real <= _zz_66;
      end
      if(_zz_45)begin
        img_reg_array_43_0_real <= _zz_66;
      end
      if(_zz_46)begin
        img_reg_array_44_0_real <= _zz_66;
      end
      if(_zz_47)begin
        img_reg_array_45_0_real <= _zz_66;
      end
      if(_zz_48)begin
        img_reg_array_46_0_real <= _zz_66;
      end
      if(_zz_49)begin
        img_reg_array_47_0_real <= _zz_66;
      end
      if(_zz_50)begin
        img_reg_array_48_0_real <= _zz_66;
      end
      if(_zz_51)begin
        img_reg_array_49_0_real <= _zz_66;
      end
      if(_zz_52)begin
        img_reg_array_50_0_real <= _zz_66;
      end
      if(_zz_53)begin
        img_reg_array_51_0_real <= _zz_66;
      end
      if(_zz_54)begin
        img_reg_array_52_0_real <= _zz_66;
      end
      if(_zz_55)begin
        img_reg_array_53_0_real <= _zz_66;
      end
      if(_zz_56)begin
        img_reg_array_54_0_real <= _zz_66;
      end
      if(_zz_57)begin
        img_reg_array_55_0_real <= _zz_66;
      end
      if(_zz_58)begin
        img_reg_array_56_0_real <= _zz_66;
      end
      if(_zz_59)begin
        img_reg_array_57_0_real <= _zz_66;
      end
      if(_zz_60)begin
        img_reg_array_58_0_real <= _zz_66;
      end
      if(_zz_61)begin
        img_reg_array_59_0_real <= _zz_66;
      end
      if(_zz_62)begin
        img_reg_array_60_0_real <= _zz_66;
      end
      if(_zz_63)begin
        img_reg_array_61_0_real <= _zz_66;
      end
      if(_zz_64)begin
        img_reg_array_62_0_real <= _zz_66;
      end
      if(_zz_65)begin
        img_reg_array_63_0_real <= _zz_66;
      end
      if(_zz_2)begin
        img_reg_array_0_0_imag <= _zz_67;
      end
      if(_zz_3)begin
        img_reg_array_1_0_imag <= _zz_67;
      end
      if(_zz_4)begin
        img_reg_array_2_0_imag <= _zz_67;
      end
      if(_zz_5)begin
        img_reg_array_3_0_imag <= _zz_67;
      end
      if(_zz_6)begin
        img_reg_array_4_0_imag <= _zz_67;
      end
      if(_zz_7)begin
        img_reg_array_5_0_imag <= _zz_67;
      end
      if(_zz_8)begin
        img_reg_array_6_0_imag <= _zz_67;
      end
      if(_zz_9)begin
        img_reg_array_7_0_imag <= _zz_67;
      end
      if(_zz_10)begin
        img_reg_array_8_0_imag <= _zz_67;
      end
      if(_zz_11)begin
        img_reg_array_9_0_imag <= _zz_67;
      end
      if(_zz_12)begin
        img_reg_array_10_0_imag <= _zz_67;
      end
      if(_zz_13)begin
        img_reg_array_11_0_imag <= _zz_67;
      end
      if(_zz_14)begin
        img_reg_array_12_0_imag <= _zz_67;
      end
      if(_zz_15)begin
        img_reg_array_13_0_imag <= _zz_67;
      end
      if(_zz_16)begin
        img_reg_array_14_0_imag <= _zz_67;
      end
      if(_zz_17)begin
        img_reg_array_15_0_imag <= _zz_67;
      end
      if(_zz_18)begin
        img_reg_array_16_0_imag <= _zz_67;
      end
      if(_zz_19)begin
        img_reg_array_17_0_imag <= _zz_67;
      end
      if(_zz_20)begin
        img_reg_array_18_0_imag <= _zz_67;
      end
      if(_zz_21)begin
        img_reg_array_19_0_imag <= _zz_67;
      end
      if(_zz_22)begin
        img_reg_array_20_0_imag <= _zz_67;
      end
      if(_zz_23)begin
        img_reg_array_21_0_imag <= _zz_67;
      end
      if(_zz_24)begin
        img_reg_array_22_0_imag <= _zz_67;
      end
      if(_zz_25)begin
        img_reg_array_23_0_imag <= _zz_67;
      end
      if(_zz_26)begin
        img_reg_array_24_0_imag <= _zz_67;
      end
      if(_zz_27)begin
        img_reg_array_25_0_imag <= _zz_67;
      end
      if(_zz_28)begin
        img_reg_array_26_0_imag <= _zz_67;
      end
      if(_zz_29)begin
        img_reg_array_27_0_imag <= _zz_67;
      end
      if(_zz_30)begin
        img_reg_array_28_0_imag <= _zz_67;
      end
      if(_zz_31)begin
        img_reg_array_29_0_imag <= _zz_67;
      end
      if(_zz_32)begin
        img_reg_array_30_0_imag <= _zz_67;
      end
      if(_zz_33)begin
        img_reg_array_31_0_imag <= _zz_67;
      end
      if(_zz_34)begin
        img_reg_array_32_0_imag <= _zz_67;
      end
      if(_zz_35)begin
        img_reg_array_33_0_imag <= _zz_67;
      end
      if(_zz_36)begin
        img_reg_array_34_0_imag <= _zz_67;
      end
      if(_zz_37)begin
        img_reg_array_35_0_imag <= _zz_67;
      end
      if(_zz_38)begin
        img_reg_array_36_0_imag <= _zz_67;
      end
      if(_zz_39)begin
        img_reg_array_37_0_imag <= _zz_67;
      end
      if(_zz_40)begin
        img_reg_array_38_0_imag <= _zz_67;
      end
      if(_zz_41)begin
        img_reg_array_39_0_imag <= _zz_67;
      end
      if(_zz_42)begin
        img_reg_array_40_0_imag <= _zz_67;
      end
      if(_zz_43)begin
        img_reg_array_41_0_imag <= _zz_67;
      end
      if(_zz_44)begin
        img_reg_array_42_0_imag <= _zz_67;
      end
      if(_zz_45)begin
        img_reg_array_43_0_imag <= _zz_67;
      end
      if(_zz_46)begin
        img_reg_array_44_0_imag <= _zz_67;
      end
      if(_zz_47)begin
        img_reg_array_45_0_imag <= _zz_67;
      end
      if(_zz_48)begin
        img_reg_array_46_0_imag <= _zz_67;
      end
      if(_zz_49)begin
        img_reg_array_47_0_imag <= _zz_67;
      end
      if(_zz_50)begin
        img_reg_array_48_0_imag <= _zz_67;
      end
      if(_zz_51)begin
        img_reg_array_49_0_imag <= _zz_67;
      end
      if(_zz_52)begin
        img_reg_array_50_0_imag <= _zz_67;
      end
      if(_zz_53)begin
        img_reg_array_51_0_imag <= _zz_67;
      end
      if(_zz_54)begin
        img_reg_array_52_0_imag <= _zz_67;
      end
      if(_zz_55)begin
        img_reg_array_53_0_imag <= _zz_67;
      end
      if(_zz_56)begin
        img_reg_array_54_0_imag <= _zz_67;
      end
      if(_zz_57)begin
        img_reg_array_55_0_imag <= _zz_67;
      end
      if(_zz_58)begin
        img_reg_array_56_0_imag <= _zz_67;
      end
      if(_zz_59)begin
        img_reg_array_57_0_imag <= _zz_67;
      end
      if(_zz_60)begin
        img_reg_array_58_0_imag <= _zz_67;
      end
      if(_zz_61)begin
        img_reg_array_59_0_imag <= _zz_67;
      end
      if(_zz_62)begin
        img_reg_array_60_0_imag <= _zz_67;
      end
      if(_zz_63)begin
        img_reg_array_61_0_imag <= _zz_67;
      end
      if(_zz_64)begin
        img_reg_array_62_0_imag <= _zz_67;
      end
      if(_zz_65)begin
        img_reg_array_63_0_imag <= _zz_67;
      end
      if(_zz_2)begin
        img_reg_array_0_1_real <= _zz_68;
      end
      if(_zz_3)begin
        img_reg_array_1_1_real <= _zz_68;
      end
      if(_zz_4)begin
        img_reg_array_2_1_real <= _zz_68;
      end
      if(_zz_5)begin
        img_reg_array_3_1_real <= _zz_68;
      end
      if(_zz_6)begin
        img_reg_array_4_1_real <= _zz_68;
      end
      if(_zz_7)begin
        img_reg_array_5_1_real <= _zz_68;
      end
      if(_zz_8)begin
        img_reg_array_6_1_real <= _zz_68;
      end
      if(_zz_9)begin
        img_reg_array_7_1_real <= _zz_68;
      end
      if(_zz_10)begin
        img_reg_array_8_1_real <= _zz_68;
      end
      if(_zz_11)begin
        img_reg_array_9_1_real <= _zz_68;
      end
      if(_zz_12)begin
        img_reg_array_10_1_real <= _zz_68;
      end
      if(_zz_13)begin
        img_reg_array_11_1_real <= _zz_68;
      end
      if(_zz_14)begin
        img_reg_array_12_1_real <= _zz_68;
      end
      if(_zz_15)begin
        img_reg_array_13_1_real <= _zz_68;
      end
      if(_zz_16)begin
        img_reg_array_14_1_real <= _zz_68;
      end
      if(_zz_17)begin
        img_reg_array_15_1_real <= _zz_68;
      end
      if(_zz_18)begin
        img_reg_array_16_1_real <= _zz_68;
      end
      if(_zz_19)begin
        img_reg_array_17_1_real <= _zz_68;
      end
      if(_zz_20)begin
        img_reg_array_18_1_real <= _zz_68;
      end
      if(_zz_21)begin
        img_reg_array_19_1_real <= _zz_68;
      end
      if(_zz_22)begin
        img_reg_array_20_1_real <= _zz_68;
      end
      if(_zz_23)begin
        img_reg_array_21_1_real <= _zz_68;
      end
      if(_zz_24)begin
        img_reg_array_22_1_real <= _zz_68;
      end
      if(_zz_25)begin
        img_reg_array_23_1_real <= _zz_68;
      end
      if(_zz_26)begin
        img_reg_array_24_1_real <= _zz_68;
      end
      if(_zz_27)begin
        img_reg_array_25_1_real <= _zz_68;
      end
      if(_zz_28)begin
        img_reg_array_26_1_real <= _zz_68;
      end
      if(_zz_29)begin
        img_reg_array_27_1_real <= _zz_68;
      end
      if(_zz_30)begin
        img_reg_array_28_1_real <= _zz_68;
      end
      if(_zz_31)begin
        img_reg_array_29_1_real <= _zz_68;
      end
      if(_zz_32)begin
        img_reg_array_30_1_real <= _zz_68;
      end
      if(_zz_33)begin
        img_reg_array_31_1_real <= _zz_68;
      end
      if(_zz_34)begin
        img_reg_array_32_1_real <= _zz_68;
      end
      if(_zz_35)begin
        img_reg_array_33_1_real <= _zz_68;
      end
      if(_zz_36)begin
        img_reg_array_34_1_real <= _zz_68;
      end
      if(_zz_37)begin
        img_reg_array_35_1_real <= _zz_68;
      end
      if(_zz_38)begin
        img_reg_array_36_1_real <= _zz_68;
      end
      if(_zz_39)begin
        img_reg_array_37_1_real <= _zz_68;
      end
      if(_zz_40)begin
        img_reg_array_38_1_real <= _zz_68;
      end
      if(_zz_41)begin
        img_reg_array_39_1_real <= _zz_68;
      end
      if(_zz_42)begin
        img_reg_array_40_1_real <= _zz_68;
      end
      if(_zz_43)begin
        img_reg_array_41_1_real <= _zz_68;
      end
      if(_zz_44)begin
        img_reg_array_42_1_real <= _zz_68;
      end
      if(_zz_45)begin
        img_reg_array_43_1_real <= _zz_68;
      end
      if(_zz_46)begin
        img_reg_array_44_1_real <= _zz_68;
      end
      if(_zz_47)begin
        img_reg_array_45_1_real <= _zz_68;
      end
      if(_zz_48)begin
        img_reg_array_46_1_real <= _zz_68;
      end
      if(_zz_49)begin
        img_reg_array_47_1_real <= _zz_68;
      end
      if(_zz_50)begin
        img_reg_array_48_1_real <= _zz_68;
      end
      if(_zz_51)begin
        img_reg_array_49_1_real <= _zz_68;
      end
      if(_zz_52)begin
        img_reg_array_50_1_real <= _zz_68;
      end
      if(_zz_53)begin
        img_reg_array_51_1_real <= _zz_68;
      end
      if(_zz_54)begin
        img_reg_array_52_1_real <= _zz_68;
      end
      if(_zz_55)begin
        img_reg_array_53_1_real <= _zz_68;
      end
      if(_zz_56)begin
        img_reg_array_54_1_real <= _zz_68;
      end
      if(_zz_57)begin
        img_reg_array_55_1_real <= _zz_68;
      end
      if(_zz_58)begin
        img_reg_array_56_1_real <= _zz_68;
      end
      if(_zz_59)begin
        img_reg_array_57_1_real <= _zz_68;
      end
      if(_zz_60)begin
        img_reg_array_58_1_real <= _zz_68;
      end
      if(_zz_61)begin
        img_reg_array_59_1_real <= _zz_68;
      end
      if(_zz_62)begin
        img_reg_array_60_1_real <= _zz_68;
      end
      if(_zz_63)begin
        img_reg_array_61_1_real <= _zz_68;
      end
      if(_zz_64)begin
        img_reg_array_62_1_real <= _zz_68;
      end
      if(_zz_65)begin
        img_reg_array_63_1_real <= _zz_68;
      end
      if(_zz_2)begin
        img_reg_array_0_1_imag <= _zz_69;
      end
      if(_zz_3)begin
        img_reg_array_1_1_imag <= _zz_69;
      end
      if(_zz_4)begin
        img_reg_array_2_1_imag <= _zz_69;
      end
      if(_zz_5)begin
        img_reg_array_3_1_imag <= _zz_69;
      end
      if(_zz_6)begin
        img_reg_array_4_1_imag <= _zz_69;
      end
      if(_zz_7)begin
        img_reg_array_5_1_imag <= _zz_69;
      end
      if(_zz_8)begin
        img_reg_array_6_1_imag <= _zz_69;
      end
      if(_zz_9)begin
        img_reg_array_7_1_imag <= _zz_69;
      end
      if(_zz_10)begin
        img_reg_array_8_1_imag <= _zz_69;
      end
      if(_zz_11)begin
        img_reg_array_9_1_imag <= _zz_69;
      end
      if(_zz_12)begin
        img_reg_array_10_1_imag <= _zz_69;
      end
      if(_zz_13)begin
        img_reg_array_11_1_imag <= _zz_69;
      end
      if(_zz_14)begin
        img_reg_array_12_1_imag <= _zz_69;
      end
      if(_zz_15)begin
        img_reg_array_13_1_imag <= _zz_69;
      end
      if(_zz_16)begin
        img_reg_array_14_1_imag <= _zz_69;
      end
      if(_zz_17)begin
        img_reg_array_15_1_imag <= _zz_69;
      end
      if(_zz_18)begin
        img_reg_array_16_1_imag <= _zz_69;
      end
      if(_zz_19)begin
        img_reg_array_17_1_imag <= _zz_69;
      end
      if(_zz_20)begin
        img_reg_array_18_1_imag <= _zz_69;
      end
      if(_zz_21)begin
        img_reg_array_19_1_imag <= _zz_69;
      end
      if(_zz_22)begin
        img_reg_array_20_1_imag <= _zz_69;
      end
      if(_zz_23)begin
        img_reg_array_21_1_imag <= _zz_69;
      end
      if(_zz_24)begin
        img_reg_array_22_1_imag <= _zz_69;
      end
      if(_zz_25)begin
        img_reg_array_23_1_imag <= _zz_69;
      end
      if(_zz_26)begin
        img_reg_array_24_1_imag <= _zz_69;
      end
      if(_zz_27)begin
        img_reg_array_25_1_imag <= _zz_69;
      end
      if(_zz_28)begin
        img_reg_array_26_1_imag <= _zz_69;
      end
      if(_zz_29)begin
        img_reg_array_27_1_imag <= _zz_69;
      end
      if(_zz_30)begin
        img_reg_array_28_1_imag <= _zz_69;
      end
      if(_zz_31)begin
        img_reg_array_29_1_imag <= _zz_69;
      end
      if(_zz_32)begin
        img_reg_array_30_1_imag <= _zz_69;
      end
      if(_zz_33)begin
        img_reg_array_31_1_imag <= _zz_69;
      end
      if(_zz_34)begin
        img_reg_array_32_1_imag <= _zz_69;
      end
      if(_zz_35)begin
        img_reg_array_33_1_imag <= _zz_69;
      end
      if(_zz_36)begin
        img_reg_array_34_1_imag <= _zz_69;
      end
      if(_zz_37)begin
        img_reg_array_35_1_imag <= _zz_69;
      end
      if(_zz_38)begin
        img_reg_array_36_1_imag <= _zz_69;
      end
      if(_zz_39)begin
        img_reg_array_37_1_imag <= _zz_69;
      end
      if(_zz_40)begin
        img_reg_array_38_1_imag <= _zz_69;
      end
      if(_zz_41)begin
        img_reg_array_39_1_imag <= _zz_69;
      end
      if(_zz_42)begin
        img_reg_array_40_1_imag <= _zz_69;
      end
      if(_zz_43)begin
        img_reg_array_41_1_imag <= _zz_69;
      end
      if(_zz_44)begin
        img_reg_array_42_1_imag <= _zz_69;
      end
      if(_zz_45)begin
        img_reg_array_43_1_imag <= _zz_69;
      end
      if(_zz_46)begin
        img_reg_array_44_1_imag <= _zz_69;
      end
      if(_zz_47)begin
        img_reg_array_45_1_imag <= _zz_69;
      end
      if(_zz_48)begin
        img_reg_array_46_1_imag <= _zz_69;
      end
      if(_zz_49)begin
        img_reg_array_47_1_imag <= _zz_69;
      end
      if(_zz_50)begin
        img_reg_array_48_1_imag <= _zz_69;
      end
      if(_zz_51)begin
        img_reg_array_49_1_imag <= _zz_69;
      end
      if(_zz_52)begin
        img_reg_array_50_1_imag <= _zz_69;
      end
      if(_zz_53)begin
        img_reg_array_51_1_imag <= _zz_69;
      end
      if(_zz_54)begin
        img_reg_array_52_1_imag <= _zz_69;
      end
      if(_zz_55)begin
        img_reg_array_53_1_imag <= _zz_69;
      end
      if(_zz_56)begin
        img_reg_array_54_1_imag <= _zz_69;
      end
      if(_zz_57)begin
        img_reg_array_55_1_imag <= _zz_69;
      end
      if(_zz_58)begin
        img_reg_array_56_1_imag <= _zz_69;
      end
      if(_zz_59)begin
        img_reg_array_57_1_imag <= _zz_69;
      end
      if(_zz_60)begin
        img_reg_array_58_1_imag <= _zz_69;
      end
      if(_zz_61)begin
        img_reg_array_59_1_imag <= _zz_69;
      end
      if(_zz_62)begin
        img_reg_array_60_1_imag <= _zz_69;
      end
      if(_zz_63)begin
        img_reg_array_61_1_imag <= _zz_69;
      end
      if(_zz_64)begin
        img_reg_array_62_1_imag <= _zz_69;
      end
      if(_zz_65)begin
        img_reg_array_63_1_imag <= _zz_69;
      end
      if(_zz_2)begin
        img_reg_array_0_2_real <= _zz_70;
      end
      if(_zz_3)begin
        img_reg_array_1_2_real <= _zz_70;
      end
      if(_zz_4)begin
        img_reg_array_2_2_real <= _zz_70;
      end
      if(_zz_5)begin
        img_reg_array_3_2_real <= _zz_70;
      end
      if(_zz_6)begin
        img_reg_array_4_2_real <= _zz_70;
      end
      if(_zz_7)begin
        img_reg_array_5_2_real <= _zz_70;
      end
      if(_zz_8)begin
        img_reg_array_6_2_real <= _zz_70;
      end
      if(_zz_9)begin
        img_reg_array_7_2_real <= _zz_70;
      end
      if(_zz_10)begin
        img_reg_array_8_2_real <= _zz_70;
      end
      if(_zz_11)begin
        img_reg_array_9_2_real <= _zz_70;
      end
      if(_zz_12)begin
        img_reg_array_10_2_real <= _zz_70;
      end
      if(_zz_13)begin
        img_reg_array_11_2_real <= _zz_70;
      end
      if(_zz_14)begin
        img_reg_array_12_2_real <= _zz_70;
      end
      if(_zz_15)begin
        img_reg_array_13_2_real <= _zz_70;
      end
      if(_zz_16)begin
        img_reg_array_14_2_real <= _zz_70;
      end
      if(_zz_17)begin
        img_reg_array_15_2_real <= _zz_70;
      end
      if(_zz_18)begin
        img_reg_array_16_2_real <= _zz_70;
      end
      if(_zz_19)begin
        img_reg_array_17_2_real <= _zz_70;
      end
      if(_zz_20)begin
        img_reg_array_18_2_real <= _zz_70;
      end
      if(_zz_21)begin
        img_reg_array_19_2_real <= _zz_70;
      end
      if(_zz_22)begin
        img_reg_array_20_2_real <= _zz_70;
      end
      if(_zz_23)begin
        img_reg_array_21_2_real <= _zz_70;
      end
      if(_zz_24)begin
        img_reg_array_22_2_real <= _zz_70;
      end
      if(_zz_25)begin
        img_reg_array_23_2_real <= _zz_70;
      end
      if(_zz_26)begin
        img_reg_array_24_2_real <= _zz_70;
      end
      if(_zz_27)begin
        img_reg_array_25_2_real <= _zz_70;
      end
      if(_zz_28)begin
        img_reg_array_26_2_real <= _zz_70;
      end
      if(_zz_29)begin
        img_reg_array_27_2_real <= _zz_70;
      end
      if(_zz_30)begin
        img_reg_array_28_2_real <= _zz_70;
      end
      if(_zz_31)begin
        img_reg_array_29_2_real <= _zz_70;
      end
      if(_zz_32)begin
        img_reg_array_30_2_real <= _zz_70;
      end
      if(_zz_33)begin
        img_reg_array_31_2_real <= _zz_70;
      end
      if(_zz_34)begin
        img_reg_array_32_2_real <= _zz_70;
      end
      if(_zz_35)begin
        img_reg_array_33_2_real <= _zz_70;
      end
      if(_zz_36)begin
        img_reg_array_34_2_real <= _zz_70;
      end
      if(_zz_37)begin
        img_reg_array_35_2_real <= _zz_70;
      end
      if(_zz_38)begin
        img_reg_array_36_2_real <= _zz_70;
      end
      if(_zz_39)begin
        img_reg_array_37_2_real <= _zz_70;
      end
      if(_zz_40)begin
        img_reg_array_38_2_real <= _zz_70;
      end
      if(_zz_41)begin
        img_reg_array_39_2_real <= _zz_70;
      end
      if(_zz_42)begin
        img_reg_array_40_2_real <= _zz_70;
      end
      if(_zz_43)begin
        img_reg_array_41_2_real <= _zz_70;
      end
      if(_zz_44)begin
        img_reg_array_42_2_real <= _zz_70;
      end
      if(_zz_45)begin
        img_reg_array_43_2_real <= _zz_70;
      end
      if(_zz_46)begin
        img_reg_array_44_2_real <= _zz_70;
      end
      if(_zz_47)begin
        img_reg_array_45_2_real <= _zz_70;
      end
      if(_zz_48)begin
        img_reg_array_46_2_real <= _zz_70;
      end
      if(_zz_49)begin
        img_reg_array_47_2_real <= _zz_70;
      end
      if(_zz_50)begin
        img_reg_array_48_2_real <= _zz_70;
      end
      if(_zz_51)begin
        img_reg_array_49_2_real <= _zz_70;
      end
      if(_zz_52)begin
        img_reg_array_50_2_real <= _zz_70;
      end
      if(_zz_53)begin
        img_reg_array_51_2_real <= _zz_70;
      end
      if(_zz_54)begin
        img_reg_array_52_2_real <= _zz_70;
      end
      if(_zz_55)begin
        img_reg_array_53_2_real <= _zz_70;
      end
      if(_zz_56)begin
        img_reg_array_54_2_real <= _zz_70;
      end
      if(_zz_57)begin
        img_reg_array_55_2_real <= _zz_70;
      end
      if(_zz_58)begin
        img_reg_array_56_2_real <= _zz_70;
      end
      if(_zz_59)begin
        img_reg_array_57_2_real <= _zz_70;
      end
      if(_zz_60)begin
        img_reg_array_58_2_real <= _zz_70;
      end
      if(_zz_61)begin
        img_reg_array_59_2_real <= _zz_70;
      end
      if(_zz_62)begin
        img_reg_array_60_2_real <= _zz_70;
      end
      if(_zz_63)begin
        img_reg_array_61_2_real <= _zz_70;
      end
      if(_zz_64)begin
        img_reg_array_62_2_real <= _zz_70;
      end
      if(_zz_65)begin
        img_reg_array_63_2_real <= _zz_70;
      end
      if(_zz_2)begin
        img_reg_array_0_2_imag <= _zz_71;
      end
      if(_zz_3)begin
        img_reg_array_1_2_imag <= _zz_71;
      end
      if(_zz_4)begin
        img_reg_array_2_2_imag <= _zz_71;
      end
      if(_zz_5)begin
        img_reg_array_3_2_imag <= _zz_71;
      end
      if(_zz_6)begin
        img_reg_array_4_2_imag <= _zz_71;
      end
      if(_zz_7)begin
        img_reg_array_5_2_imag <= _zz_71;
      end
      if(_zz_8)begin
        img_reg_array_6_2_imag <= _zz_71;
      end
      if(_zz_9)begin
        img_reg_array_7_2_imag <= _zz_71;
      end
      if(_zz_10)begin
        img_reg_array_8_2_imag <= _zz_71;
      end
      if(_zz_11)begin
        img_reg_array_9_2_imag <= _zz_71;
      end
      if(_zz_12)begin
        img_reg_array_10_2_imag <= _zz_71;
      end
      if(_zz_13)begin
        img_reg_array_11_2_imag <= _zz_71;
      end
      if(_zz_14)begin
        img_reg_array_12_2_imag <= _zz_71;
      end
      if(_zz_15)begin
        img_reg_array_13_2_imag <= _zz_71;
      end
      if(_zz_16)begin
        img_reg_array_14_2_imag <= _zz_71;
      end
      if(_zz_17)begin
        img_reg_array_15_2_imag <= _zz_71;
      end
      if(_zz_18)begin
        img_reg_array_16_2_imag <= _zz_71;
      end
      if(_zz_19)begin
        img_reg_array_17_2_imag <= _zz_71;
      end
      if(_zz_20)begin
        img_reg_array_18_2_imag <= _zz_71;
      end
      if(_zz_21)begin
        img_reg_array_19_2_imag <= _zz_71;
      end
      if(_zz_22)begin
        img_reg_array_20_2_imag <= _zz_71;
      end
      if(_zz_23)begin
        img_reg_array_21_2_imag <= _zz_71;
      end
      if(_zz_24)begin
        img_reg_array_22_2_imag <= _zz_71;
      end
      if(_zz_25)begin
        img_reg_array_23_2_imag <= _zz_71;
      end
      if(_zz_26)begin
        img_reg_array_24_2_imag <= _zz_71;
      end
      if(_zz_27)begin
        img_reg_array_25_2_imag <= _zz_71;
      end
      if(_zz_28)begin
        img_reg_array_26_2_imag <= _zz_71;
      end
      if(_zz_29)begin
        img_reg_array_27_2_imag <= _zz_71;
      end
      if(_zz_30)begin
        img_reg_array_28_2_imag <= _zz_71;
      end
      if(_zz_31)begin
        img_reg_array_29_2_imag <= _zz_71;
      end
      if(_zz_32)begin
        img_reg_array_30_2_imag <= _zz_71;
      end
      if(_zz_33)begin
        img_reg_array_31_2_imag <= _zz_71;
      end
      if(_zz_34)begin
        img_reg_array_32_2_imag <= _zz_71;
      end
      if(_zz_35)begin
        img_reg_array_33_2_imag <= _zz_71;
      end
      if(_zz_36)begin
        img_reg_array_34_2_imag <= _zz_71;
      end
      if(_zz_37)begin
        img_reg_array_35_2_imag <= _zz_71;
      end
      if(_zz_38)begin
        img_reg_array_36_2_imag <= _zz_71;
      end
      if(_zz_39)begin
        img_reg_array_37_2_imag <= _zz_71;
      end
      if(_zz_40)begin
        img_reg_array_38_2_imag <= _zz_71;
      end
      if(_zz_41)begin
        img_reg_array_39_2_imag <= _zz_71;
      end
      if(_zz_42)begin
        img_reg_array_40_2_imag <= _zz_71;
      end
      if(_zz_43)begin
        img_reg_array_41_2_imag <= _zz_71;
      end
      if(_zz_44)begin
        img_reg_array_42_2_imag <= _zz_71;
      end
      if(_zz_45)begin
        img_reg_array_43_2_imag <= _zz_71;
      end
      if(_zz_46)begin
        img_reg_array_44_2_imag <= _zz_71;
      end
      if(_zz_47)begin
        img_reg_array_45_2_imag <= _zz_71;
      end
      if(_zz_48)begin
        img_reg_array_46_2_imag <= _zz_71;
      end
      if(_zz_49)begin
        img_reg_array_47_2_imag <= _zz_71;
      end
      if(_zz_50)begin
        img_reg_array_48_2_imag <= _zz_71;
      end
      if(_zz_51)begin
        img_reg_array_49_2_imag <= _zz_71;
      end
      if(_zz_52)begin
        img_reg_array_50_2_imag <= _zz_71;
      end
      if(_zz_53)begin
        img_reg_array_51_2_imag <= _zz_71;
      end
      if(_zz_54)begin
        img_reg_array_52_2_imag <= _zz_71;
      end
      if(_zz_55)begin
        img_reg_array_53_2_imag <= _zz_71;
      end
      if(_zz_56)begin
        img_reg_array_54_2_imag <= _zz_71;
      end
      if(_zz_57)begin
        img_reg_array_55_2_imag <= _zz_71;
      end
      if(_zz_58)begin
        img_reg_array_56_2_imag <= _zz_71;
      end
      if(_zz_59)begin
        img_reg_array_57_2_imag <= _zz_71;
      end
      if(_zz_60)begin
        img_reg_array_58_2_imag <= _zz_71;
      end
      if(_zz_61)begin
        img_reg_array_59_2_imag <= _zz_71;
      end
      if(_zz_62)begin
        img_reg_array_60_2_imag <= _zz_71;
      end
      if(_zz_63)begin
        img_reg_array_61_2_imag <= _zz_71;
      end
      if(_zz_64)begin
        img_reg_array_62_2_imag <= _zz_71;
      end
      if(_zz_65)begin
        img_reg_array_63_2_imag <= _zz_71;
      end
      if(_zz_2)begin
        img_reg_array_0_3_real <= _zz_72;
      end
      if(_zz_3)begin
        img_reg_array_1_3_real <= _zz_72;
      end
      if(_zz_4)begin
        img_reg_array_2_3_real <= _zz_72;
      end
      if(_zz_5)begin
        img_reg_array_3_3_real <= _zz_72;
      end
      if(_zz_6)begin
        img_reg_array_4_3_real <= _zz_72;
      end
      if(_zz_7)begin
        img_reg_array_5_3_real <= _zz_72;
      end
      if(_zz_8)begin
        img_reg_array_6_3_real <= _zz_72;
      end
      if(_zz_9)begin
        img_reg_array_7_3_real <= _zz_72;
      end
      if(_zz_10)begin
        img_reg_array_8_3_real <= _zz_72;
      end
      if(_zz_11)begin
        img_reg_array_9_3_real <= _zz_72;
      end
      if(_zz_12)begin
        img_reg_array_10_3_real <= _zz_72;
      end
      if(_zz_13)begin
        img_reg_array_11_3_real <= _zz_72;
      end
      if(_zz_14)begin
        img_reg_array_12_3_real <= _zz_72;
      end
      if(_zz_15)begin
        img_reg_array_13_3_real <= _zz_72;
      end
      if(_zz_16)begin
        img_reg_array_14_3_real <= _zz_72;
      end
      if(_zz_17)begin
        img_reg_array_15_3_real <= _zz_72;
      end
      if(_zz_18)begin
        img_reg_array_16_3_real <= _zz_72;
      end
      if(_zz_19)begin
        img_reg_array_17_3_real <= _zz_72;
      end
      if(_zz_20)begin
        img_reg_array_18_3_real <= _zz_72;
      end
      if(_zz_21)begin
        img_reg_array_19_3_real <= _zz_72;
      end
      if(_zz_22)begin
        img_reg_array_20_3_real <= _zz_72;
      end
      if(_zz_23)begin
        img_reg_array_21_3_real <= _zz_72;
      end
      if(_zz_24)begin
        img_reg_array_22_3_real <= _zz_72;
      end
      if(_zz_25)begin
        img_reg_array_23_3_real <= _zz_72;
      end
      if(_zz_26)begin
        img_reg_array_24_3_real <= _zz_72;
      end
      if(_zz_27)begin
        img_reg_array_25_3_real <= _zz_72;
      end
      if(_zz_28)begin
        img_reg_array_26_3_real <= _zz_72;
      end
      if(_zz_29)begin
        img_reg_array_27_3_real <= _zz_72;
      end
      if(_zz_30)begin
        img_reg_array_28_3_real <= _zz_72;
      end
      if(_zz_31)begin
        img_reg_array_29_3_real <= _zz_72;
      end
      if(_zz_32)begin
        img_reg_array_30_3_real <= _zz_72;
      end
      if(_zz_33)begin
        img_reg_array_31_3_real <= _zz_72;
      end
      if(_zz_34)begin
        img_reg_array_32_3_real <= _zz_72;
      end
      if(_zz_35)begin
        img_reg_array_33_3_real <= _zz_72;
      end
      if(_zz_36)begin
        img_reg_array_34_3_real <= _zz_72;
      end
      if(_zz_37)begin
        img_reg_array_35_3_real <= _zz_72;
      end
      if(_zz_38)begin
        img_reg_array_36_3_real <= _zz_72;
      end
      if(_zz_39)begin
        img_reg_array_37_3_real <= _zz_72;
      end
      if(_zz_40)begin
        img_reg_array_38_3_real <= _zz_72;
      end
      if(_zz_41)begin
        img_reg_array_39_3_real <= _zz_72;
      end
      if(_zz_42)begin
        img_reg_array_40_3_real <= _zz_72;
      end
      if(_zz_43)begin
        img_reg_array_41_3_real <= _zz_72;
      end
      if(_zz_44)begin
        img_reg_array_42_3_real <= _zz_72;
      end
      if(_zz_45)begin
        img_reg_array_43_3_real <= _zz_72;
      end
      if(_zz_46)begin
        img_reg_array_44_3_real <= _zz_72;
      end
      if(_zz_47)begin
        img_reg_array_45_3_real <= _zz_72;
      end
      if(_zz_48)begin
        img_reg_array_46_3_real <= _zz_72;
      end
      if(_zz_49)begin
        img_reg_array_47_3_real <= _zz_72;
      end
      if(_zz_50)begin
        img_reg_array_48_3_real <= _zz_72;
      end
      if(_zz_51)begin
        img_reg_array_49_3_real <= _zz_72;
      end
      if(_zz_52)begin
        img_reg_array_50_3_real <= _zz_72;
      end
      if(_zz_53)begin
        img_reg_array_51_3_real <= _zz_72;
      end
      if(_zz_54)begin
        img_reg_array_52_3_real <= _zz_72;
      end
      if(_zz_55)begin
        img_reg_array_53_3_real <= _zz_72;
      end
      if(_zz_56)begin
        img_reg_array_54_3_real <= _zz_72;
      end
      if(_zz_57)begin
        img_reg_array_55_3_real <= _zz_72;
      end
      if(_zz_58)begin
        img_reg_array_56_3_real <= _zz_72;
      end
      if(_zz_59)begin
        img_reg_array_57_3_real <= _zz_72;
      end
      if(_zz_60)begin
        img_reg_array_58_3_real <= _zz_72;
      end
      if(_zz_61)begin
        img_reg_array_59_3_real <= _zz_72;
      end
      if(_zz_62)begin
        img_reg_array_60_3_real <= _zz_72;
      end
      if(_zz_63)begin
        img_reg_array_61_3_real <= _zz_72;
      end
      if(_zz_64)begin
        img_reg_array_62_3_real <= _zz_72;
      end
      if(_zz_65)begin
        img_reg_array_63_3_real <= _zz_72;
      end
      if(_zz_2)begin
        img_reg_array_0_3_imag <= _zz_73;
      end
      if(_zz_3)begin
        img_reg_array_1_3_imag <= _zz_73;
      end
      if(_zz_4)begin
        img_reg_array_2_3_imag <= _zz_73;
      end
      if(_zz_5)begin
        img_reg_array_3_3_imag <= _zz_73;
      end
      if(_zz_6)begin
        img_reg_array_4_3_imag <= _zz_73;
      end
      if(_zz_7)begin
        img_reg_array_5_3_imag <= _zz_73;
      end
      if(_zz_8)begin
        img_reg_array_6_3_imag <= _zz_73;
      end
      if(_zz_9)begin
        img_reg_array_7_3_imag <= _zz_73;
      end
      if(_zz_10)begin
        img_reg_array_8_3_imag <= _zz_73;
      end
      if(_zz_11)begin
        img_reg_array_9_3_imag <= _zz_73;
      end
      if(_zz_12)begin
        img_reg_array_10_3_imag <= _zz_73;
      end
      if(_zz_13)begin
        img_reg_array_11_3_imag <= _zz_73;
      end
      if(_zz_14)begin
        img_reg_array_12_3_imag <= _zz_73;
      end
      if(_zz_15)begin
        img_reg_array_13_3_imag <= _zz_73;
      end
      if(_zz_16)begin
        img_reg_array_14_3_imag <= _zz_73;
      end
      if(_zz_17)begin
        img_reg_array_15_3_imag <= _zz_73;
      end
      if(_zz_18)begin
        img_reg_array_16_3_imag <= _zz_73;
      end
      if(_zz_19)begin
        img_reg_array_17_3_imag <= _zz_73;
      end
      if(_zz_20)begin
        img_reg_array_18_3_imag <= _zz_73;
      end
      if(_zz_21)begin
        img_reg_array_19_3_imag <= _zz_73;
      end
      if(_zz_22)begin
        img_reg_array_20_3_imag <= _zz_73;
      end
      if(_zz_23)begin
        img_reg_array_21_3_imag <= _zz_73;
      end
      if(_zz_24)begin
        img_reg_array_22_3_imag <= _zz_73;
      end
      if(_zz_25)begin
        img_reg_array_23_3_imag <= _zz_73;
      end
      if(_zz_26)begin
        img_reg_array_24_3_imag <= _zz_73;
      end
      if(_zz_27)begin
        img_reg_array_25_3_imag <= _zz_73;
      end
      if(_zz_28)begin
        img_reg_array_26_3_imag <= _zz_73;
      end
      if(_zz_29)begin
        img_reg_array_27_3_imag <= _zz_73;
      end
      if(_zz_30)begin
        img_reg_array_28_3_imag <= _zz_73;
      end
      if(_zz_31)begin
        img_reg_array_29_3_imag <= _zz_73;
      end
      if(_zz_32)begin
        img_reg_array_30_3_imag <= _zz_73;
      end
      if(_zz_33)begin
        img_reg_array_31_3_imag <= _zz_73;
      end
      if(_zz_34)begin
        img_reg_array_32_3_imag <= _zz_73;
      end
      if(_zz_35)begin
        img_reg_array_33_3_imag <= _zz_73;
      end
      if(_zz_36)begin
        img_reg_array_34_3_imag <= _zz_73;
      end
      if(_zz_37)begin
        img_reg_array_35_3_imag <= _zz_73;
      end
      if(_zz_38)begin
        img_reg_array_36_3_imag <= _zz_73;
      end
      if(_zz_39)begin
        img_reg_array_37_3_imag <= _zz_73;
      end
      if(_zz_40)begin
        img_reg_array_38_3_imag <= _zz_73;
      end
      if(_zz_41)begin
        img_reg_array_39_3_imag <= _zz_73;
      end
      if(_zz_42)begin
        img_reg_array_40_3_imag <= _zz_73;
      end
      if(_zz_43)begin
        img_reg_array_41_3_imag <= _zz_73;
      end
      if(_zz_44)begin
        img_reg_array_42_3_imag <= _zz_73;
      end
      if(_zz_45)begin
        img_reg_array_43_3_imag <= _zz_73;
      end
      if(_zz_46)begin
        img_reg_array_44_3_imag <= _zz_73;
      end
      if(_zz_47)begin
        img_reg_array_45_3_imag <= _zz_73;
      end
      if(_zz_48)begin
        img_reg_array_46_3_imag <= _zz_73;
      end
      if(_zz_49)begin
        img_reg_array_47_3_imag <= _zz_73;
      end
      if(_zz_50)begin
        img_reg_array_48_3_imag <= _zz_73;
      end
      if(_zz_51)begin
        img_reg_array_49_3_imag <= _zz_73;
      end
      if(_zz_52)begin
        img_reg_array_50_3_imag <= _zz_73;
      end
      if(_zz_53)begin
        img_reg_array_51_3_imag <= _zz_73;
      end
      if(_zz_54)begin
        img_reg_array_52_3_imag <= _zz_73;
      end
      if(_zz_55)begin
        img_reg_array_53_3_imag <= _zz_73;
      end
      if(_zz_56)begin
        img_reg_array_54_3_imag <= _zz_73;
      end
      if(_zz_57)begin
        img_reg_array_55_3_imag <= _zz_73;
      end
      if(_zz_58)begin
        img_reg_array_56_3_imag <= _zz_73;
      end
      if(_zz_59)begin
        img_reg_array_57_3_imag <= _zz_73;
      end
      if(_zz_60)begin
        img_reg_array_58_3_imag <= _zz_73;
      end
      if(_zz_61)begin
        img_reg_array_59_3_imag <= _zz_73;
      end
      if(_zz_62)begin
        img_reg_array_60_3_imag <= _zz_73;
      end
      if(_zz_63)begin
        img_reg_array_61_3_imag <= _zz_73;
      end
      if(_zz_64)begin
        img_reg_array_62_3_imag <= _zz_73;
      end
      if(_zz_65)begin
        img_reg_array_63_3_imag <= _zz_73;
      end
      if(_zz_2)begin
        img_reg_array_0_4_real <= _zz_74;
      end
      if(_zz_3)begin
        img_reg_array_1_4_real <= _zz_74;
      end
      if(_zz_4)begin
        img_reg_array_2_4_real <= _zz_74;
      end
      if(_zz_5)begin
        img_reg_array_3_4_real <= _zz_74;
      end
      if(_zz_6)begin
        img_reg_array_4_4_real <= _zz_74;
      end
      if(_zz_7)begin
        img_reg_array_5_4_real <= _zz_74;
      end
      if(_zz_8)begin
        img_reg_array_6_4_real <= _zz_74;
      end
      if(_zz_9)begin
        img_reg_array_7_4_real <= _zz_74;
      end
      if(_zz_10)begin
        img_reg_array_8_4_real <= _zz_74;
      end
      if(_zz_11)begin
        img_reg_array_9_4_real <= _zz_74;
      end
      if(_zz_12)begin
        img_reg_array_10_4_real <= _zz_74;
      end
      if(_zz_13)begin
        img_reg_array_11_4_real <= _zz_74;
      end
      if(_zz_14)begin
        img_reg_array_12_4_real <= _zz_74;
      end
      if(_zz_15)begin
        img_reg_array_13_4_real <= _zz_74;
      end
      if(_zz_16)begin
        img_reg_array_14_4_real <= _zz_74;
      end
      if(_zz_17)begin
        img_reg_array_15_4_real <= _zz_74;
      end
      if(_zz_18)begin
        img_reg_array_16_4_real <= _zz_74;
      end
      if(_zz_19)begin
        img_reg_array_17_4_real <= _zz_74;
      end
      if(_zz_20)begin
        img_reg_array_18_4_real <= _zz_74;
      end
      if(_zz_21)begin
        img_reg_array_19_4_real <= _zz_74;
      end
      if(_zz_22)begin
        img_reg_array_20_4_real <= _zz_74;
      end
      if(_zz_23)begin
        img_reg_array_21_4_real <= _zz_74;
      end
      if(_zz_24)begin
        img_reg_array_22_4_real <= _zz_74;
      end
      if(_zz_25)begin
        img_reg_array_23_4_real <= _zz_74;
      end
      if(_zz_26)begin
        img_reg_array_24_4_real <= _zz_74;
      end
      if(_zz_27)begin
        img_reg_array_25_4_real <= _zz_74;
      end
      if(_zz_28)begin
        img_reg_array_26_4_real <= _zz_74;
      end
      if(_zz_29)begin
        img_reg_array_27_4_real <= _zz_74;
      end
      if(_zz_30)begin
        img_reg_array_28_4_real <= _zz_74;
      end
      if(_zz_31)begin
        img_reg_array_29_4_real <= _zz_74;
      end
      if(_zz_32)begin
        img_reg_array_30_4_real <= _zz_74;
      end
      if(_zz_33)begin
        img_reg_array_31_4_real <= _zz_74;
      end
      if(_zz_34)begin
        img_reg_array_32_4_real <= _zz_74;
      end
      if(_zz_35)begin
        img_reg_array_33_4_real <= _zz_74;
      end
      if(_zz_36)begin
        img_reg_array_34_4_real <= _zz_74;
      end
      if(_zz_37)begin
        img_reg_array_35_4_real <= _zz_74;
      end
      if(_zz_38)begin
        img_reg_array_36_4_real <= _zz_74;
      end
      if(_zz_39)begin
        img_reg_array_37_4_real <= _zz_74;
      end
      if(_zz_40)begin
        img_reg_array_38_4_real <= _zz_74;
      end
      if(_zz_41)begin
        img_reg_array_39_4_real <= _zz_74;
      end
      if(_zz_42)begin
        img_reg_array_40_4_real <= _zz_74;
      end
      if(_zz_43)begin
        img_reg_array_41_4_real <= _zz_74;
      end
      if(_zz_44)begin
        img_reg_array_42_4_real <= _zz_74;
      end
      if(_zz_45)begin
        img_reg_array_43_4_real <= _zz_74;
      end
      if(_zz_46)begin
        img_reg_array_44_4_real <= _zz_74;
      end
      if(_zz_47)begin
        img_reg_array_45_4_real <= _zz_74;
      end
      if(_zz_48)begin
        img_reg_array_46_4_real <= _zz_74;
      end
      if(_zz_49)begin
        img_reg_array_47_4_real <= _zz_74;
      end
      if(_zz_50)begin
        img_reg_array_48_4_real <= _zz_74;
      end
      if(_zz_51)begin
        img_reg_array_49_4_real <= _zz_74;
      end
      if(_zz_52)begin
        img_reg_array_50_4_real <= _zz_74;
      end
      if(_zz_53)begin
        img_reg_array_51_4_real <= _zz_74;
      end
      if(_zz_54)begin
        img_reg_array_52_4_real <= _zz_74;
      end
      if(_zz_55)begin
        img_reg_array_53_4_real <= _zz_74;
      end
      if(_zz_56)begin
        img_reg_array_54_4_real <= _zz_74;
      end
      if(_zz_57)begin
        img_reg_array_55_4_real <= _zz_74;
      end
      if(_zz_58)begin
        img_reg_array_56_4_real <= _zz_74;
      end
      if(_zz_59)begin
        img_reg_array_57_4_real <= _zz_74;
      end
      if(_zz_60)begin
        img_reg_array_58_4_real <= _zz_74;
      end
      if(_zz_61)begin
        img_reg_array_59_4_real <= _zz_74;
      end
      if(_zz_62)begin
        img_reg_array_60_4_real <= _zz_74;
      end
      if(_zz_63)begin
        img_reg_array_61_4_real <= _zz_74;
      end
      if(_zz_64)begin
        img_reg_array_62_4_real <= _zz_74;
      end
      if(_zz_65)begin
        img_reg_array_63_4_real <= _zz_74;
      end
      if(_zz_2)begin
        img_reg_array_0_4_imag <= _zz_75;
      end
      if(_zz_3)begin
        img_reg_array_1_4_imag <= _zz_75;
      end
      if(_zz_4)begin
        img_reg_array_2_4_imag <= _zz_75;
      end
      if(_zz_5)begin
        img_reg_array_3_4_imag <= _zz_75;
      end
      if(_zz_6)begin
        img_reg_array_4_4_imag <= _zz_75;
      end
      if(_zz_7)begin
        img_reg_array_5_4_imag <= _zz_75;
      end
      if(_zz_8)begin
        img_reg_array_6_4_imag <= _zz_75;
      end
      if(_zz_9)begin
        img_reg_array_7_4_imag <= _zz_75;
      end
      if(_zz_10)begin
        img_reg_array_8_4_imag <= _zz_75;
      end
      if(_zz_11)begin
        img_reg_array_9_4_imag <= _zz_75;
      end
      if(_zz_12)begin
        img_reg_array_10_4_imag <= _zz_75;
      end
      if(_zz_13)begin
        img_reg_array_11_4_imag <= _zz_75;
      end
      if(_zz_14)begin
        img_reg_array_12_4_imag <= _zz_75;
      end
      if(_zz_15)begin
        img_reg_array_13_4_imag <= _zz_75;
      end
      if(_zz_16)begin
        img_reg_array_14_4_imag <= _zz_75;
      end
      if(_zz_17)begin
        img_reg_array_15_4_imag <= _zz_75;
      end
      if(_zz_18)begin
        img_reg_array_16_4_imag <= _zz_75;
      end
      if(_zz_19)begin
        img_reg_array_17_4_imag <= _zz_75;
      end
      if(_zz_20)begin
        img_reg_array_18_4_imag <= _zz_75;
      end
      if(_zz_21)begin
        img_reg_array_19_4_imag <= _zz_75;
      end
      if(_zz_22)begin
        img_reg_array_20_4_imag <= _zz_75;
      end
      if(_zz_23)begin
        img_reg_array_21_4_imag <= _zz_75;
      end
      if(_zz_24)begin
        img_reg_array_22_4_imag <= _zz_75;
      end
      if(_zz_25)begin
        img_reg_array_23_4_imag <= _zz_75;
      end
      if(_zz_26)begin
        img_reg_array_24_4_imag <= _zz_75;
      end
      if(_zz_27)begin
        img_reg_array_25_4_imag <= _zz_75;
      end
      if(_zz_28)begin
        img_reg_array_26_4_imag <= _zz_75;
      end
      if(_zz_29)begin
        img_reg_array_27_4_imag <= _zz_75;
      end
      if(_zz_30)begin
        img_reg_array_28_4_imag <= _zz_75;
      end
      if(_zz_31)begin
        img_reg_array_29_4_imag <= _zz_75;
      end
      if(_zz_32)begin
        img_reg_array_30_4_imag <= _zz_75;
      end
      if(_zz_33)begin
        img_reg_array_31_4_imag <= _zz_75;
      end
      if(_zz_34)begin
        img_reg_array_32_4_imag <= _zz_75;
      end
      if(_zz_35)begin
        img_reg_array_33_4_imag <= _zz_75;
      end
      if(_zz_36)begin
        img_reg_array_34_4_imag <= _zz_75;
      end
      if(_zz_37)begin
        img_reg_array_35_4_imag <= _zz_75;
      end
      if(_zz_38)begin
        img_reg_array_36_4_imag <= _zz_75;
      end
      if(_zz_39)begin
        img_reg_array_37_4_imag <= _zz_75;
      end
      if(_zz_40)begin
        img_reg_array_38_4_imag <= _zz_75;
      end
      if(_zz_41)begin
        img_reg_array_39_4_imag <= _zz_75;
      end
      if(_zz_42)begin
        img_reg_array_40_4_imag <= _zz_75;
      end
      if(_zz_43)begin
        img_reg_array_41_4_imag <= _zz_75;
      end
      if(_zz_44)begin
        img_reg_array_42_4_imag <= _zz_75;
      end
      if(_zz_45)begin
        img_reg_array_43_4_imag <= _zz_75;
      end
      if(_zz_46)begin
        img_reg_array_44_4_imag <= _zz_75;
      end
      if(_zz_47)begin
        img_reg_array_45_4_imag <= _zz_75;
      end
      if(_zz_48)begin
        img_reg_array_46_4_imag <= _zz_75;
      end
      if(_zz_49)begin
        img_reg_array_47_4_imag <= _zz_75;
      end
      if(_zz_50)begin
        img_reg_array_48_4_imag <= _zz_75;
      end
      if(_zz_51)begin
        img_reg_array_49_4_imag <= _zz_75;
      end
      if(_zz_52)begin
        img_reg_array_50_4_imag <= _zz_75;
      end
      if(_zz_53)begin
        img_reg_array_51_4_imag <= _zz_75;
      end
      if(_zz_54)begin
        img_reg_array_52_4_imag <= _zz_75;
      end
      if(_zz_55)begin
        img_reg_array_53_4_imag <= _zz_75;
      end
      if(_zz_56)begin
        img_reg_array_54_4_imag <= _zz_75;
      end
      if(_zz_57)begin
        img_reg_array_55_4_imag <= _zz_75;
      end
      if(_zz_58)begin
        img_reg_array_56_4_imag <= _zz_75;
      end
      if(_zz_59)begin
        img_reg_array_57_4_imag <= _zz_75;
      end
      if(_zz_60)begin
        img_reg_array_58_4_imag <= _zz_75;
      end
      if(_zz_61)begin
        img_reg_array_59_4_imag <= _zz_75;
      end
      if(_zz_62)begin
        img_reg_array_60_4_imag <= _zz_75;
      end
      if(_zz_63)begin
        img_reg_array_61_4_imag <= _zz_75;
      end
      if(_zz_64)begin
        img_reg_array_62_4_imag <= _zz_75;
      end
      if(_zz_65)begin
        img_reg_array_63_4_imag <= _zz_75;
      end
      if(_zz_2)begin
        img_reg_array_0_5_real <= _zz_76;
      end
      if(_zz_3)begin
        img_reg_array_1_5_real <= _zz_76;
      end
      if(_zz_4)begin
        img_reg_array_2_5_real <= _zz_76;
      end
      if(_zz_5)begin
        img_reg_array_3_5_real <= _zz_76;
      end
      if(_zz_6)begin
        img_reg_array_4_5_real <= _zz_76;
      end
      if(_zz_7)begin
        img_reg_array_5_5_real <= _zz_76;
      end
      if(_zz_8)begin
        img_reg_array_6_5_real <= _zz_76;
      end
      if(_zz_9)begin
        img_reg_array_7_5_real <= _zz_76;
      end
      if(_zz_10)begin
        img_reg_array_8_5_real <= _zz_76;
      end
      if(_zz_11)begin
        img_reg_array_9_5_real <= _zz_76;
      end
      if(_zz_12)begin
        img_reg_array_10_5_real <= _zz_76;
      end
      if(_zz_13)begin
        img_reg_array_11_5_real <= _zz_76;
      end
      if(_zz_14)begin
        img_reg_array_12_5_real <= _zz_76;
      end
      if(_zz_15)begin
        img_reg_array_13_5_real <= _zz_76;
      end
      if(_zz_16)begin
        img_reg_array_14_5_real <= _zz_76;
      end
      if(_zz_17)begin
        img_reg_array_15_5_real <= _zz_76;
      end
      if(_zz_18)begin
        img_reg_array_16_5_real <= _zz_76;
      end
      if(_zz_19)begin
        img_reg_array_17_5_real <= _zz_76;
      end
      if(_zz_20)begin
        img_reg_array_18_5_real <= _zz_76;
      end
      if(_zz_21)begin
        img_reg_array_19_5_real <= _zz_76;
      end
      if(_zz_22)begin
        img_reg_array_20_5_real <= _zz_76;
      end
      if(_zz_23)begin
        img_reg_array_21_5_real <= _zz_76;
      end
      if(_zz_24)begin
        img_reg_array_22_5_real <= _zz_76;
      end
      if(_zz_25)begin
        img_reg_array_23_5_real <= _zz_76;
      end
      if(_zz_26)begin
        img_reg_array_24_5_real <= _zz_76;
      end
      if(_zz_27)begin
        img_reg_array_25_5_real <= _zz_76;
      end
      if(_zz_28)begin
        img_reg_array_26_5_real <= _zz_76;
      end
      if(_zz_29)begin
        img_reg_array_27_5_real <= _zz_76;
      end
      if(_zz_30)begin
        img_reg_array_28_5_real <= _zz_76;
      end
      if(_zz_31)begin
        img_reg_array_29_5_real <= _zz_76;
      end
      if(_zz_32)begin
        img_reg_array_30_5_real <= _zz_76;
      end
      if(_zz_33)begin
        img_reg_array_31_5_real <= _zz_76;
      end
      if(_zz_34)begin
        img_reg_array_32_5_real <= _zz_76;
      end
      if(_zz_35)begin
        img_reg_array_33_5_real <= _zz_76;
      end
      if(_zz_36)begin
        img_reg_array_34_5_real <= _zz_76;
      end
      if(_zz_37)begin
        img_reg_array_35_5_real <= _zz_76;
      end
      if(_zz_38)begin
        img_reg_array_36_5_real <= _zz_76;
      end
      if(_zz_39)begin
        img_reg_array_37_5_real <= _zz_76;
      end
      if(_zz_40)begin
        img_reg_array_38_5_real <= _zz_76;
      end
      if(_zz_41)begin
        img_reg_array_39_5_real <= _zz_76;
      end
      if(_zz_42)begin
        img_reg_array_40_5_real <= _zz_76;
      end
      if(_zz_43)begin
        img_reg_array_41_5_real <= _zz_76;
      end
      if(_zz_44)begin
        img_reg_array_42_5_real <= _zz_76;
      end
      if(_zz_45)begin
        img_reg_array_43_5_real <= _zz_76;
      end
      if(_zz_46)begin
        img_reg_array_44_5_real <= _zz_76;
      end
      if(_zz_47)begin
        img_reg_array_45_5_real <= _zz_76;
      end
      if(_zz_48)begin
        img_reg_array_46_5_real <= _zz_76;
      end
      if(_zz_49)begin
        img_reg_array_47_5_real <= _zz_76;
      end
      if(_zz_50)begin
        img_reg_array_48_5_real <= _zz_76;
      end
      if(_zz_51)begin
        img_reg_array_49_5_real <= _zz_76;
      end
      if(_zz_52)begin
        img_reg_array_50_5_real <= _zz_76;
      end
      if(_zz_53)begin
        img_reg_array_51_5_real <= _zz_76;
      end
      if(_zz_54)begin
        img_reg_array_52_5_real <= _zz_76;
      end
      if(_zz_55)begin
        img_reg_array_53_5_real <= _zz_76;
      end
      if(_zz_56)begin
        img_reg_array_54_5_real <= _zz_76;
      end
      if(_zz_57)begin
        img_reg_array_55_5_real <= _zz_76;
      end
      if(_zz_58)begin
        img_reg_array_56_5_real <= _zz_76;
      end
      if(_zz_59)begin
        img_reg_array_57_5_real <= _zz_76;
      end
      if(_zz_60)begin
        img_reg_array_58_5_real <= _zz_76;
      end
      if(_zz_61)begin
        img_reg_array_59_5_real <= _zz_76;
      end
      if(_zz_62)begin
        img_reg_array_60_5_real <= _zz_76;
      end
      if(_zz_63)begin
        img_reg_array_61_5_real <= _zz_76;
      end
      if(_zz_64)begin
        img_reg_array_62_5_real <= _zz_76;
      end
      if(_zz_65)begin
        img_reg_array_63_5_real <= _zz_76;
      end
      if(_zz_2)begin
        img_reg_array_0_5_imag <= _zz_77;
      end
      if(_zz_3)begin
        img_reg_array_1_5_imag <= _zz_77;
      end
      if(_zz_4)begin
        img_reg_array_2_5_imag <= _zz_77;
      end
      if(_zz_5)begin
        img_reg_array_3_5_imag <= _zz_77;
      end
      if(_zz_6)begin
        img_reg_array_4_5_imag <= _zz_77;
      end
      if(_zz_7)begin
        img_reg_array_5_5_imag <= _zz_77;
      end
      if(_zz_8)begin
        img_reg_array_6_5_imag <= _zz_77;
      end
      if(_zz_9)begin
        img_reg_array_7_5_imag <= _zz_77;
      end
      if(_zz_10)begin
        img_reg_array_8_5_imag <= _zz_77;
      end
      if(_zz_11)begin
        img_reg_array_9_5_imag <= _zz_77;
      end
      if(_zz_12)begin
        img_reg_array_10_5_imag <= _zz_77;
      end
      if(_zz_13)begin
        img_reg_array_11_5_imag <= _zz_77;
      end
      if(_zz_14)begin
        img_reg_array_12_5_imag <= _zz_77;
      end
      if(_zz_15)begin
        img_reg_array_13_5_imag <= _zz_77;
      end
      if(_zz_16)begin
        img_reg_array_14_5_imag <= _zz_77;
      end
      if(_zz_17)begin
        img_reg_array_15_5_imag <= _zz_77;
      end
      if(_zz_18)begin
        img_reg_array_16_5_imag <= _zz_77;
      end
      if(_zz_19)begin
        img_reg_array_17_5_imag <= _zz_77;
      end
      if(_zz_20)begin
        img_reg_array_18_5_imag <= _zz_77;
      end
      if(_zz_21)begin
        img_reg_array_19_5_imag <= _zz_77;
      end
      if(_zz_22)begin
        img_reg_array_20_5_imag <= _zz_77;
      end
      if(_zz_23)begin
        img_reg_array_21_5_imag <= _zz_77;
      end
      if(_zz_24)begin
        img_reg_array_22_5_imag <= _zz_77;
      end
      if(_zz_25)begin
        img_reg_array_23_5_imag <= _zz_77;
      end
      if(_zz_26)begin
        img_reg_array_24_5_imag <= _zz_77;
      end
      if(_zz_27)begin
        img_reg_array_25_5_imag <= _zz_77;
      end
      if(_zz_28)begin
        img_reg_array_26_5_imag <= _zz_77;
      end
      if(_zz_29)begin
        img_reg_array_27_5_imag <= _zz_77;
      end
      if(_zz_30)begin
        img_reg_array_28_5_imag <= _zz_77;
      end
      if(_zz_31)begin
        img_reg_array_29_5_imag <= _zz_77;
      end
      if(_zz_32)begin
        img_reg_array_30_5_imag <= _zz_77;
      end
      if(_zz_33)begin
        img_reg_array_31_5_imag <= _zz_77;
      end
      if(_zz_34)begin
        img_reg_array_32_5_imag <= _zz_77;
      end
      if(_zz_35)begin
        img_reg_array_33_5_imag <= _zz_77;
      end
      if(_zz_36)begin
        img_reg_array_34_5_imag <= _zz_77;
      end
      if(_zz_37)begin
        img_reg_array_35_5_imag <= _zz_77;
      end
      if(_zz_38)begin
        img_reg_array_36_5_imag <= _zz_77;
      end
      if(_zz_39)begin
        img_reg_array_37_5_imag <= _zz_77;
      end
      if(_zz_40)begin
        img_reg_array_38_5_imag <= _zz_77;
      end
      if(_zz_41)begin
        img_reg_array_39_5_imag <= _zz_77;
      end
      if(_zz_42)begin
        img_reg_array_40_5_imag <= _zz_77;
      end
      if(_zz_43)begin
        img_reg_array_41_5_imag <= _zz_77;
      end
      if(_zz_44)begin
        img_reg_array_42_5_imag <= _zz_77;
      end
      if(_zz_45)begin
        img_reg_array_43_5_imag <= _zz_77;
      end
      if(_zz_46)begin
        img_reg_array_44_5_imag <= _zz_77;
      end
      if(_zz_47)begin
        img_reg_array_45_5_imag <= _zz_77;
      end
      if(_zz_48)begin
        img_reg_array_46_5_imag <= _zz_77;
      end
      if(_zz_49)begin
        img_reg_array_47_5_imag <= _zz_77;
      end
      if(_zz_50)begin
        img_reg_array_48_5_imag <= _zz_77;
      end
      if(_zz_51)begin
        img_reg_array_49_5_imag <= _zz_77;
      end
      if(_zz_52)begin
        img_reg_array_50_5_imag <= _zz_77;
      end
      if(_zz_53)begin
        img_reg_array_51_5_imag <= _zz_77;
      end
      if(_zz_54)begin
        img_reg_array_52_5_imag <= _zz_77;
      end
      if(_zz_55)begin
        img_reg_array_53_5_imag <= _zz_77;
      end
      if(_zz_56)begin
        img_reg_array_54_5_imag <= _zz_77;
      end
      if(_zz_57)begin
        img_reg_array_55_5_imag <= _zz_77;
      end
      if(_zz_58)begin
        img_reg_array_56_5_imag <= _zz_77;
      end
      if(_zz_59)begin
        img_reg_array_57_5_imag <= _zz_77;
      end
      if(_zz_60)begin
        img_reg_array_58_5_imag <= _zz_77;
      end
      if(_zz_61)begin
        img_reg_array_59_5_imag <= _zz_77;
      end
      if(_zz_62)begin
        img_reg_array_60_5_imag <= _zz_77;
      end
      if(_zz_63)begin
        img_reg_array_61_5_imag <= _zz_77;
      end
      if(_zz_64)begin
        img_reg_array_62_5_imag <= _zz_77;
      end
      if(_zz_65)begin
        img_reg_array_63_5_imag <= _zz_77;
      end
      if(_zz_2)begin
        img_reg_array_0_6_real <= _zz_78;
      end
      if(_zz_3)begin
        img_reg_array_1_6_real <= _zz_78;
      end
      if(_zz_4)begin
        img_reg_array_2_6_real <= _zz_78;
      end
      if(_zz_5)begin
        img_reg_array_3_6_real <= _zz_78;
      end
      if(_zz_6)begin
        img_reg_array_4_6_real <= _zz_78;
      end
      if(_zz_7)begin
        img_reg_array_5_6_real <= _zz_78;
      end
      if(_zz_8)begin
        img_reg_array_6_6_real <= _zz_78;
      end
      if(_zz_9)begin
        img_reg_array_7_6_real <= _zz_78;
      end
      if(_zz_10)begin
        img_reg_array_8_6_real <= _zz_78;
      end
      if(_zz_11)begin
        img_reg_array_9_6_real <= _zz_78;
      end
      if(_zz_12)begin
        img_reg_array_10_6_real <= _zz_78;
      end
      if(_zz_13)begin
        img_reg_array_11_6_real <= _zz_78;
      end
      if(_zz_14)begin
        img_reg_array_12_6_real <= _zz_78;
      end
      if(_zz_15)begin
        img_reg_array_13_6_real <= _zz_78;
      end
      if(_zz_16)begin
        img_reg_array_14_6_real <= _zz_78;
      end
      if(_zz_17)begin
        img_reg_array_15_6_real <= _zz_78;
      end
      if(_zz_18)begin
        img_reg_array_16_6_real <= _zz_78;
      end
      if(_zz_19)begin
        img_reg_array_17_6_real <= _zz_78;
      end
      if(_zz_20)begin
        img_reg_array_18_6_real <= _zz_78;
      end
      if(_zz_21)begin
        img_reg_array_19_6_real <= _zz_78;
      end
      if(_zz_22)begin
        img_reg_array_20_6_real <= _zz_78;
      end
      if(_zz_23)begin
        img_reg_array_21_6_real <= _zz_78;
      end
      if(_zz_24)begin
        img_reg_array_22_6_real <= _zz_78;
      end
      if(_zz_25)begin
        img_reg_array_23_6_real <= _zz_78;
      end
      if(_zz_26)begin
        img_reg_array_24_6_real <= _zz_78;
      end
      if(_zz_27)begin
        img_reg_array_25_6_real <= _zz_78;
      end
      if(_zz_28)begin
        img_reg_array_26_6_real <= _zz_78;
      end
      if(_zz_29)begin
        img_reg_array_27_6_real <= _zz_78;
      end
      if(_zz_30)begin
        img_reg_array_28_6_real <= _zz_78;
      end
      if(_zz_31)begin
        img_reg_array_29_6_real <= _zz_78;
      end
      if(_zz_32)begin
        img_reg_array_30_6_real <= _zz_78;
      end
      if(_zz_33)begin
        img_reg_array_31_6_real <= _zz_78;
      end
      if(_zz_34)begin
        img_reg_array_32_6_real <= _zz_78;
      end
      if(_zz_35)begin
        img_reg_array_33_6_real <= _zz_78;
      end
      if(_zz_36)begin
        img_reg_array_34_6_real <= _zz_78;
      end
      if(_zz_37)begin
        img_reg_array_35_6_real <= _zz_78;
      end
      if(_zz_38)begin
        img_reg_array_36_6_real <= _zz_78;
      end
      if(_zz_39)begin
        img_reg_array_37_6_real <= _zz_78;
      end
      if(_zz_40)begin
        img_reg_array_38_6_real <= _zz_78;
      end
      if(_zz_41)begin
        img_reg_array_39_6_real <= _zz_78;
      end
      if(_zz_42)begin
        img_reg_array_40_6_real <= _zz_78;
      end
      if(_zz_43)begin
        img_reg_array_41_6_real <= _zz_78;
      end
      if(_zz_44)begin
        img_reg_array_42_6_real <= _zz_78;
      end
      if(_zz_45)begin
        img_reg_array_43_6_real <= _zz_78;
      end
      if(_zz_46)begin
        img_reg_array_44_6_real <= _zz_78;
      end
      if(_zz_47)begin
        img_reg_array_45_6_real <= _zz_78;
      end
      if(_zz_48)begin
        img_reg_array_46_6_real <= _zz_78;
      end
      if(_zz_49)begin
        img_reg_array_47_6_real <= _zz_78;
      end
      if(_zz_50)begin
        img_reg_array_48_6_real <= _zz_78;
      end
      if(_zz_51)begin
        img_reg_array_49_6_real <= _zz_78;
      end
      if(_zz_52)begin
        img_reg_array_50_6_real <= _zz_78;
      end
      if(_zz_53)begin
        img_reg_array_51_6_real <= _zz_78;
      end
      if(_zz_54)begin
        img_reg_array_52_6_real <= _zz_78;
      end
      if(_zz_55)begin
        img_reg_array_53_6_real <= _zz_78;
      end
      if(_zz_56)begin
        img_reg_array_54_6_real <= _zz_78;
      end
      if(_zz_57)begin
        img_reg_array_55_6_real <= _zz_78;
      end
      if(_zz_58)begin
        img_reg_array_56_6_real <= _zz_78;
      end
      if(_zz_59)begin
        img_reg_array_57_6_real <= _zz_78;
      end
      if(_zz_60)begin
        img_reg_array_58_6_real <= _zz_78;
      end
      if(_zz_61)begin
        img_reg_array_59_6_real <= _zz_78;
      end
      if(_zz_62)begin
        img_reg_array_60_6_real <= _zz_78;
      end
      if(_zz_63)begin
        img_reg_array_61_6_real <= _zz_78;
      end
      if(_zz_64)begin
        img_reg_array_62_6_real <= _zz_78;
      end
      if(_zz_65)begin
        img_reg_array_63_6_real <= _zz_78;
      end
      if(_zz_2)begin
        img_reg_array_0_6_imag <= _zz_79;
      end
      if(_zz_3)begin
        img_reg_array_1_6_imag <= _zz_79;
      end
      if(_zz_4)begin
        img_reg_array_2_6_imag <= _zz_79;
      end
      if(_zz_5)begin
        img_reg_array_3_6_imag <= _zz_79;
      end
      if(_zz_6)begin
        img_reg_array_4_6_imag <= _zz_79;
      end
      if(_zz_7)begin
        img_reg_array_5_6_imag <= _zz_79;
      end
      if(_zz_8)begin
        img_reg_array_6_6_imag <= _zz_79;
      end
      if(_zz_9)begin
        img_reg_array_7_6_imag <= _zz_79;
      end
      if(_zz_10)begin
        img_reg_array_8_6_imag <= _zz_79;
      end
      if(_zz_11)begin
        img_reg_array_9_6_imag <= _zz_79;
      end
      if(_zz_12)begin
        img_reg_array_10_6_imag <= _zz_79;
      end
      if(_zz_13)begin
        img_reg_array_11_6_imag <= _zz_79;
      end
      if(_zz_14)begin
        img_reg_array_12_6_imag <= _zz_79;
      end
      if(_zz_15)begin
        img_reg_array_13_6_imag <= _zz_79;
      end
      if(_zz_16)begin
        img_reg_array_14_6_imag <= _zz_79;
      end
      if(_zz_17)begin
        img_reg_array_15_6_imag <= _zz_79;
      end
      if(_zz_18)begin
        img_reg_array_16_6_imag <= _zz_79;
      end
      if(_zz_19)begin
        img_reg_array_17_6_imag <= _zz_79;
      end
      if(_zz_20)begin
        img_reg_array_18_6_imag <= _zz_79;
      end
      if(_zz_21)begin
        img_reg_array_19_6_imag <= _zz_79;
      end
      if(_zz_22)begin
        img_reg_array_20_6_imag <= _zz_79;
      end
      if(_zz_23)begin
        img_reg_array_21_6_imag <= _zz_79;
      end
      if(_zz_24)begin
        img_reg_array_22_6_imag <= _zz_79;
      end
      if(_zz_25)begin
        img_reg_array_23_6_imag <= _zz_79;
      end
      if(_zz_26)begin
        img_reg_array_24_6_imag <= _zz_79;
      end
      if(_zz_27)begin
        img_reg_array_25_6_imag <= _zz_79;
      end
      if(_zz_28)begin
        img_reg_array_26_6_imag <= _zz_79;
      end
      if(_zz_29)begin
        img_reg_array_27_6_imag <= _zz_79;
      end
      if(_zz_30)begin
        img_reg_array_28_6_imag <= _zz_79;
      end
      if(_zz_31)begin
        img_reg_array_29_6_imag <= _zz_79;
      end
      if(_zz_32)begin
        img_reg_array_30_6_imag <= _zz_79;
      end
      if(_zz_33)begin
        img_reg_array_31_6_imag <= _zz_79;
      end
      if(_zz_34)begin
        img_reg_array_32_6_imag <= _zz_79;
      end
      if(_zz_35)begin
        img_reg_array_33_6_imag <= _zz_79;
      end
      if(_zz_36)begin
        img_reg_array_34_6_imag <= _zz_79;
      end
      if(_zz_37)begin
        img_reg_array_35_6_imag <= _zz_79;
      end
      if(_zz_38)begin
        img_reg_array_36_6_imag <= _zz_79;
      end
      if(_zz_39)begin
        img_reg_array_37_6_imag <= _zz_79;
      end
      if(_zz_40)begin
        img_reg_array_38_6_imag <= _zz_79;
      end
      if(_zz_41)begin
        img_reg_array_39_6_imag <= _zz_79;
      end
      if(_zz_42)begin
        img_reg_array_40_6_imag <= _zz_79;
      end
      if(_zz_43)begin
        img_reg_array_41_6_imag <= _zz_79;
      end
      if(_zz_44)begin
        img_reg_array_42_6_imag <= _zz_79;
      end
      if(_zz_45)begin
        img_reg_array_43_6_imag <= _zz_79;
      end
      if(_zz_46)begin
        img_reg_array_44_6_imag <= _zz_79;
      end
      if(_zz_47)begin
        img_reg_array_45_6_imag <= _zz_79;
      end
      if(_zz_48)begin
        img_reg_array_46_6_imag <= _zz_79;
      end
      if(_zz_49)begin
        img_reg_array_47_6_imag <= _zz_79;
      end
      if(_zz_50)begin
        img_reg_array_48_6_imag <= _zz_79;
      end
      if(_zz_51)begin
        img_reg_array_49_6_imag <= _zz_79;
      end
      if(_zz_52)begin
        img_reg_array_50_6_imag <= _zz_79;
      end
      if(_zz_53)begin
        img_reg_array_51_6_imag <= _zz_79;
      end
      if(_zz_54)begin
        img_reg_array_52_6_imag <= _zz_79;
      end
      if(_zz_55)begin
        img_reg_array_53_6_imag <= _zz_79;
      end
      if(_zz_56)begin
        img_reg_array_54_6_imag <= _zz_79;
      end
      if(_zz_57)begin
        img_reg_array_55_6_imag <= _zz_79;
      end
      if(_zz_58)begin
        img_reg_array_56_6_imag <= _zz_79;
      end
      if(_zz_59)begin
        img_reg_array_57_6_imag <= _zz_79;
      end
      if(_zz_60)begin
        img_reg_array_58_6_imag <= _zz_79;
      end
      if(_zz_61)begin
        img_reg_array_59_6_imag <= _zz_79;
      end
      if(_zz_62)begin
        img_reg_array_60_6_imag <= _zz_79;
      end
      if(_zz_63)begin
        img_reg_array_61_6_imag <= _zz_79;
      end
      if(_zz_64)begin
        img_reg_array_62_6_imag <= _zz_79;
      end
      if(_zz_65)begin
        img_reg_array_63_6_imag <= _zz_79;
      end
      if(_zz_2)begin
        img_reg_array_0_7_real <= _zz_80;
      end
      if(_zz_3)begin
        img_reg_array_1_7_real <= _zz_80;
      end
      if(_zz_4)begin
        img_reg_array_2_7_real <= _zz_80;
      end
      if(_zz_5)begin
        img_reg_array_3_7_real <= _zz_80;
      end
      if(_zz_6)begin
        img_reg_array_4_7_real <= _zz_80;
      end
      if(_zz_7)begin
        img_reg_array_5_7_real <= _zz_80;
      end
      if(_zz_8)begin
        img_reg_array_6_7_real <= _zz_80;
      end
      if(_zz_9)begin
        img_reg_array_7_7_real <= _zz_80;
      end
      if(_zz_10)begin
        img_reg_array_8_7_real <= _zz_80;
      end
      if(_zz_11)begin
        img_reg_array_9_7_real <= _zz_80;
      end
      if(_zz_12)begin
        img_reg_array_10_7_real <= _zz_80;
      end
      if(_zz_13)begin
        img_reg_array_11_7_real <= _zz_80;
      end
      if(_zz_14)begin
        img_reg_array_12_7_real <= _zz_80;
      end
      if(_zz_15)begin
        img_reg_array_13_7_real <= _zz_80;
      end
      if(_zz_16)begin
        img_reg_array_14_7_real <= _zz_80;
      end
      if(_zz_17)begin
        img_reg_array_15_7_real <= _zz_80;
      end
      if(_zz_18)begin
        img_reg_array_16_7_real <= _zz_80;
      end
      if(_zz_19)begin
        img_reg_array_17_7_real <= _zz_80;
      end
      if(_zz_20)begin
        img_reg_array_18_7_real <= _zz_80;
      end
      if(_zz_21)begin
        img_reg_array_19_7_real <= _zz_80;
      end
      if(_zz_22)begin
        img_reg_array_20_7_real <= _zz_80;
      end
      if(_zz_23)begin
        img_reg_array_21_7_real <= _zz_80;
      end
      if(_zz_24)begin
        img_reg_array_22_7_real <= _zz_80;
      end
      if(_zz_25)begin
        img_reg_array_23_7_real <= _zz_80;
      end
      if(_zz_26)begin
        img_reg_array_24_7_real <= _zz_80;
      end
      if(_zz_27)begin
        img_reg_array_25_7_real <= _zz_80;
      end
      if(_zz_28)begin
        img_reg_array_26_7_real <= _zz_80;
      end
      if(_zz_29)begin
        img_reg_array_27_7_real <= _zz_80;
      end
      if(_zz_30)begin
        img_reg_array_28_7_real <= _zz_80;
      end
      if(_zz_31)begin
        img_reg_array_29_7_real <= _zz_80;
      end
      if(_zz_32)begin
        img_reg_array_30_7_real <= _zz_80;
      end
      if(_zz_33)begin
        img_reg_array_31_7_real <= _zz_80;
      end
      if(_zz_34)begin
        img_reg_array_32_7_real <= _zz_80;
      end
      if(_zz_35)begin
        img_reg_array_33_7_real <= _zz_80;
      end
      if(_zz_36)begin
        img_reg_array_34_7_real <= _zz_80;
      end
      if(_zz_37)begin
        img_reg_array_35_7_real <= _zz_80;
      end
      if(_zz_38)begin
        img_reg_array_36_7_real <= _zz_80;
      end
      if(_zz_39)begin
        img_reg_array_37_7_real <= _zz_80;
      end
      if(_zz_40)begin
        img_reg_array_38_7_real <= _zz_80;
      end
      if(_zz_41)begin
        img_reg_array_39_7_real <= _zz_80;
      end
      if(_zz_42)begin
        img_reg_array_40_7_real <= _zz_80;
      end
      if(_zz_43)begin
        img_reg_array_41_7_real <= _zz_80;
      end
      if(_zz_44)begin
        img_reg_array_42_7_real <= _zz_80;
      end
      if(_zz_45)begin
        img_reg_array_43_7_real <= _zz_80;
      end
      if(_zz_46)begin
        img_reg_array_44_7_real <= _zz_80;
      end
      if(_zz_47)begin
        img_reg_array_45_7_real <= _zz_80;
      end
      if(_zz_48)begin
        img_reg_array_46_7_real <= _zz_80;
      end
      if(_zz_49)begin
        img_reg_array_47_7_real <= _zz_80;
      end
      if(_zz_50)begin
        img_reg_array_48_7_real <= _zz_80;
      end
      if(_zz_51)begin
        img_reg_array_49_7_real <= _zz_80;
      end
      if(_zz_52)begin
        img_reg_array_50_7_real <= _zz_80;
      end
      if(_zz_53)begin
        img_reg_array_51_7_real <= _zz_80;
      end
      if(_zz_54)begin
        img_reg_array_52_7_real <= _zz_80;
      end
      if(_zz_55)begin
        img_reg_array_53_7_real <= _zz_80;
      end
      if(_zz_56)begin
        img_reg_array_54_7_real <= _zz_80;
      end
      if(_zz_57)begin
        img_reg_array_55_7_real <= _zz_80;
      end
      if(_zz_58)begin
        img_reg_array_56_7_real <= _zz_80;
      end
      if(_zz_59)begin
        img_reg_array_57_7_real <= _zz_80;
      end
      if(_zz_60)begin
        img_reg_array_58_7_real <= _zz_80;
      end
      if(_zz_61)begin
        img_reg_array_59_7_real <= _zz_80;
      end
      if(_zz_62)begin
        img_reg_array_60_7_real <= _zz_80;
      end
      if(_zz_63)begin
        img_reg_array_61_7_real <= _zz_80;
      end
      if(_zz_64)begin
        img_reg_array_62_7_real <= _zz_80;
      end
      if(_zz_65)begin
        img_reg_array_63_7_real <= _zz_80;
      end
      if(_zz_2)begin
        img_reg_array_0_7_imag <= _zz_81;
      end
      if(_zz_3)begin
        img_reg_array_1_7_imag <= _zz_81;
      end
      if(_zz_4)begin
        img_reg_array_2_7_imag <= _zz_81;
      end
      if(_zz_5)begin
        img_reg_array_3_7_imag <= _zz_81;
      end
      if(_zz_6)begin
        img_reg_array_4_7_imag <= _zz_81;
      end
      if(_zz_7)begin
        img_reg_array_5_7_imag <= _zz_81;
      end
      if(_zz_8)begin
        img_reg_array_6_7_imag <= _zz_81;
      end
      if(_zz_9)begin
        img_reg_array_7_7_imag <= _zz_81;
      end
      if(_zz_10)begin
        img_reg_array_8_7_imag <= _zz_81;
      end
      if(_zz_11)begin
        img_reg_array_9_7_imag <= _zz_81;
      end
      if(_zz_12)begin
        img_reg_array_10_7_imag <= _zz_81;
      end
      if(_zz_13)begin
        img_reg_array_11_7_imag <= _zz_81;
      end
      if(_zz_14)begin
        img_reg_array_12_7_imag <= _zz_81;
      end
      if(_zz_15)begin
        img_reg_array_13_7_imag <= _zz_81;
      end
      if(_zz_16)begin
        img_reg_array_14_7_imag <= _zz_81;
      end
      if(_zz_17)begin
        img_reg_array_15_7_imag <= _zz_81;
      end
      if(_zz_18)begin
        img_reg_array_16_7_imag <= _zz_81;
      end
      if(_zz_19)begin
        img_reg_array_17_7_imag <= _zz_81;
      end
      if(_zz_20)begin
        img_reg_array_18_7_imag <= _zz_81;
      end
      if(_zz_21)begin
        img_reg_array_19_7_imag <= _zz_81;
      end
      if(_zz_22)begin
        img_reg_array_20_7_imag <= _zz_81;
      end
      if(_zz_23)begin
        img_reg_array_21_7_imag <= _zz_81;
      end
      if(_zz_24)begin
        img_reg_array_22_7_imag <= _zz_81;
      end
      if(_zz_25)begin
        img_reg_array_23_7_imag <= _zz_81;
      end
      if(_zz_26)begin
        img_reg_array_24_7_imag <= _zz_81;
      end
      if(_zz_27)begin
        img_reg_array_25_7_imag <= _zz_81;
      end
      if(_zz_28)begin
        img_reg_array_26_7_imag <= _zz_81;
      end
      if(_zz_29)begin
        img_reg_array_27_7_imag <= _zz_81;
      end
      if(_zz_30)begin
        img_reg_array_28_7_imag <= _zz_81;
      end
      if(_zz_31)begin
        img_reg_array_29_7_imag <= _zz_81;
      end
      if(_zz_32)begin
        img_reg_array_30_7_imag <= _zz_81;
      end
      if(_zz_33)begin
        img_reg_array_31_7_imag <= _zz_81;
      end
      if(_zz_34)begin
        img_reg_array_32_7_imag <= _zz_81;
      end
      if(_zz_35)begin
        img_reg_array_33_7_imag <= _zz_81;
      end
      if(_zz_36)begin
        img_reg_array_34_7_imag <= _zz_81;
      end
      if(_zz_37)begin
        img_reg_array_35_7_imag <= _zz_81;
      end
      if(_zz_38)begin
        img_reg_array_36_7_imag <= _zz_81;
      end
      if(_zz_39)begin
        img_reg_array_37_7_imag <= _zz_81;
      end
      if(_zz_40)begin
        img_reg_array_38_7_imag <= _zz_81;
      end
      if(_zz_41)begin
        img_reg_array_39_7_imag <= _zz_81;
      end
      if(_zz_42)begin
        img_reg_array_40_7_imag <= _zz_81;
      end
      if(_zz_43)begin
        img_reg_array_41_7_imag <= _zz_81;
      end
      if(_zz_44)begin
        img_reg_array_42_7_imag <= _zz_81;
      end
      if(_zz_45)begin
        img_reg_array_43_7_imag <= _zz_81;
      end
      if(_zz_46)begin
        img_reg_array_44_7_imag <= _zz_81;
      end
      if(_zz_47)begin
        img_reg_array_45_7_imag <= _zz_81;
      end
      if(_zz_48)begin
        img_reg_array_46_7_imag <= _zz_81;
      end
      if(_zz_49)begin
        img_reg_array_47_7_imag <= _zz_81;
      end
      if(_zz_50)begin
        img_reg_array_48_7_imag <= _zz_81;
      end
      if(_zz_51)begin
        img_reg_array_49_7_imag <= _zz_81;
      end
      if(_zz_52)begin
        img_reg_array_50_7_imag <= _zz_81;
      end
      if(_zz_53)begin
        img_reg_array_51_7_imag <= _zz_81;
      end
      if(_zz_54)begin
        img_reg_array_52_7_imag <= _zz_81;
      end
      if(_zz_55)begin
        img_reg_array_53_7_imag <= _zz_81;
      end
      if(_zz_56)begin
        img_reg_array_54_7_imag <= _zz_81;
      end
      if(_zz_57)begin
        img_reg_array_55_7_imag <= _zz_81;
      end
      if(_zz_58)begin
        img_reg_array_56_7_imag <= _zz_81;
      end
      if(_zz_59)begin
        img_reg_array_57_7_imag <= _zz_81;
      end
      if(_zz_60)begin
        img_reg_array_58_7_imag <= _zz_81;
      end
      if(_zz_61)begin
        img_reg_array_59_7_imag <= _zz_81;
      end
      if(_zz_62)begin
        img_reg_array_60_7_imag <= _zz_81;
      end
      if(_zz_63)begin
        img_reg_array_61_7_imag <= _zz_81;
      end
      if(_zz_64)begin
        img_reg_array_62_7_imag <= _zz_81;
      end
      if(_zz_65)begin
        img_reg_array_63_7_imag <= _zz_81;
      end
      if(_zz_2)begin
        img_reg_array_0_8_real <= _zz_82;
      end
      if(_zz_3)begin
        img_reg_array_1_8_real <= _zz_82;
      end
      if(_zz_4)begin
        img_reg_array_2_8_real <= _zz_82;
      end
      if(_zz_5)begin
        img_reg_array_3_8_real <= _zz_82;
      end
      if(_zz_6)begin
        img_reg_array_4_8_real <= _zz_82;
      end
      if(_zz_7)begin
        img_reg_array_5_8_real <= _zz_82;
      end
      if(_zz_8)begin
        img_reg_array_6_8_real <= _zz_82;
      end
      if(_zz_9)begin
        img_reg_array_7_8_real <= _zz_82;
      end
      if(_zz_10)begin
        img_reg_array_8_8_real <= _zz_82;
      end
      if(_zz_11)begin
        img_reg_array_9_8_real <= _zz_82;
      end
      if(_zz_12)begin
        img_reg_array_10_8_real <= _zz_82;
      end
      if(_zz_13)begin
        img_reg_array_11_8_real <= _zz_82;
      end
      if(_zz_14)begin
        img_reg_array_12_8_real <= _zz_82;
      end
      if(_zz_15)begin
        img_reg_array_13_8_real <= _zz_82;
      end
      if(_zz_16)begin
        img_reg_array_14_8_real <= _zz_82;
      end
      if(_zz_17)begin
        img_reg_array_15_8_real <= _zz_82;
      end
      if(_zz_18)begin
        img_reg_array_16_8_real <= _zz_82;
      end
      if(_zz_19)begin
        img_reg_array_17_8_real <= _zz_82;
      end
      if(_zz_20)begin
        img_reg_array_18_8_real <= _zz_82;
      end
      if(_zz_21)begin
        img_reg_array_19_8_real <= _zz_82;
      end
      if(_zz_22)begin
        img_reg_array_20_8_real <= _zz_82;
      end
      if(_zz_23)begin
        img_reg_array_21_8_real <= _zz_82;
      end
      if(_zz_24)begin
        img_reg_array_22_8_real <= _zz_82;
      end
      if(_zz_25)begin
        img_reg_array_23_8_real <= _zz_82;
      end
      if(_zz_26)begin
        img_reg_array_24_8_real <= _zz_82;
      end
      if(_zz_27)begin
        img_reg_array_25_8_real <= _zz_82;
      end
      if(_zz_28)begin
        img_reg_array_26_8_real <= _zz_82;
      end
      if(_zz_29)begin
        img_reg_array_27_8_real <= _zz_82;
      end
      if(_zz_30)begin
        img_reg_array_28_8_real <= _zz_82;
      end
      if(_zz_31)begin
        img_reg_array_29_8_real <= _zz_82;
      end
      if(_zz_32)begin
        img_reg_array_30_8_real <= _zz_82;
      end
      if(_zz_33)begin
        img_reg_array_31_8_real <= _zz_82;
      end
      if(_zz_34)begin
        img_reg_array_32_8_real <= _zz_82;
      end
      if(_zz_35)begin
        img_reg_array_33_8_real <= _zz_82;
      end
      if(_zz_36)begin
        img_reg_array_34_8_real <= _zz_82;
      end
      if(_zz_37)begin
        img_reg_array_35_8_real <= _zz_82;
      end
      if(_zz_38)begin
        img_reg_array_36_8_real <= _zz_82;
      end
      if(_zz_39)begin
        img_reg_array_37_8_real <= _zz_82;
      end
      if(_zz_40)begin
        img_reg_array_38_8_real <= _zz_82;
      end
      if(_zz_41)begin
        img_reg_array_39_8_real <= _zz_82;
      end
      if(_zz_42)begin
        img_reg_array_40_8_real <= _zz_82;
      end
      if(_zz_43)begin
        img_reg_array_41_8_real <= _zz_82;
      end
      if(_zz_44)begin
        img_reg_array_42_8_real <= _zz_82;
      end
      if(_zz_45)begin
        img_reg_array_43_8_real <= _zz_82;
      end
      if(_zz_46)begin
        img_reg_array_44_8_real <= _zz_82;
      end
      if(_zz_47)begin
        img_reg_array_45_8_real <= _zz_82;
      end
      if(_zz_48)begin
        img_reg_array_46_8_real <= _zz_82;
      end
      if(_zz_49)begin
        img_reg_array_47_8_real <= _zz_82;
      end
      if(_zz_50)begin
        img_reg_array_48_8_real <= _zz_82;
      end
      if(_zz_51)begin
        img_reg_array_49_8_real <= _zz_82;
      end
      if(_zz_52)begin
        img_reg_array_50_8_real <= _zz_82;
      end
      if(_zz_53)begin
        img_reg_array_51_8_real <= _zz_82;
      end
      if(_zz_54)begin
        img_reg_array_52_8_real <= _zz_82;
      end
      if(_zz_55)begin
        img_reg_array_53_8_real <= _zz_82;
      end
      if(_zz_56)begin
        img_reg_array_54_8_real <= _zz_82;
      end
      if(_zz_57)begin
        img_reg_array_55_8_real <= _zz_82;
      end
      if(_zz_58)begin
        img_reg_array_56_8_real <= _zz_82;
      end
      if(_zz_59)begin
        img_reg_array_57_8_real <= _zz_82;
      end
      if(_zz_60)begin
        img_reg_array_58_8_real <= _zz_82;
      end
      if(_zz_61)begin
        img_reg_array_59_8_real <= _zz_82;
      end
      if(_zz_62)begin
        img_reg_array_60_8_real <= _zz_82;
      end
      if(_zz_63)begin
        img_reg_array_61_8_real <= _zz_82;
      end
      if(_zz_64)begin
        img_reg_array_62_8_real <= _zz_82;
      end
      if(_zz_65)begin
        img_reg_array_63_8_real <= _zz_82;
      end
      if(_zz_2)begin
        img_reg_array_0_8_imag <= _zz_83;
      end
      if(_zz_3)begin
        img_reg_array_1_8_imag <= _zz_83;
      end
      if(_zz_4)begin
        img_reg_array_2_8_imag <= _zz_83;
      end
      if(_zz_5)begin
        img_reg_array_3_8_imag <= _zz_83;
      end
      if(_zz_6)begin
        img_reg_array_4_8_imag <= _zz_83;
      end
      if(_zz_7)begin
        img_reg_array_5_8_imag <= _zz_83;
      end
      if(_zz_8)begin
        img_reg_array_6_8_imag <= _zz_83;
      end
      if(_zz_9)begin
        img_reg_array_7_8_imag <= _zz_83;
      end
      if(_zz_10)begin
        img_reg_array_8_8_imag <= _zz_83;
      end
      if(_zz_11)begin
        img_reg_array_9_8_imag <= _zz_83;
      end
      if(_zz_12)begin
        img_reg_array_10_8_imag <= _zz_83;
      end
      if(_zz_13)begin
        img_reg_array_11_8_imag <= _zz_83;
      end
      if(_zz_14)begin
        img_reg_array_12_8_imag <= _zz_83;
      end
      if(_zz_15)begin
        img_reg_array_13_8_imag <= _zz_83;
      end
      if(_zz_16)begin
        img_reg_array_14_8_imag <= _zz_83;
      end
      if(_zz_17)begin
        img_reg_array_15_8_imag <= _zz_83;
      end
      if(_zz_18)begin
        img_reg_array_16_8_imag <= _zz_83;
      end
      if(_zz_19)begin
        img_reg_array_17_8_imag <= _zz_83;
      end
      if(_zz_20)begin
        img_reg_array_18_8_imag <= _zz_83;
      end
      if(_zz_21)begin
        img_reg_array_19_8_imag <= _zz_83;
      end
      if(_zz_22)begin
        img_reg_array_20_8_imag <= _zz_83;
      end
      if(_zz_23)begin
        img_reg_array_21_8_imag <= _zz_83;
      end
      if(_zz_24)begin
        img_reg_array_22_8_imag <= _zz_83;
      end
      if(_zz_25)begin
        img_reg_array_23_8_imag <= _zz_83;
      end
      if(_zz_26)begin
        img_reg_array_24_8_imag <= _zz_83;
      end
      if(_zz_27)begin
        img_reg_array_25_8_imag <= _zz_83;
      end
      if(_zz_28)begin
        img_reg_array_26_8_imag <= _zz_83;
      end
      if(_zz_29)begin
        img_reg_array_27_8_imag <= _zz_83;
      end
      if(_zz_30)begin
        img_reg_array_28_8_imag <= _zz_83;
      end
      if(_zz_31)begin
        img_reg_array_29_8_imag <= _zz_83;
      end
      if(_zz_32)begin
        img_reg_array_30_8_imag <= _zz_83;
      end
      if(_zz_33)begin
        img_reg_array_31_8_imag <= _zz_83;
      end
      if(_zz_34)begin
        img_reg_array_32_8_imag <= _zz_83;
      end
      if(_zz_35)begin
        img_reg_array_33_8_imag <= _zz_83;
      end
      if(_zz_36)begin
        img_reg_array_34_8_imag <= _zz_83;
      end
      if(_zz_37)begin
        img_reg_array_35_8_imag <= _zz_83;
      end
      if(_zz_38)begin
        img_reg_array_36_8_imag <= _zz_83;
      end
      if(_zz_39)begin
        img_reg_array_37_8_imag <= _zz_83;
      end
      if(_zz_40)begin
        img_reg_array_38_8_imag <= _zz_83;
      end
      if(_zz_41)begin
        img_reg_array_39_8_imag <= _zz_83;
      end
      if(_zz_42)begin
        img_reg_array_40_8_imag <= _zz_83;
      end
      if(_zz_43)begin
        img_reg_array_41_8_imag <= _zz_83;
      end
      if(_zz_44)begin
        img_reg_array_42_8_imag <= _zz_83;
      end
      if(_zz_45)begin
        img_reg_array_43_8_imag <= _zz_83;
      end
      if(_zz_46)begin
        img_reg_array_44_8_imag <= _zz_83;
      end
      if(_zz_47)begin
        img_reg_array_45_8_imag <= _zz_83;
      end
      if(_zz_48)begin
        img_reg_array_46_8_imag <= _zz_83;
      end
      if(_zz_49)begin
        img_reg_array_47_8_imag <= _zz_83;
      end
      if(_zz_50)begin
        img_reg_array_48_8_imag <= _zz_83;
      end
      if(_zz_51)begin
        img_reg_array_49_8_imag <= _zz_83;
      end
      if(_zz_52)begin
        img_reg_array_50_8_imag <= _zz_83;
      end
      if(_zz_53)begin
        img_reg_array_51_8_imag <= _zz_83;
      end
      if(_zz_54)begin
        img_reg_array_52_8_imag <= _zz_83;
      end
      if(_zz_55)begin
        img_reg_array_53_8_imag <= _zz_83;
      end
      if(_zz_56)begin
        img_reg_array_54_8_imag <= _zz_83;
      end
      if(_zz_57)begin
        img_reg_array_55_8_imag <= _zz_83;
      end
      if(_zz_58)begin
        img_reg_array_56_8_imag <= _zz_83;
      end
      if(_zz_59)begin
        img_reg_array_57_8_imag <= _zz_83;
      end
      if(_zz_60)begin
        img_reg_array_58_8_imag <= _zz_83;
      end
      if(_zz_61)begin
        img_reg_array_59_8_imag <= _zz_83;
      end
      if(_zz_62)begin
        img_reg_array_60_8_imag <= _zz_83;
      end
      if(_zz_63)begin
        img_reg_array_61_8_imag <= _zz_83;
      end
      if(_zz_64)begin
        img_reg_array_62_8_imag <= _zz_83;
      end
      if(_zz_65)begin
        img_reg_array_63_8_imag <= _zz_83;
      end
      if(_zz_2)begin
        img_reg_array_0_9_real <= _zz_84;
      end
      if(_zz_3)begin
        img_reg_array_1_9_real <= _zz_84;
      end
      if(_zz_4)begin
        img_reg_array_2_9_real <= _zz_84;
      end
      if(_zz_5)begin
        img_reg_array_3_9_real <= _zz_84;
      end
      if(_zz_6)begin
        img_reg_array_4_9_real <= _zz_84;
      end
      if(_zz_7)begin
        img_reg_array_5_9_real <= _zz_84;
      end
      if(_zz_8)begin
        img_reg_array_6_9_real <= _zz_84;
      end
      if(_zz_9)begin
        img_reg_array_7_9_real <= _zz_84;
      end
      if(_zz_10)begin
        img_reg_array_8_9_real <= _zz_84;
      end
      if(_zz_11)begin
        img_reg_array_9_9_real <= _zz_84;
      end
      if(_zz_12)begin
        img_reg_array_10_9_real <= _zz_84;
      end
      if(_zz_13)begin
        img_reg_array_11_9_real <= _zz_84;
      end
      if(_zz_14)begin
        img_reg_array_12_9_real <= _zz_84;
      end
      if(_zz_15)begin
        img_reg_array_13_9_real <= _zz_84;
      end
      if(_zz_16)begin
        img_reg_array_14_9_real <= _zz_84;
      end
      if(_zz_17)begin
        img_reg_array_15_9_real <= _zz_84;
      end
      if(_zz_18)begin
        img_reg_array_16_9_real <= _zz_84;
      end
      if(_zz_19)begin
        img_reg_array_17_9_real <= _zz_84;
      end
      if(_zz_20)begin
        img_reg_array_18_9_real <= _zz_84;
      end
      if(_zz_21)begin
        img_reg_array_19_9_real <= _zz_84;
      end
      if(_zz_22)begin
        img_reg_array_20_9_real <= _zz_84;
      end
      if(_zz_23)begin
        img_reg_array_21_9_real <= _zz_84;
      end
      if(_zz_24)begin
        img_reg_array_22_9_real <= _zz_84;
      end
      if(_zz_25)begin
        img_reg_array_23_9_real <= _zz_84;
      end
      if(_zz_26)begin
        img_reg_array_24_9_real <= _zz_84;
      end
      if(_zz_27)begin
        img_reg_array_25_9_real <= _zz_84;
      end
      if(_zz_28)begin
        img_reg_array_26_9_real <= _zz_84;
      end
      if(_zz_29)begin
        img_reg_array_27_9_real <= _zz_84;
      end
      if(_zz_30)begin
        img_reg_array_28_9_real <= _zz_84;
      end
      if(_zz_31)begin
        img_reg_array_29_9_real <= _zz_84;
      end
      if(_zz_32)begin
        img_reg_array_30_9_real <= _zz_84;
      end
      if(_zz_33)begin
        img_reg_array_31_9_real <= _zz_84;
      end
      if(_zz_34)begin
        img_reg_array_32_9_real <= _zz_84;
      end
      if(_zz_35)begin
        img_reg_array_33_9_real <= _zz_84;
      end
      if(_zz_36)begin
        img_reg_array_34_9_real <= _zz_84;
      end
      if(_zz_37)begin
        img_reg_array_35_9_real <= _zz_84;
      end
      if(_zz_38)begin
        img_reg_array_36_9_real <= _zz_84;
      end
      if(_zz_39)begin
        img_reg_array_37_9_real <= _zz_84;
      end
      if(_zz_40)begin
        img_reg_array_38_9_real <= _zz_84;
      end
      if(_zz_41)begin
        img_reg_array_39_9_real <= _zz_84;
      end
      if(_zz_42)begin
        img_reg_array_40_9_real <= _zz_84;
      end
      if(_zz_43)begin
        img_reg_array_41_9_real <= _zz_84;
      end
      if(_zz_44)begin
        img_reg_array_42_9_real <= _zz_84;
      end
      if(_zz_45)begin
        img_reg_array_43_9_real <= _zz_84;
      end
      if(_zz_46)begin
        img_reg_array_44_9_real <= _zz_84;
      end
      if(_zz_47)begin
        img_reg_array_45_9_real <= _zz_84;
      end
      if(_zz_48)begin
        img_reg_array_46_9_real <= _zz_84;
      end
      if(_zz_49)begin
        img_reg_array_47_9_real <= _zz_84;
      end
      if(_zz_50)begin
        img_reg_array_48_9_real <= _zz_84;
      end
      if(_zz_51)begin
        img_reg_array_49_9_real <= _zz_84;
      end
      if(_zz_52)begin
        img_reg_array_50_9_real <= _zz_84;
      end
      if(_zz_53)begin
        img_reg_array_51_9_real <= _zz_84;
      end
      if(_zz_54)begin
        img_reg_array_52_9_real <= _zz_84;
      end
      if(_zz_55)begin
        img_reg_array_53_9_real <= _zz_84;
      end
      if(_zz_56)begin
        img_reg_array_54_9_real <= _zz_84;
      end
      if(_zz_57)begin
        img_reg_array_55_9_real <= _zz_84;
      end
      if(_zz_58)begin
        img_reg_array_56_9_real <= _zz_84;
      end
      if(_zz_59)begin
        img_reg_array_57_9_real <= _zz_84;
      end
      if(_zz_60)begin
        img_reg_array_58_9_real <= _zz_84;
      end
      if(_zz_61)begin
        img_reg_array_59_9_real <= _zz_84;
      end
      if(_zz_62)begin
        img_reg_array_60_9_real <= _zz_84;
      end
      if(_zz_63)begin
        img_reg_array_61_9_real <= _zz_84;
      end
      if(_zz_64)begin
        img_reg_array_62_9_real <= _zz_84;
      end
      if(_zz_65)begin
        img_reg_array_63_9_real <= _zz_84;
      end
      if(_zz_2)begin
        img_reg_array_0_9_imag <= _zz_85;
      end
      if(_zz_3)begin
        img_reg_array_1_9_imag <= _zz_85;
      end
      if(_zz_4)begin
        img_reg_array_2_9_imag <= _zz_85;
      end
      if(_zz_5)begin
        img_reg_array_3_9_imag <= _zz_85;
      end
      if(_zz_6)begin
        img_reg_array_4_9_imag <= _zz_85;
      end
      if(_zz_7)begin
        img_reg_array_5_9_imag <= _zz_85;
      end
      if(_zz_8)begin
        img_reg_array_6_9_imag <= _zz_85;
      end
      if(_zz_9)begin
        img_reg_array_7_9_imag <= _zz_85;
      end
      if(_zz_10)begin
        img_reg_array_8_9_imag <= _zz_85;
      end
      if(_zz_11)begin
        img_reg_array_9_9_imag <= _zz_85;
      end
      if(_zz_12)begin
        img_reg_array_10_9_imag <= _zz_85;
      end
      if(_zz_13)begin
        img_reg_array_11_9_imag <= _zz_85;
      end
      if(_zz_14)begin
        img_reg_array_12_9_imag <= _zz_85;
      end
      if(_zz_15)begin
        img_reg_array_13_9_imag <= _zz_85;
      end
      if(_zz_16)begin
        img_reg_array_14_9_imag <= _zz_85;
      end
      if(_zz_17)begin
        img_reg_array_15_9_imag <= _zz_85;
      end
      if(_zz_18)begin
        img_reg_array_16_9_imag <= _zz_85;
      end
      if(_zz_19)begin
        img_reg_array_17_9_imag <= _zz_85;
      end
      if(_zz_20)begin
        img_reg_array_18_9_imag <= _zz_85;
      end
      if(_zz_21)begin
        img_reg_array_19_9_imag <= _zz_85;
      end
      if(_zz_22)begin
        img_reg_array_20_9_imag <= _zz_85;
      end
      if(_zz_23)begin
        img_reg_array_21_9_imag <= _zz_85;
      end
      if(_zz_24)begin
        img_reg_array_22_9_imag <= _zz_85;
      end
      if(_zz_25)begin
        img_reg_array_23_9_imag <= _zz_85;
      end
      if(_zz_26)begin
        img_reg_array_24_9_imag <= _zz_85;
      end
      if(_zz_27)begin
        img_reg_array_25_9_imag <= _zz_85;
      end
      if(_zz_28)begin
        img_reg_array_26_9_imag <= _zz_85;
      end
      if(_zz_29)begin
        img_reg_array_27_9_imag <= _zz_85;
      end
      if(_zz_30)begin
        img_reg_array_28_9_imag <= _zz_85;
      end
      if(_zz_31)begin
        img_reg_array_29_9_imag <= _zz_85;
      end
      if(_zz_32)begin
        img_reg_array_30_9_imag <= _zz_85;
      end
      if(_zz_33)begin
        img_reg_array_31_9_imag <= _zz_85;
      end
      if(_zz_34)begin
        img_reg_array_32_9_imag <= _zz_85;
      end
      if(_zz_35)begin
        img_reg_array_33_9_imag <= _zz_85;
      end
      if(_zz_36)begin
        img_reg_array_34_9_imag <= _zz_85;
      end
      if(_zz_37)begin
        img_reg_array_35_9_imag <= _zz_85;
      end
      if(_zz_38)begin
        img_reg_array_36_9_imag <= _zz_85;
      end
      if(_zz_39)begin
        img_reg_array_37_9_imag <= _zz_85;
      end
      if(_zz_40)begin
        img_reg_array_38_9_imag <= _zz_85;
      end
      if(_zz_41)begin
        img_reg_array_39_9_imag <= _zz_85;
      end
      if(_zz_42)begin
        img_reg_array_40_9_imag <= _zz_85;
      end
      if(_zz_43)begin
        img_reg_array_41_9_imag <= _zz_85;
      end
      if(_zz_44)begin
        img_reg_array_42_9_imag <= _zz_85;
      end
      if(_zz_45)begin
        img_reg_array_43_9_imag <= _zz_85;
      end
      if(_zz_46)begin
        img_reg_array_44_9_imag <= _zz_85;
      end
      if(_zz_47)begin
        img_reg_array_45_9_imag <= _zz_85;
      end
      if(_zz_48)begin
        img_reg_array_46_9_imag <= _zz_85;
      end
      if(_zz_49)begin
        img_reg_array_47_9_imag <= _zz_85;
      end
      if(_zz_50)begin
        img_reg_array_48_9_imag <= _zz_85;
      end
      if(_zz_51)begin
        img_reg_array_49_9_imag <= _zz_85;
      end
      if(_zz_52)begin
        img_reg_array_50_9_imag <= _zz_85;
      end
      if(_zz_53)begin
        img_reg_array_51_9_imag <= _zz_85;
      end
      if(_zz_54)begin
        img_reg_array_52_9_imag <= _zz_85;
      end
      if(_zz_55)begin
        img_reg_array_53_9_imag <= _zz_85;
      end
      if(_zz_56)begin
        img_reg_array_54_9_imag <= _zz_85;
      end
      if(_zz_57)begin
        img_reg_array_55_9_imag <= _zz_85;
      end
      if(_zz_58)begin
        img_reg_array_56_9_imag <= _zz_85;
      end
      if(_zz_59)begin
        img_reg_array_57_9_imag <= _zz_85;
      end
      if(_zz_60)begin
        img_reg_array_58_9_imag <= _zz_85;
      end
      if(_zz_61)begin
        img_reg_array_59_9_imag <= _zz_85;
      end
      if(_zz_62)begin
        img_reg_array_60_9_imag <= _zz_85;
      end
      if(_zz_63)begin
        img_reg_array_61_9_imag <= _zz_85;
      end
      if(_zz_64)begin
        img_reg_array_62_9_imag <= _zz_85;
      end
      if(_zz_65)begin
        img_reg_array_63_9_imag <= _zz_85;
      end
      if(_zz_2)begin
        img_reg_array_0_10_real <= _zz_86;
      end
      if(_zz_3)begin
        img_reg_array_1_10_real <= _zz_86;
      end
      if(_zz_4)begin
        img_reg_array_2_10_real <= _zz_86;
      end
      if(_zz_5)begin
        img_reg_array_3_10_real <= _zz_86;
      end
      if(_zz_6)begin
        img_reg_array_4_10_real <= _zz_86;
      end
      if(_zz_7)begin
        img_reg_array_5_10_real <= _zz_86;
      end
      if(_zz_8)begin
        img_reg_array_6_10_real <= _zz_86;
      end
      if(_zz_9)begin
        img_reg_array_7_10_real <= _zz_86;
      end
      if(_zz_10)begin
        img_reg_array_8_10_real <= _zz_86;
      end
      if(_zz_11)begin
        img_reg_array_9_10_real <= _zz_86;
      end
      if(_zz_12)begin
        img_reg_array_10_10_real <= _zz_86;
      end
      if(_zz_13)begin
        img_reg_array_11_10_real <= _zz_86;
      end
      if(_zz_14)begin
        img_reg_array_12_10_real <= _zz_86;
      end
      if(_zz_15)begin
        img_reg_array_13_10_real <= _zz_86;
      end
      if(_zz_16)begin
        img_reg_array_14_10_real <= _zz_86;
      end
      if(_zz_17)begin
        img_reg_array_15_10_real <= _zz_86;
      end
      if(_zz_18)begin
        img_reg_array_16_10_real <= _zz_86;
      end
      if(_zz_19)begin
        img_reg_array_17_10_real <= _zz_86;
      end
      if(_zz_20)begin
        img_reg_array_18_10_real <= _zz_86;
      end
      if(_zz_21)begin
        img_reg_array_19_10_real <= _zz_86;
      end
      if(_zz_22)begin
        img_reg_array_20_10_real <= _zz_86;
      end
      if(_zz_23)begin
        img_reg_array_21_10_real <= _zz_86;
      end
      if(_zz_24)begin
        img_reg_array_22_10_real <= _zz_86;
      end
      if(_zz_25)begin
        img_reg_array_23_10_real <= _zz_86;
      end
      if(_zz_26)begin
        img_reg_array_24_10_real <= _zz_86;
      end
      if(_zz_27)begin
        img_reg_array_25_10_real <= _zz_86;
      end
      if(_zz_28)begin
        img_reg_array_26_10_real <= _zz_86;
      end
      if(_zz_29)begin
        img_reg_array_27_10_real <= _zz_86;
      end
      if(_zz_30)begin
        img_reg_array_28_10_real <= _zz_86;
      end
      if(_zz_31)begin
        img_reg_array_29_10_real <= _zz_86;
      end
      if(_zz_32)begin
        img_reg_array_30_10_real <= _zz_86;
      end
      if(_zz_33)begin
        img_reg_array_31_10_real <= _zz_86;
      end
      if(_zz_34)begin
        img_reg_array_32_10_real <= _zz_86;
      end
      if(_zz_35)begin
        img_reg_array_33_10_real <= _zz_86;
      end
      if(_zz_36)begin
        img_reg_array_34_10_real <= _zz_86;
      end
      if(_zz_37)begin
        img_reg_array_35_10_real <= _zz_86;
      end
      if(_zz_38)begin
        img_reg_array_36_10_real <= _zz_86;
      end
      if(_zz_39)begin
        img_reg_array_37_10_real <= _zz_86;
      end
      if(_zz_40)begin
        img_reg_array_38_10_real <= _zz_86;
      end
      if(_zz_41)begin
        img_reg_array_39_10_real <= _zz_86;
      end
      if(_zz_42)begin
        img_reg_array_40_10_real <= _zz_86;
      end
      if(_zz_43)begin
        img_reg_array_41_10_real <= _zz_86;
      end
      if(_zz_44)begin
        img_reg_array_42_10_real <= _zz_86;
      end
      if(_zz_45)begin
        img_reg_array_43_10_real <= _zz_86;
      end
      if(_zz_46)begin
        img_reg_array_44_10_real <= _zz_86;
      end
      if(_zz_47)begin
        img_reg_array_45_10_real <= _zz_86;
      end
      if(_zz_48)begin
        img_reg_array_46_10_real <= _zz_86;
      end
      if(_zz_49)begin
        img_reg_array_47_10_real <= _zz_86;
      end
      if(_zz_50)begin
        img_reg_array_48_10_real <= _zz_86;
      end
      if(_zz_51)begin
        img_reg_array_49_10_real <= _zz_86;
      end
      if(_zz_52)begin
        img_reg_array_50_10_real <= _zz_86;
      end
      if(_zz_53)begin
        img_reg_array_51_10_real <= _zz_86;
      end
      if(_zz_54)begin
        img_reg_array_52_10_real <= _zz_86;
      end
      if(_zz_55)begin
        img_reg_array_53_10_real <= _zz_86;
      end
      if(_zz_56)begin
        img_reg_array_54_10_real <= _zz_86;
      end
      if(_zz_57)begin
        img_reg_array_55_10_real <= _zz_86;
      end
      if(_zz_58)begin
        img_reg_array_56_10_real <= _zz_86;
      end
      if(_zz_59)begin
        img_reg_array_57_10_real <= _zz_86;
      end
      if(_zz_60)begin
        img_reg_array_58_10_real <= _zz_86;
      end
      if(_zz_61)begin
        img_reg_array_59_10_real <= _zz_86;
      end
      if(_zz_62)begin
        img_reg_array_60_10_real <= _zz_86;
      end
      if(_zz_63)begin
        img_reg_array_61_10_real <= _zz_86;
      end
      if(_zz_64)begin
        img_reg_array_62_10_real <= _zz_86;
      end
      if(_zz_65)begin
        img_reg_array_63_10_real <= _zz_86;
      end
      if(_zz_2)begin
        img_reg_array_0_10_imag <= _zz_87;
      end
      if(_zz_3)begin
        img_reg_array_1_10_imag <= _zz_87;
      end
      if(_zz_4)begin
        img_reg_array_2_10_imag <= _zz_87;
      end
      if(_zz_5)begin
        img_reg_array_3_10_imag <= _zz_87;
      end
      if(_zz_6)begin
        img_reg_array_4_10_imag <= _zz_87;
      end
      if(_zz_7)begin
        img_reg_array_5_10_imag <= _zz_87;
      end
      if(_zz_8)begin
        img_reg_array_6_10_imag <= _zz_87;
      end
      if(_zz_9)begin
        img_reg_array_7_10_imag <= _zz_87;
      end
      if(_zz_10)begin
        img_reg_array_8_10_imag <= _zz_87;
      end
      if(_zz_11)begin
        img_reg_array_9_10_imag <= _zz_87;
      end
      if(_zz_12)begin
        img_reg_array_10_10_imag <= _zz_87;
      end
      if(_zz_13)begin
        img_reg_array_11_10_imag <= _zz_87;
      end
      if(_zz_14)begin
        img_reg_array_12_10_imag <= _zz_87;
      end
      if(_zz_15)begin
        img_reg_array_13_10_imag <= _zz_87;
      end
      if(_zz_16)begin
        img_reg_array_14_10_imag <= _zz_87;
      end
      if(_zz_17)begin
        img_reg_array_15_10_imag <= _zz_87;
      end
      if(_zz_18)begin
        img_reg_array_16_10_imag <= _zz_87;
      end
      if(_zz_19)begin
        img_reg_array_17_10_imag <= _zz_87;
      end
      if(_zz_20)begin
        img_reg_array_18_10_imag <= _zz_87;
      end
      if(_zz_21)begin
        img_reg_array_19_10_imag <= _zz_87;
      end
      if(_zz_22)begin
        img_reg_array_20_10_imag <= _zz_87;
      end
      if(_zz_23)begin
        img_reg_array_21_10_imag <= _zz_87;
      end
      if(_zz_24)begin
        img_reg_array_22_10_imag <= _zz_87;
      end
      if(_zz_25)begin
        img_reg_array_23_10_imag <= _zz_87;
      end
      if(_zz_26)begin
        img_reg_array_24_10_imag <= _zz_87;
      end
      if(_zz_27)begin
        img_reg_array_25_10_imag <= _zz_87;
      end
      if(_zz_28)begin
        img_reg_array_26_10_imag <= _zz_87;
      end
      if(_zz_29)begin
        img_reg_array_27_10_imag <= _zz_87;
      end
      if(_zz_30)begin
        img_reg_array_28_10_imag <= _zz_87;
      end
      if(_zz_31)begin
        img_reg_array_29_10_imag <= _zz_87;
      end
      if(_zz_32)begin
        img_reg_array_30_10_imag <= _zz_87;
      end
      if(_zz_33)begin
        img_reg_array_31_10_imag <= _zz_87;
      end
      if(_zz_34)begin
        img_reg_array_32_10_imag <= _zz_87;
      end
      if(_zz_35)begin
        img_reg_array_33_10_imag <= _zz_87;
      end
      if(_zz_36)begin
        img_reg_array_34_10_imag <= _zz_87;
      end
      if(_zz_37)begin
        img_reg_array_35_10_imag <= _zz_87;
      end
      if(_zz_38)begin
        img_reg_array_36_10_imag <= _zz_87;
      end
      if(_zz_39)begin
        img_reg_array_37_10_imag <= _zz_87;
      end
      if(_zz_40)begin
        img_reg_array_38_10_imag <= _zz_87;
      end
      if(_zz_41)begin
        img_reg_array_39_10_imag <= _zz_87;
      end
      if(_zz_42)begin
        img_reg_array_40_10_imag <= _zz_87;
      end
      if(_zz_43)begin
        img_reg_array_41_10_imag <= _zz_87;
      end
      if(_zz_44)begin
        img_reg_array_42_10_imag <= _zz_87;
      end
      if(_zz_45)begin
        img_reg_array_43_10_imag <= _zz_87;
      end
      if(_zz_46)begin
        img_reg_array_44_10_imag <= _zz_87;
      end
      if(_zz_47)begin
        img_reg_array_45_10_imag <= _zz_87;
      end
      if(_zz_48)begin
        img_reg_array_46_10_imag <= _zz_87;
      end
      if(_zz_49)begin
        img_reg_array_47_10_imag <= _zz_87;
      end
      if(_zz_50)begin
        img_reg_array_48_10_imag <= _zz_87;
      end
      if(_zz_51)begin
        img_reg_array_49_10_imag <= _zz_87;
      end
      if(_zz_52)begin
        img_reg_array_50_10_imag <= _zz_87;
      end
      if(_zz_53)begin
        img_reg_array_51_10_imag <= _zz_87;
      end
      if(_zz_54)begin
        img_reg_array_52_10_imag <= _zz_87;
      end
      if(_zz_55)begin
        img_reg_array_53_10_imag <= _zz_87;
      end
      if(_zz_56)begin
        img_reg_array_54_10_imag <= _zz_87;
      end
      if(_zz_57)begin
        img_reg_array_55_10_imag <= _zz_87;
      end
      if(_zz_58)begin
        img_reg_array_56_10_imag <= _zz_87;
      end
      if(_zz_59)begin
        img_reg_array_57_10_imag <= _zz_87;
      end
      if(_zz_60)begin
        img_reg_array_58_10_imag <= _zz_87;
      end
      if(_zz_61)begin
        img_reg_array_59_10_imag <= _zz_87;
      end
      if(_zz_62)begin
        img_reg_array_60_10_imag <= _zz_87;
      end
      if(_zz_63)begin
        img_reg_array_61_10_imag <= _zz_87;
      end
      if(_zz_64)begin
        img_reg_array_62_10_imag <= _zz_87;
      end
      if(_zz_65)begin
        img_reg_array_63_10_imag <= _zz_87;
      end
      if(_zz_2)begin
        img_reg_array_0_11_real <= _zz_88;
      end
      if(_zz_3)begin
        img_reg_array_1_11_real <= _zz_88;
      end
      if(_zz_4)begin
        img_reg_array_2_11_real <= _zz_88;
      end
      if(_zz_5)begin
        img_reg_array_3_11_real <= _zz_88;
      end
      if(_zz_6)begin
        img_reg_array_4_11_real <= _zz_88;
      end
      if(_zz_7)begin
        img_reg_array_5_11_real <= _zz_88;
      end
      if(_zz_8)begin
        img_reg_array_6_11_real <= _zz_88;
      end
      if(_zz_9)begin
        img_reg_array_7_11_real <= _zz_88;
      end
      if(_zz_10)begin
        img_reg_array_8_11_real <= _zz_88;
      end
      if(_zz_11)begin
        img_reg_array_9_11_real <= _zz_88;
      end
      if(_zz_12)begin
        img_reg_array_10_11_real <= _zz_88;
      end
      if(_zz_13)begin
        img_reg_array_11_11_real <= _zz_88;
      end
      if(_zz_14)begin
        img_reg_array_12_11_real <= _zz_88;
      end
      if(_zz_15)begin
        img_reg_array_13_11_real <= _zz_88;
      end
      if(_zz_16)begin
        img_reg_array_14_11_real <= _zz_88;
      end
      if(_zz_17)begin
        img_reg_array_15_11_real <= _zz_88;
      end
      if(_zz_18)begin
        img_reg_array_16_11_real <= _zz_88;
      end
      if(_zz_19)begin
        img_reg_array_17_11_real <= _zz_88;
      end
      if(_zz_20)begin
        img_reg_array_18_11_real <= _zz_88;
      end
      if(_zz_21)begin
        img_reg_array_19_11_real <= _zz_88;
      end
      if(_zz_22)begin
        img_reg_array_20_11_real <= _zz_88;
      end
      if(_zz_23)begin
        img_reg_array_21_11_real <= _zz_88;
      end
      if(_zz_24)begin
        img_reg_array_22_11_real <= _zz_88;
      end
      if(_zz_25)begin
        img_reg_array_23_11_real <= _zz_88;
      end
      if(_zz_26)begin
        img_reg_array_24_11_real <= _zz_88;
      end
      if(_zz_27)begin
        img_reg_array_25_11_real <= _zz_88;
      end
      if(_zz_28)begin
        img_reg_array_26_11_real <= _zz_88;
      end
      if(_zz_29)begin
        img_reg_array_27_11_real <= _zz_88;
      end
      if(_zz_30)begin
        img_reg_array_28_11_real <= _zz_88;
      end
      if(_zz_31)begin
        img_reg_array_29_11_real <= _zz_88;
      end
      if(_zz_32)begin
        img_reg_array_30_11_real <= _zz_88;
      end
      if(_zz_33)begin
        img_reg_array_31_11_real <= _zz_88;
      end
      if(_zz_34)begin
        img_reg_array_32_11_real <= _zz_88;
      end
      if(_zz_35)begin
        img_reg_array_33_11_real <= _zz_88;
      end
      if(_zz_36)begin
        img_reg_array_34_11_real <= _zz_88;
      end
      if(_zz_37)begin
        img_reg_array_35_11_real <= _zz_88;
      end
      if(_zz_38)begin
        img_reg_array_36_11_real <= _zz_88;
      end
      if(_zz_39)begin
        img_reg_array_37_11_real <= _zz_88;
      end
      if(_zz_40)begin
        img_reg_array_38_11_real <= _zz_88;
      end
      if(_zz_41)begin
        img_reg_array_39_11_real <= _zz_88;
      end
      if(_zz_42)begin
        img_reg_array_40_11_real <= _zz_88;
      end
      if(_zz_43)begin
        img_reg_array_41_11_real <= _zz_88;
      end
      if(_zz_44)begin
        img_reg_array_42_11_real <= _zz_88;
      end
      if(_zz_45)begin
        img_reg_array_43_11_real <= _zz_88;
      end
      if(_zz_46)begin
        img_reg_array_44_11_real <= _zz_88;
      end
      if(_zz_47)begin
        img_reg_array_45_11_real <= _zz_88;
      end
      if(_zz_48)begin
        img_reg_array_46_11_real <= _zz_88;
      end
      if(_zz_49)begin
        img_reg_array_47_11_real <= _zz_88;
      end
      if(_zz_50)begin
        img_reg_array_48_11_real <= _zz_88;
      end
      if(_zz_51)begin
        img_reg_array_49_11_real <= _zz_88;
      end
      if(_zz_52)begin
        img_reg_array_50_11_real <= _zz_88;
      end
      if(_zz_53)begin
        img_reg_array_51_11_real <= _zz_88;
      end
      if(_zz_54)begin
        img_reg_array_52_11_real <= _zz_88;
      end
      if(_zz_55)begin
        img_reg_array_53_11_real <= _zz_88;
      end
      if(_zz_56)begin
        img_reg_array_54_11_real <= _zz_88;
      end
      if(_zz_57)begin
        img_reg_array_55_11_real <= _zz_88;
      end
      if(_zz_58)begin
        img_reg_array_56_11_real <= _zz_88;
      end
      if(_zz_59)begin
        img_reg_array_57_11_real <= _zz_88;
      end
      if(_zz_60)begin
        img_reg_array_58_11_real <= _zz_88;
      end
      if(_zz_61)begin
        img_reg_array_59_11_real <= _zz_88;
      end
      if(_zz_62)begin
        img_reg_array_60_11_real <= _zz_88;
      end
      if(_zz_63)begin
        img_reg_array_61_11_real <= _zz_88;
      end
      if(_zz_64)begin
        img_reg_array_62_11_real <= _zz_88;
      end
      if(_zz_65)begin
        img_reg_array_63_11_real <= _zz_88;
      end
      if(_zz_2)begin
        img_reg_array_0_11_imag <= _zz_89;
      end
      if(_zz_3)begin
        img_reg_array_1_11_imag <= _zz_89;
      end
      if(_zz_4)begin
        img_reg_array_2_11_imag <= _zz_89;
      end
      if(_zz_5)begin
        img_reg_array_3_11_imag <= _zz_89;
      end
      if(_zz_6)begin
        img_reg_array_4_11_imag <= _zz_89;
      end
      if(_zz_7)begin
        img_reg_array_5_11_imag <= _zz_89;
      end
      if(_zz_8)begin
        img_reg_array_6_11_imag <= _zz_89;
      end
      if(_zz_9)begin
        img_reg_array_7_11_imag <= _zz_89;
      end
      if(_zz_10)begin
        img_reg_array_8_11_imag <= _zz_89;
      end
      if(_zz_11)begin
        img_reg_array_9_11_imag <= _zz_89;
      end
      if(_zz_12)begin
        img_reg_array_10_11_imag <= _zz_89;
      end
      if(_zz_13)begin
        img_reg_array_11_11_imag <= _zz_89;
      end
      if(_zz_14)begin
        img_reg_array_12_11_imag <= _zz_89;
      end
      if(_zz_15)begin
        img_reg_array_13_11_imag <= _zz_89;
      end
      if(_zz_16)begin
        img_reg_array_14_11_imag <= _zz_89;
      end
      if(_zz_17)begin
        img_reg_array_15_11_imag <= _zz_89;
      end
      if(_zz_18)begin
        img_reg_array_16_11_imag <= _zz_89;
      end
      if(_zz_19)begin
        img_reg_array_17_11_imag <= _zz_89;
      end
      if(_zz_20)begin
        img_reg_array_18_11_imag <= _zz_89;
      end
      if(_zz_21)begin
        img_reg_array_19_11_imag <= _zz_89;
      end
      if(_zz_22)begin
        img_reg_array_20_11_imag <= _zz_89;
      end
      if(_zz_23)begin
        img_reg_array_21_11_imag <= _zz_89;
      end
      if(_zz_24)begin
        img_reg_array_22_11_imag <= _zz_89;
      end
      if(_zz_25)begin
        img_reg_array_23_11_imag <= _zz_89;
      end
      if(_zz_26)begin
        img_reg_array_24_11_imag <= _zz_89;
      end
      if(_zz_27)begin
        img_reg_array_25_11_imag <= _zz_89;
      end
      if(_zz_28)begin
        img_reg_array_26_11_imag <= _zz_89;
      end
      if(_zz_29)begin
        img_reg_array_27_11_imag <= _zz_89;
      end
      if(_zz_30)begin
        img_reg_array_28_11_imag <= _zz_89;
      end
      if(_zz_31)begin
        img_reg_array_29_11_imag <= _zz_89;
      end
      if(_zz_32)begin
        img_reg_array_30_11_imag <= _zz_89;
      end
      if(_zz_33)begin
        img_reg_array_31_11_imag <= _zz_89;
      end
      if(_zz_34)begin
        img_reg_array_32_11_imag <= _zz_89;
      end
      if(_zz_35)begin
        img_reg_array_33_11_imag <= _zz_89;
      end
      if(_zz_36)begin
        img_reg_array_34_11_imag <= _zz_89;
      end
      if(_zz_37)begin
        img_reg_array_35_11_imag <= _zz_89;
      end
      if(_zz_38)begin
        img_reg_array_36_11_imag <= _zz_89;
      end
      if(_zz_39)begin
        img_reg_array_37_11_imag <= _zz_89;
      end
      if(_zz_40)begin
        img_reg_array_38_11_imag <= _zz_89;
      end
      if(_zz_41)begin
        img_reg_array_39_11_imag <= _zz_89;
      end
      if(_zz_42)begin
        img_reg_array_40_11_imag <= _zz_89;
      end
      if(_zz_43)begin
        img_reg_array_41_11_imag <= _zz_89;
      end
      if(_zz_44)begin
        img_reg_array_42_11_imag <= _zz_89;
      end
      if(_zz_45)begin
        img_reg_array_43_11_imag <= _zz_89;
      end
      if(_zz_46)begin
        img_reg_array_44_11_imag <= _zz_89;
      end
      if(_zz_47)begin
        img_reg_array_45_11_imag <= _zz_89;
      end
      if(_zz_48)begin
        img_reg_array_46_11_imag <= _zz_89;
      end
      if(_zz_49)begin
        img_reg_array_47_11_imag <= _zz_89;
      end
      if(_zz_50)begin
        img_reg_array_48_11_imag <= _zz_89;
      end
      if(_zz_51)begin
        img_reg_array_49_11_imag <= _zz_89;
      end
      if(_zz_52)begin
        img_reg_array_50_11_imag <= _zz_89;
      end
      if(_zz_53)begin
        img_reg_array_51_11_imag <= _zz_89;
      end
      if(_zz_54)begin
        img_reg_array_52_11_imag <= _zz_89;
      end
      if(_zz_55)begin
        img_reg_array_53_11_imag <= _zz_89;
      end
      if(_zz_56)begin
        img_reg_array_54_11_imag <= _zz_89;
      end
      if(_zz_57)begin
        img_reg_array_55_11_imag <= _zz_89;
      end
      if(_zz_58)begin
        img_reg_array_56_11_imag <= _zz_89;
      end
      if(_zz_59)begin
        img_reg_array_57_11_imag <= _zz_89;
      end
      if(_zz_60)begin
        img_reg_array_58_11_imag <= _zz_89;
      end
      if(_zz_61)begin
        img_reg_array_59_11_imag <= _zz_89;
      end
      if(_zz_62)begin
        img_reg_array_60_11_imag <= _zz_89;
      end
      if(_zz_63)begin
        img_reg_array_61_11_imag <= _zz_89;
      end
      if(_zz_64)begin
        img_reg_array_62_11_imag <= _zz_89;
      end
      if(_zz_65)begin
        img_reg_array_63_11_imag <= _zz_89;
      end
      if(_zz_2)begin
        img_reg_array_0_12_real <= _zz_90;
      end
      if(_zz_3)begin
        img_reg_array_1_12_real <= _zz_90;
      end
      if(_zz_4)begin
        img_reg_array_2_12_real <= _zz_90;
      end
      if(_zz_5)begin
        img_reg_array_3_12_real <= _zz_90;
      end
      if(_zz_6)begin
        img_reg_array_4_12_real <= _zz_90;
      end
      if(_zz_7)begin
        img_reg_array_5_12_real <= _zz_90;
      end
      if(_zz_8)begin
        img_reg_array_6_12_real <= _zz_90;
      end
      if(_zz_9)begin
        img_reg_array_7_12_real <= _zz_90;
      end
      if(_zz_10)begin
        img_reg_array_8_12_real <= _zz_90;
      end
      if(_zz_11)begin
        img_reg_array_9_12_real <= _zz_90;
      end
      if(_zz_12)begin
        img_reg_array_10_12_real <= _zz_90;
      end
      if(_zz_13)begin
        img_reg_array_11_12_real <= _zz_90;
      end
      if(_zz_14)begin
        img_reg_array_12_12_real <= _zz_90;
      end
      if(_zz_15)begin
        img_reg_array_13_12_real <= _zz_90;
      end
      if(_zz_16)begin
        img_reg_array_14_12_real <= _zz_90;
      end
      if(_zz_17)begin
        img_reg_array_15_12_real <= _zz_90;
      end
      if(_zz_18)begin
        img_reg_array_16_12_real <= _zz_90;
      end
      if(_zz_19)begin
        img_reg_array_17_12_real <= _zz_90;
      end
      if(_zz_20)begin
        img_reg_array_18_12_real <= _zz_90;
      end
      if(_zz_21)begin
        img_reg_array_19_12_real <= _zz_90;
      end
      if(_zz_22)begin
        img_reg_array_20_12_real <= _zz_90;
      end
      if(_zz_23)begin
        img_reg_array_21_12_real <= _zz_90;
      end
      if(_zz_24)begin
        img_reg_array_22_12_real <= _zz_90;
      end
      if(_zz_25)begin
        img_reg_array_23_12_real <= _zz_90;
      end
      if(_zz_26)begin
        img_reg_array_24_12_real <= _zz_90;
      end
      if(_zz_27)begin
        img_reg_array_25_12_real <= _zz_90;
      end
      if(_zz_28)begin
        img_reg_array_26_12_real <= _zz_90;
      end
      if(_zz_29)begin
        img_reg_array_27_12_real <= _zz_90;
      end
      if(_zz_30)begin
        img_reg_array_28_12_real <= _zz_90;
      end
      if(_zz_31)begin
        img_reg_array_29_12_real <= _zz_90;
      end
      if(_zz_32)begin
        img_reg_array_30_12_real <= _zz_90;
      end
      if(_zz_33)begin
        img_reg_array_31_12_real <= _zz_90;
      end
      if(_zz_34)begin
        img_reg_array_32_12_real <= _zz_90;
      end
      if(_zz_35)begin
        img_reg_array_33_12_real <= _zz_90;
      end
      if(_zz_36)begin
        img_reg_array_34_12_real <= _zz_90;
      end
      if(_zz_37)begin
        img_reg_array_35_12_real <= _zz_90;
      end
      if(_zz_38)begin
        img_reg_array_36_12_real <= _zz_90;
      end
      if(_zz_39)begin
        img_reg_array_37_12_real <= _zz_90;
      end
      if(_zz_40)begin
        img_reg_array_38_12_real <= _zz_90;
      end
      if(_zz_41)begin
        img_reg_array_39_12_real <= _zz_90;
      end
      if(_zz_42)begin
        img_reg_array_40_12_real <= _zz_90;
      end
      if(_zz_43)begin
        img_reg_array_41_12_real <= _zz_90;
      end
      if(_zz_44)begin
        img_reg_array_42_12_real <= _zz_90;
      end
      if(_zz_45)begin
        img_reg_array_43_12_real <= _zz_90;
      end
      if(_zz_46)begin
        img_reg_array_44_12_real <= _zz_90;
      end
      if(_zz_47)begin
        img_reg_array_45_12_real <= _zz_90;
      end
      if(_zz_48)begin
        img_reg_array_46_12_real <= _zz_90;
      end
      if(_zz_49)begin
        img_reg_array_47_12_real <= _zz_90;
      end
      if(_zz_50)begin
        img_reg_array_48_12_real <= _zz_90;
      end
      if(_zz_51)begin
        img_reg_array_49_12_real <= _zz_90;
      end
      if(_zz_52)begin
        img_reg_array_50_12_real <= _zz_90;
      end
      if(_zz_53)begin
        img_reg_array_51_12_real <= _zz_90;
      end
      if(_zz_54)begin
        img_reg_array_52_12_real <= _zz_90;
      end
      if(_zz_55)begin
        img_reg_array_53_12_real <= _zz_90;
      end
      if(_zz_56)begin
        img_reg_array_54_12_real <= _zz_90;
      end
      if(_zz_57)begin
        img_reg_array_55_12_real <= _zz_90;
      end
      if(_zz_58)begin
        img_reg_array_56_12_real <= _zz_90;
      end
      if(_zz_59)begin
        img_reg_array_57_12_real <= _zz_90;
      end
      if(_zz_60)begin
        img_reg_array_58_12_real <= _zz_90;
      end
      if(_zz_61)begin
        img_reg_array_59_12_real <= _zz_90;
      end
      if(_zz_62)begin
        img_reg_array_60_12_real <= _zz_90;
      end
      if(_zz_63)begin
        img_reg_array_61_12_real <= _zz_90;
      end
      if(_zz_64)begin
        img_reg_array_62_12_real <= _zz_90;
      end
      if(_zz_65)begin
        img_reg_array_63_12_real <= _zz_90;
      end
      if(_zz_2)begin
        img_reg_array_0_12_imag <= _zz_91;
      end
      if(_zz_3)begin
        img_reg_array_1_12_imag <= _zz_91;
      end
      if(_zz_4)begin
        img_reg_array_2_12_imag <= _zz_91;
      end
      if(_zz_5)begin
        img_reg_array_3_12_imag <= _zz_91;
      end
      if(_zz_6)begin
        img_reg_array_4_12_imag <= _zz_91;
      end
      if(_zz_7)begin
        img_reg_array_5_12_imag <= _zz_91;
      end
      if(_zz_8)begin
        img_reg_array_6_12_imag <= _zz_91;
      end
      if(_zz_9)begin
        img_reg_array_7_12_imag <= _zz_91;
      end
      if(_zz_10)begin
        img_reg_array_8_12_imag <= _zz_91;
      end
      if(_zz_11)begin
        img_reg_array_9_12_imag <= _zz_91;
      end
      if(_zz_12)begin
        img_reg_array_10_12_imag <= _zz_91;
      end
      if(_zz_13)begin
        img_reg_array_11_12_imag <= _zz_91;
      end
      if(_zz_14)begin
        img_reg_array_12_12_imag <= _zz_91;
      end
      if(_zz_15)begin
        img_reg_array_13_12_imag <= _zz_91;
      end
      if(_zz_16)begin
        img_reg_array_14_12_imag <= _zz_91;
      end
      if(_zz_17)begin
        img_reg_array_15_12_imag <= _zz_91;
      end
      if(_zz_18)begin
        img_reg_array_16_12_imag <= _zz_91;
      end
      if(_zz_19)begin
        img_reg_array_17_12_imag <= _zz_91;
      end
      if(_zz_20)begin
        img_reg_array_18_12_imag <= _zz_91;
      end
      if(_zz_21)begin
        img_reg_array_19_12_imag <= _zz_91;
      end
      if(_zz_22)begin
        img_reg_array_20_12_imag <= _zz_91;
      end
      if(_zz_23)begin
        img_reg_array_21_12_imag <= _zz_91;
      end
      if(_zz_24)begin
        img_reg_array_22_12_imag <= _zz_91;
      end
      if(_zz_25)begin
        img_reg_array_23_12_imag <= _zz_91;
      end
      if(_zz_26)begin
        img_reg_array_24_12_imag <= _zz_91;
      end
      if(_zz_27)begin
        img_reg_array_25_12_imag <= _zz_91;
      end
      if(_zz_28)begin
        img_reg_array_26_12_imag <= _zz_91;
      end
      if(_zz_29)begin
        img_reg_array_27_12_imag <= _zz_91;
      end
      if(_zz_30)begin
        img_reg_array_28_12_imag <= _zz_91;
      end
      if(_zz_31)begin
        img_reg_array_29_12_imag <= _zz_91;
      end
      if(_zz_32)begin
        img_reg_array_30_12_imag <= _zz_91;
      end
      if(_zz_33)begin
        img_reg_array_31_12_imag <= _zz_91;
      end
      if(_zz_34)begin
        img_reg_array_32_12_imag <= _zz_91;
      end
      if(_zz_35)begin
        img_reg_array_33_12_imag <= _zz_91;
      end
      if(_zz_36)begin
        img_reg_array_34_12_imag <= _zz_91;
      end
      if(_zz_37)begin
        img_reg_array_35_12_imag <= _zz_91;
      end
      if(_zz_38)begin
        img_reg_array_36_12_imag <= _zz_91;
      end
      if(_zz_39)begin
        img_reg_array_37_12_imag <= _zz_91;
      end
      if(_zz_40)begin
        img_reg_array_38_12_imag <= _zz_91;
      end
      if(_zz_41)begin
        img_reg_array_39_12_imag <= _zz_91;
      end
      if(_zz_42)begin
        img_reg_array_40_12_imag <= _zz_91;
      end
      if(_zz_43)begin
        img_reg_array_41_12_imag <= _zz_91;
      end
      if(_zz_44)begin
        img_reg_array_42_12_imag <= _zz_91;
      end
      if(_zz_45)begin
        img_reg_array_43_12_imag <= _zz_91;
      end
      if(_zz_46)begin
        img_reg_array_44_12_imag <= _zz_91;
      end
      if(_zz_47)begin
        img_reg_array_45_12_imag <= _zz_91;
      end
      if(_zz_48)begin
        img_reg_array_46_12_imag <= _zz_91;
      end
      if(_zz_49)begin
        img_reg_array_47_12_imag <= _zz_91;
      end
      if(_zz_50)begin
        img_reg_array_48_12_imag <= _zz_91;
      end
      if(_zz_51)begin
        img_reg_array_49_12_imag <= _zz_91;
      end
      if(_zz_52)begin
        img_reg_array_50_12_imag <= _zz_91;
      end
      if(_zz_53)begin
        img_reg_array_51_12_imag <= _zz_91;
      end
      if(_zz_54)begin
        img_reg_array_52_12_imag <= _zz_91;
      end
      if(_zz_55)begin
        img_reg_array_53_12_imag <= _zz_91;
      end
      if(_zz_56)begin
        img_reg_array_54_12_imag <= _zz_91;
      end
      if(_zz_57)begin
        img_reg_array_55_12_imag <= _zz_91;
      end
      if(_zz_58)begin
        img_reg_array_56_12_imag <= _zz_91;
      end
      if(_zz_59)begin
        img_reg_array_57_12_imag <= _zz_91;
      end
      if(_zz_60)begin
        img_reg_array_58_12_imag <= _zz_91;
      end
      if(_zz_61)begin
        img_reg_array_59_12_imag <= _zz_91;
      end
      if(_zz_62)begin
        img_reg_array_60_12_imag <= _zz_91;
      end
      if(_zz_63)begin
        img_reg_array_61_12_imag <= _zz_91;
      end
      if(_zz_64)begin
        img_reg_array_62_12_imag <= _zz_91;
      end
      if(_zz_65)begin
        img_reg_array_63_12_imag <= _zz_91;
      end
      if(_zz_2)begin
        img_reg_array_0_13_real <= _zz_92;
      end
      if(_zz_3)begin
        img_reg_array_1_13_real <= _zz_92;
      end
      if(_zz_4)begin
        img_reg_array_2_13_real <= _zz_92;
      end
      if(_zz_5)begin
        img_reg_array_3_13_real <= _zz_92;
      end
      if(_zz_6)begin
        img_reg_array_4_13_real <= _zz_92;
      end
      if(_zz_7)begin
        img_reg_array_5_13_real <= _zz_92;
      end
      if(_zz_8)begin
        img_reg_array_6_13_real <= _zz_92;
      end
      if(_zz_9)begin
        img_reg_array_7_13_real <= _zz_92;
      end
      if(_zz_10)begin
        img_reg_array_8_13_real <= _zz_92;
      end
      if(_zz_11)begin
        img_reg_array_9_13_real <= _zz_92;
      end
      if(_zz_12)begin
        img_reg_array_10_13_real <= _zz_92;
      end
      if(_zz_13)begin
        img_reg_array_11_13_real <= _zz_92;
      end
      if(_zz_14)begin
        img_reg_array_12_13_real <= _zz_92;
      end
      if(_zz_15)begin
        img_reg_array_13_13_real <= _zz_92;
      end
      if(_zz_16)begin
        img_reg_array_14_13_real <= _zz_92;
      end
      if(_zz_17)begin
        img_reg_array_15_13_real <= _zz_92;
      end
      if(_zz_18)begin
        img_reg_array_16_13_real <= _zz_92;
      end
      if(_zz_19)begin
        img_reg_array_17_13_real <= _zz_92;
      end
      if(_zz_20)begin
        img_reg_array_18_13_real <= _zz_92;
      end
      if(_zz_21)begin
        img_reg_array_19_13_real <= _zz_92;
      end
      if(_zz_22)begin
        img_reg_array_20_13_real <= _zz_92;
      end
      if(_zz_23)begin
        img_reg_array_21_13_real <= _zz_92;
      end
      if(_zz_24)begin
        img_reg_array_22_13_real <= _zz_92;
      end
      if(_zz_25)begin
        img_reg_array_23_13_real <= _zz_92;
      end
      if(_zz_26)begin
        img_reg_array_24_13_real <= _zz_92;
      end
      if(_zz_27)begin
        img_reg_array_25_13_real <= _zz_92;
      end
      if(_zz_28)begin
        img_reg_array_26_13_real <= _zz_92;
      end
      if(_zz_29)begin
        img_reg_array_27_13_real <= _zz_92;
      end
      if(_zz_30)begin
        img_reg_array_28_13_real <= _zz_92;
      end
      if(_zz_31)begin
        img_reg_array_29_13_real <= _zz_92;
      end
      if(_zz_32)begin
        img_reg_array_30_13_real <= _zz_92;
      end
      if(_zz_33)begin
        img_reg_array_31_13_real <= _zz_92;
      end
      if(_zz_34)begin
        img_reg_array_32_13_real <= _zz_92;
      end
      if(_zz_35)begin
        img_reg_array_33_13_real <= _zz_92;
      end
      if(_zz_36)begin
        img_reg_array_34_13_real <= _zz_92;
      end
      if(_zz_37)begin
        img_reg_array_35_13_real <= _zz_92;
      end
      if(_zz_38)begin
        img_reg_array_36_13_real <= _zz_92;
      end
      if(_zz_39)begin
        img_reg_array_37_13_real <= _zz_92;
      end
      if(_zz_40)begin
        img_reg_array_38_13_real <= _zz_92;
      end
      if(_zz_41)begin
        img_reg_array_39_13_real <= _zz_92;
      end
      if(_zz_42)begin
        img_reg_array_40_13_real <= _zz_92;
      end
      if(_zz_43)begin
        img_reg_array_41_13_real <= _zz_92;
      end
      if(_zz_44)begin
        img_reg_array_42_13_real <= _zz_92;
      end
      if(_zz_45)begin
        img_reg_array_43_13_real <= _zz_92;
      end
      if(_zz_46)begin
        img_reg_array_44_13_real <= _zz_92;
      end
      if(_zz_47)begin
        img_reg_array_45_13_real <= _zz_92;
      end
      if(_zz_48)begin
        img_reg_array_46_13_real <= _zz_92;
      end
      if(_zz_49)begin
        img_reg_array_47_13_real <= _zz_92;
      end
      if(_zz_50)begin
        img_reg_array_48_13_real <= _zz_92;
      end
      if(_zz_51)begin
        img_reg_array_49_13_real <= _zz_92;
      end
      if(_zz_52)begin
        img_reg_array_50_13_real <= _zz_92;
      end
      if(_zz_53)begin
        img_reg_array_51_13_real <= _zz_92;
      end
      if(_zz_54)begin
        img_reg_array_52_13_real <= _zz_92;
      end
      if(_zz_55)begin
        img_reg_array_53_13_real <= _zz_92;
      end
      if(_zz_56)begin
        img_reg_array_54_13_real <= _zz_92;
      end
      if(_zz_57)begin
        img_reg_array_55_13_real <= _zz_92;
      end
      if(_zz_58)begin
        img_reg_array_56_13_real <= _zz_92;
      end
      if(_zz_59)begin
        img_reg_array_57_13_real <= _zz_92;
      end
      if(_zz_60)begin
        img_reg_array_58_13_real <= _zz_92;
      end
      if(_zz_61)begin
        img_reg_array_59_13_real <= _zz_92;
      end
      if(_zz_62)begin
        img_reg_array_60_13_real <= _zz_92;
      end
      if(_zz_63)begin
        img_reg_array_61_13_real <= _zz_92;
      end
      if(_zz_64)begin
        img_reg_array_62_13_real <= _zz_92;
      end
      if(_zz_65)begin
        img_reg_array_63_13_real <= _zz_92;
      end
      if(_zz_2)begin
        img_reg_array_0_13_imag <= _zz_93;
      end
      if(_zz_3)begin
        img_reg_array_1_13_imag <= _zz_93;
      end
      if(_zz_4)begin
        img_reg_array_2_13_imag <= _zz_93;
      end
      if(_zz_5)begin
        img_reg_array_3_13_imag <= _zz_93;
      end
      if(_zz_6)begin
        img_reg_array_4_13_imag <= _zz_93;
      end
      if(_zz_7)begin
        img_reg_array_5_13_imag <= _zz_93;
      end
      if(_zz_8)begin
        img_reg_array_6_13_imag <= _zz_93;
      end
      if(_zz_9)begin
        img_reg_array_7_13_imag <= _zz_93;
      end
      if(_zz_10)begin
        img_reg_array_8_13_imag <= _zz_93;
      end
      if(_zz_11)begin
        img_reg_array_9_13_imag <= _zz_93;
      end
      if(_zz_12)begin
        img_reg_array_10_13_imag <= _zz_93;
      end
      if(_zz_13)begin
        img_reg_array_11_13_imag <= _zz_93;
      end
      if(_zz_14)begin
        img_reg_array_12_13_imag <= _zz_93;
      end
      if(_zz_15)begin
        img_reg_array_13_13_imag <= _zz_93;
      end
      if(_zz_16)begin
        img_reg_array_14_13_imag <= _zz_93;
      end
      if(_zz_17)begin
        img_reg_array_15_13_imag <= _zz_93;
      end
      if(_zz_18)begin
        img_reg_array_16_13_imag <= _zz_93;
      end
      if(_zz_19)begin
        img_reg_array_17_13_imag <= _zz_93;
      end
      if(_zz_20)begin
        img_reg_array_18_13_imag <= _zz_93;
      end
      if(_zz_21)begin
        img_reg_array_19_13_imag <= _zz_93;
      end
      if(_zz_22)begin
        img_reg_array_20_13_imag <= _zz_93;
      end
      if(_zz_23)begin
        img_reg_array_21_13_imag <= _zz_93;
      end
      if(_zz_24)begin
        img_reg_array_22_13_imag <= _zz_93;
      end
      if(_zz_25)begin
        img_reg_array_23_13_imag <= _zz_93;
      end
      if(_zz_26)begin
        img_reg_array_24_13_imag <= _zz_93;
      end
      if(_zz_27)begin
        img_reg_array_25_13_imag <= _zz_93;
      end
      if(_zz_28)begin
        img_reg_array_26_13_imag <= _zz_93;
      end
      if(_zz_29)begin
        img_reg_array_27_13_imag <= _zz_93;
      end
      if(_zz_30)begin
        img_reg_array_28_13_imag <= _zz_93;
      end
      if(_zz_31)begin
        img_reg_array_29_13_imag <= _zz_93;
      end
      if(_zz_32)begin
        img_reg_array_30_13_imag <= _zz_93;
      end
      if(_zz_33)begin
        img_reg_array_31_13_imag <= _zz_93;
      end
      if(_zz_34)begin
        img_reg_array_32_13_imag <= _zz_93;
      end
      if(_zz_35)begin
        img_reg_array_33_13_imag <= _zz_93;
      end
      if(_zz_36)begin
        img_reg_array_34_13_imag <= _zz_93;
      end
      if(_zz_37)begin
        img_reg_array_35_13_imag <= _zz_93;
      end
      if(_zz_38)begin
        img_reg_array_36_13_imag <= _zz_93;
      end
      if(_zz_39)begin
        img_reg_array_37_13_imag <= _zz_93;
      end
      if(_zz_40)begin
        img_reg_array_38_13_imag <= _zz_93;
      end
      if(_zz_41)begin
        img_reg_array_39_13_imag <= _zz_93;
      end
      if(_zz_42)begin
        img_reg_array_40_13_imag <= _zz_93;
      end
      if(_zz_43)begin
        img_reg_array_41_13_imag <= _zz_93;
      end
      if(_zz_44)begin
        img_reg_array_42_13_imag <= _zz_93;
      end
      if(_zz_45)begin
        img_reg_array_43_13_imag <= _zz_93;
      end
      if(_zz_46)begin
        img_reg_array_44_13_imag <= _zz_93;
      end
      if(_zz_47)begin
        img_reg_array_45_13_imag <= _zz_93;
      end
      if(_zz_48)begin
        img_reg_array_46_13_imag <= _zz_93;
      end
      if(_zz_49)begin
        img_reg_array_47_13_imag <= _zz_93;
      end
      if(_zz_50)begin
        img_reg_array_48_13_imag <= _zz_93;
      end
      if(_zz_51)begin
        img_reg_array_49_13_imag <= _zz_93;
      end
      if(_zz_52)begin
        img_reg_array_50_13_imag <= _zz_93;
      end
      if(_zz_53)begin
        img_reg_array_51_13_imag <= _zz_93;
      end
      if(_zz_54)begin
        img_reg_array_52_13_imag <= _zz_93;
      end
      if(_zz_55)begin
        img_reg_array_53_13_imag <= _zz_93;
      end
      if(_zz_56)begin
        img_reg_array_54_13_imag <= _zz_93;
      end
      if(_zz_57)begin
        img_reg_array_55_13_imag <= _zz_93;
      end
      if(_zz_58)begin
        img_reg_array_56_13_imag <= _zz_93;
      end
      if(_zz_59)begin
        img_reg_array_57_13_imag <= _zz_93;
      end
      if(_zz_60)begin
        img_reg_array_58_13_imag <= _zz_93;
      end
      if(_zz_61)begin
        img_reg_array_59_13_imag <= _zz_93;
      end
      if(_zz_62)begin
        img_reg_array_60_13_imag <= _zz_93;
      end
      if(_zz_63)begin
        img_reg_array_61_13_imag <= _zz_93;
      end
      if(_zz_64)begin
        img_reg_array_62_13_imag <= _zz_93;
      end
      if(_zz_65)begin
        img_reg_array_63_13_imag <= _zz_93;
      end
      if(_zz_2)begin
        img_reg_array_0_14_real <= _zz_94;
      end
      if(_zz_3)begin
        img_reg_array_1_14_real <= _zz_94;
      end
      if(_zz_4)begin
        img_reg_array_2_14_real <= _zz_94;
      end
      if(_zz_5)begin
        img_reg_array_3_14_real <= _zz_94;
      end
      if(_zz_6)begin
        img_reg_array_4_14_real <= _zz_94;
      end
      if(_zz_7)begin
        img_reg_array_5_14_real <= _zz_94;
      end
      if(_zz_8)begin
        img_reg_array_6_14_real <= _zz_94;
      end
      if(_zz_9)begin
        img_reg_array_7_14_real <= _zz_94;
      end
      if(_zz_10)begin
        img_reg_array_8_14_real <= _zz_94;
      end
      if(_zz_11)begin
        img_reg_array_9_14_real <= _zz_94;
      end
      if(_zz_12)begin
        img_reg_array_10_14_real <= _zz_94;
      end
      if(_zz_13)begin
        img_reg_array_11_14_real <= _zz_94;
      end
      if(_zz_14)begin
        img_reg_array_12_14_real <= _zz_94;
      end
      if(_zz_15)begin
        img_reg_array_13_14_real <= _zz_94;
      end
      if(_zz_16)begin
        img_reg_array_14_14_real <= _zz_94;
      end
      if(_zz_17)begin
        img_reg_array_15_14_real <= _zz_94;
      end
      if(_zz_18)begin
        img_reg_array_16_14_real <= _zz_94;
      end
      if(_zz_19)begin
        img_reg_array_17_14_real <= _zz_94;
      end
      if(_zz_20)begin
        img_reg_array_18_14_real <= _zz_94;
      end
      if(_zz_21)begin
        img_reg_array_19_14_real <= _zz_94;
      end
      if(_zz_22)begin
        img_reg_array_20_14_real <= _zz_94;
      end
      if(_zz_23)begin
        img_reg_array_21_14_real <= _zz_94;
      end
      if(_zz_24)begin
        img_reg_array_22_14_real <= _zz_94;
      end
      if(_zz_25)begin
        img_reg_array_23_14_real <= _zz_94;
      end
      if(_zz_26)begin
        img_reg_array_24_14_real <= _zz_94;
      end
      if(_zz_27)begin
        img_reg_array_25_14_real <= _zz_94;
      end
      if(_zz_28)begin
        img_reg_array_26_14_real <= _zz_94;
      end
      if(_zz_29)begin
        img_reg_array_27_14_real <= _zz_94;
      end
      if(_zz_30)begin
        img_reg_array_28_14_real <= _zz_94;
      end
      if(_zz_31)begin
        img_reg_array_29_14_real <= _zz_94;
      end
      if(_zz_32)begin
        img_reg_array_30_14_real <= _zz_94;
      end
      if(_zz_33)begin
        img_reg_array_31_14_real <= _zz_94;
      end
      if(_zz_34)begin
        img_reg_array_32_14_real <= _zz_94;
      end
      if(_zz_35)begin
        img_reg_array_33_14_real <= _zz_94;
      end
      if(_zz_36)begin
        img_reg_array_34_14_real <= _zz_94;
      end
      if(_zz_37)begin
        img_reg_array_35_14_real <= _zz_94;
      end
      if(_zz_38)begin
        img_reg_array_36_14_real <= _zz_94;
      end
      if(_zz_39)begin
        img_reg_array_37_14_real <= _zz_94;
      end
      if(_zz_40)begin
        img_reg_array_38_14_real <= _zz_94;
      end
      if(_zz_41)begin
        img_reg_array_39_14_real <= _zz_94;
      end
      if(_zz_42)begin
        img_reg_array_40_14_real <= _zz_94;
      end
      if(_zz_43)begin
        img_reg_array_41_14_real <= _zz_94;
      end
      if(_zz_44)begin
        img_reg_array_42_14_real <= _zz_94;
      end
      if(_zz_45)begin
        img_reg_array_43_14_real <= _zz_94;
      end
      if(_zz_46)begin
        img_reg_array_44_14_real <= _zz_94;
      end
      if(_zz_47)begin
        img_reg_array_45_14_real <= _zz_94;
      end
      if(_zz_48)begin
        img_reg_array_46_14_real <= _zz_94;
      end
      if(_zz_49)begin
        img_reg_array_47_14_real <= _zz_94;
      end
      if(_zz_50)begin
        img_reg_array_48_14_real <= _zz_94;
      end
      if(_zz_51)begin
        img_reg_array_49_14_real <= _zz_94;
      end
      if(_zz_52)begin
        img_reg_array_50_14_real <= _zz_94;
      end
      if(_zz_53)begin
        img_reg_array_51_14_real <= _zz_94;
      end
      if(_zz_54)begin
        img_reg_array_52_14_real <= _zz_94;
      end
      if(_zz_55)begin
        img_reg_array_53_14_real <= _zz_94;
      end
      if(_zz_56)begin
        img_reg_array_54_14_real <= _zz_94;
      end
      if(_zz_57)begin
        img_reg_array_55_14_real <= _zz_94;
      end
      if(_zz_58)begin
        img_reg_array_56_14_real <= _zz_94;
      end
      if(_zz_59)begin
        img_reg_array_57_14_real <= _zz_94;
      end
      if(_zz_60)begin
        img_reg_array_58_14_real <= _zz_94;
      end
      if(_zz_61)begin
        img_reg_array_59_14_real <= _zz_94;
      end
      if(_zz_62)begin
        img_reg_array_60_14_real <= _zz_94;
      end
      if(_zz_63)begin
        img_reg_array_61_14_real <= _zz_94;
      end
      if(_zz_64)begin
        img_reg_array_62_14_real <= _zz_94;
      end
      if(_zz_65)begin
        img_reg_array_63_14_real <= _zz_94;
      end
      if(_zz_2)begin
        img_reg_array_0_14_imag <= _zz_95;
      end
      if(_zz_3)begin
        img_reg_array_1_14_imag <= _zz_95;
      end
      if(_zz_4)begin
        img_reg_array_2_14_imag <= _zz_95;
      end
      if(_zz_5)begin
        img_reg_array_3_14_imag <= _zz_95;
      end
      if(_zz_6)begin
        img_reg_array_4_14_imag <= _zz_95;
      end
      if(_zz_7)begin
        img_reg_array_5_14_imag <= _zz_95;
      end
      if(_zz_8)begin
        img_reg_array_6_14_imag <= _zz_95;
      end
      if(_zz_9)begin
        img_reg_array_7_14_imag <= _zz_95;
      end
      if(_zz_10)begin
        img_reg_array_8_14_imag <= _zz_95;
      end
      if(_zz_11)begin
        img_reg_array_9_14_imag <= _zz_95;
      end
      if(_zz_12)begin
        img_reg_array_10_14_imag <= _zz_95;
      end
      if(_zz_13)begin
        img_reg_array_11_14_imag <= _zz_95;
      end
      if(_zz_14)begin
        img_reg_array_12_14_imag <= _zz_95;
      end
      if(_zz_15)begin
        img_reg_array_13_14_imag <= _zz_95;
      end
      if(_zz_16)begin
        img_reg_array_14_14_imag <= _zz_95;
      end
      if(_zz_17)begin
        img_reg_array_15_14_imag <= _zz_95;
      end
      if(_zz_18)begin
        img_reg_array_16_14_imag <= _zz_95;
      end
      if(_zz_19)begin
        img_reg_array_17_14_imag <= _zz_95;
      end
      if(_zz_20)begin
        img_reg_array_18_14_imag <= _zz_95;
      end
      if(_zz_21)begin
        img_reg_array_19_14_imag <= _zz_95;
      end
      if(_zz_22)begin
        img_reg_array_20_14_imag <= _zz_95;
      end
      if(_zz_23)begin
        img_reg_array_21_14_imag <= _zz_95;
      end
      if(_zz_24)begin
        img_reg_array_22_14_imag <= _zz_95;
      end
      if(_zz_25)begin
        img_reg_array_23_14_imag <= _zz_95;
      end
      if(_zz_26)begin
        img_reg_array_24_14_imag <= _zz_95;
      end
      if(_zz_27)begin
        img_reg_array_25_14_imag <= _zz_95;
      end
      if(_zz_28)begin
        img_reg_array_26_14_imag <= _zz_95;
      end
      if(_zz_29)begin
        img_reg_array_27_14_imag <= _zz_95;
      end
      if(_zz_30)begin
        img_reg_array_28_14_imag <= _zz_95;
      end
      if(_zz_31)begin
        img_reg_array_29_14_imag <= _zz_95;
      end
      if(_zz_32)begin
        img_reg_array_30_14_imag <= _zz_95;
      end
      if(_zz_33)begin
        img_reg_array_31_14_imag <= _zz_95;
      end
      if(_zz_34)begin
        img_reg_array_32_14_imag <= _zz_95;
      end
      if(_zz_35)begin
        img_reg_array_33_14_imag <= _zz_95;
      end
      if(_zz_36)begin
        img_reg_array_34_14_imag <= _zz_95;
      end
      if(_zz_37)begin
        img_reg_array_35_14_imag <= _zz_95;
      end
      if(_zz_38)begin
        img_reg_array_36_14_imag <= _zz_95;
      end
      if(_zz_39)begin
        img_reg_array_37_14_imag <= _zz_95;
      end
      if(_zz_40)begin
        img_reg_array_38_14_imag <= _zz_95;
      end
      if(_zz_41)begin
        img_reg_array_39_14_imag <= _zz_95;
      end
      if(_zz_42)begin
        img_reg_array_40_14_imag <= _zz_95;
      end
      if(_zz_43)begin
        img_reg_array_41_14_imag <= _zz_95;
      end
      if(_zz_44)begin
        img_reg_array_42_14_imag <= _zz_95;
      end
      if(_zz_45)begin
        img_reg_array_43_14_imag <= _zz_95;
      end
      if(_zz_46)begin
        img_reg_array_44_14_imag <= _zz_95;
      end
      if(_zz_47)begin
        img_reg_array_45_14_imag <= _zz_95;
      end
      if(_zz_48)begin
        img_reg_array_46_14_imag <= _zz_95;
      end
      if(_zz_49)begin
        img_reg_array_47_14_imag <= _zz_95;
      end
      if(_zz_50)begin
        img_reg_array_48_14_imag <= _zz_95;
      end
      if(_zz_51)begin
        img_reg_array_49_14_imag <= _zz_95;
      end
      if(_zz_52)begin
        img_reg_array_50_14_imag <= _zz_95;
      end
      if(_zz_53)begin
        img_reg_array_51_14_imag <= _zz_95;
      end
      if(_zz_54)begin
        img_reg_array_52_14_imag <= _zz_95;
      end
      if(_zz_55)begin
        img_reg_array_53_14_imag <= _zz_95;
      end
      if(_zz_56)begin
        img_reg_array_54_14_imag <= _zz_95;
      end
      if(_zz_57)begin
        img_reg_array_55_14_imag <= _zz_95;
      end
      if(_zz_58)begin
        img_reg_array_56_14_imag <= _zz_95;
      end
      if(_zz_59)begin
        img_reg_array_57_14_imag <= _zz_95;
      end
      if(_zz_60)begin
        img_reg_array_58_14_imag <= _zz_95;
      end
      if(_zz_61)begin
        img_reg_array_59_14_imag <= _zz_95;
      end
      if(_zz_62)begin
        img_reg_array_60_14_imag <= _zz_95;
      end
      if(_zz_63)begin
        img_reg_array_61_14_imag <= _zz_95;
      end
      if(_zz_64)begin
        img_reg_array_62_14_imag <= _zz_95;
      end
      if(_zz_65)begin
        img_reg_array_63_14_imag <= _zz_95;
      end
      if(_zz_2)begin
        img_reg_array_0_15_real <= _zz_96;
      end
      if(_zz_3)begin
        img_reg_array_1_15_real <= _zz_96;
      end
      if(_zz_4)begin
        img_reg_array_2_15_real <= _zz_96;
      end
      if(_zz_5)begin
        img_reg_array_3_15_real <= _zz_96;
      end
      if(_zz_6)begin
        img_reg_array_4_15_real <= _zz_96;
      end
      if(_zz_7)begin
        img_reg_array_5_15_real <= _zz_96;
      end
      if(_zz_8)begin
        img_reg_array_6_15_real <= _zz_96;
      end
      if(_zz_9)begin
        img_reg_array_7_15_real <= _zz_96;
      end
      if(_zz_10)begin
        img_reg_array_8_15_real <= _zz_96;
      end
      if(_zz_11)begin
        img_reg_array_9_15_real <= _zz_96;
      end
      if(_zz_12)begin
        img_reg_array_10_15_real <= _zz_96;
      end
      if(_zz_13)begin
        img_reg_array_11_15_real <= _zz_96;
      end
      if(_zz_14)begin
        img_reg_array_12_15_real <= _zz_96;
      end
      if(_zz_15)begin
        img_reg_array_13_15_real <= _zz_96;
      end
      if(_zz_16)begin
        img_reg_array_14_15_real <= _zz_96;
      end
      if(_zz_17)begin
        img_reg_array_15_15_real <= _zz_96;
      end
      if(_zz_18)begin
        img_reg_array_16_15_real <= _zz_96;
      end
      if(_zz_19)begin
        img_reg_array_17_15_real <= _zz_96;
      end
      if(_zz_20)begin
        img_reg_array_18_15_real <= _zz_96;
      end
      if(_zz_21)begin
        img_reg_array_19_15_real <= _zz_96;
      end
      if(_zz_22)begin
        img_reg_array_20_15_real <= _zz_96;
      end
      if(_zz_23)begin
        img_reg_array_21_15_real <= _zz_96;
      end
      if(_zz_24)begin
        img_reg_array_22_15_real <= _zz_96;
      end
      if(_zz_25)begin
        img_reg_array_23_15_real <= _zz_96;
      end
      if(_zz_26)begin
        img_reg_array_24_15_real <= _zz_96;
      end
      if(_zz_27)begin
        img_reg_array_25_15_real <= _zz_96;
      end
      if(_zz_28)begin
        img_reg_array_26_15_real <= _zz_96;
      end
      if(_zz_29)begin
        img_reg_array_27_15_real <= _zz_96;
      end
      if(_zz_30)begin
        img_reg_array_28_15_real <= _zz_96;
      end
      if(_zz_31)begin
        img_reg_array_29_15_real <= _zz_96;
      end
      if(_zz_32)begin
        img_reg_array_30_15_real <= _zz_96;
      end
      if(_zz_33)begin
        img_reg_array_31_15_real <= _zz_96;
      end
      if(_zz_34)begin
        img_reg_array_32_15_real <= _zz_96;
      end
      if(_zz_35)begin
        img_reg_array_33_15_real <= _zz_96;
      end
      if(_zz_36)begin
        img_reg_array_34_15_real <= _zz_96;
      end
      if(_zz_37)begin
        img_reg_array_35_15_real <= _zz_96;
      end
      if(_zz_38)begin
        img_reg_array_36_15_real <= _zz_96;
      end
      if(_zz_39)begin
        img_reg_array_37_15_real <= _zz_96;
      end
      if(_zz_40)begin
        img_reg_array_38_15_real <= _zz_96;
      end
      if(_zz_41)begin
        img_reg_array_39_15_real <= _zz_96;
      end
      if(_zz_42)begin
        img_reg_array_40_15_real <= _zz_96;
      end
      if(_zz_43)begin
        img_reg_array_41_15_real <= _zz_96;
      end
      if(_zz_44)begin
        img_reg_array_42_15_real <= _zz_96;
      end
      if(_zz_45)begin
        img_reg_array_43_15_real <= _zz_96;
      end
      if(_zz_46)begin
        img_reg_array_44_15_real <= _zz_96;
      end
      if(_zz_47)begin
        img_reg_array_45_15_real <= _zz_96;
      end
      if(_zz_48)begin
        img_reg_array_46_15_real <= _zz_96;
      end
      if(_zz_49)begin
        img_reg_array_47_15_real <= _zz_96;
      end
      if(_zz_50)begin
        img_reg_array_48_15_real <= _zz_96;
      end
      if(_zz_51)begin
        img_reg_array_49_15_real <= _zz_96;
      end
      if(_zz_52)begin
        img_reg_array_50_15_real <= _zz_96;
      end
      if(_zz_53)begin
        img_reg_array_51_15_real <= _zz_96;
      end
      if(_zz_54)begin
        img_reg_array_52_15_real <= _zz_96;
      end
      if(_zz_55)begin
        img_reg_array_53_15_real <= _zz_96;
      end
      if(_zz_56)begin
        img_reg_array_54_15_real <= _zz_96;
      end
      if(_zz_57)begin
        img_reg_array_55_15_real <= _zz_96;
      end
      if(_zz_58)begin
        img_reg_array_56_15_real <= _zz_96;
      end
      if(_zz_59)begin
        img_reg_array_57_15_real <= _zz_96;
      end
      if(_zz_60)begin
        img_reg_array_58_15_real <= _zz_96;
      end
      if(_zz_61)begin
        img_reg_array_59_15_real <= _zz_96;
      end
      if(_zz_62)begin
        img_reg_array_60_15_real <= _zz_96;
      end
      if(_zz_63)begin
        img_reg_array_61_15_real <= _zz_96;
      end
      if(_zz_64)begin
        img_reg_array_62_15_real <= _zz_96;
      end
      if(_zz_65)begin
        img_reg_array_63_15_real <= _zz_96;
      end
      if(_zz_2)begin
        img_reg_array_0_15_imag <= _zz_97;
      end
      if(_zz_3)begin
        img_reg_array_1_15_imag <= _zz_97;
      end
      if(_zz_4)begin
        img_reg_array_2_15_imag <= _zz_97;
      end
      if(_zz_5)begin
        img_reg_array_3_15_imag <= _zz_97;
      end
      if(_zz_6)begin
        img_reg_array_4_15_imag <= _zz_97;
      end
      if(_zz_7)begin
        img_reg_array_5_15_imag <= _zz_97;
      end
      if(_zz_8)begin
        img_reg_array_6_15_imag <= _zz_97;
      end
      if(_zz_9)begin
        img_reg_array_7_15_imag <= _zz_97;
      end
      if(_zz_10)begin
        img_reg_array_8_15_imag <= _zz_97;
      end
      if(_zz_11)begin
        img_reg_array_9_15_imag <= _zz_97;
      end
      if(_zz_12)begin
        img_reg_array_10_15_imag <= _zz_97;
      end
      if(_zz_13)begin
        img_reg_array_11_15_imag <= _zz_97;
      end
      if(_zz_14)begin
        img_reg_array_12_15_imag <= _zz_97;
      end
      if(_zz_15)begin
        img_reg_array_13_15_imag <= _zz_97;
      end
      if(_zz_16)begin
        img_reg_array_14_15_imag <= _zz_97;
      end
      if(_zz_17)begin
        img_reg_array_15_15_imag <= _zz_97;
      end
      if(_zz_18)begin
        img_reg_array_16_15_imag <= _zz_97;
      end
      if(_zz_19)begin
        img_reg_array_17_15_imag <= _zz_97;
      end
      if(_zz_20)begin
        img_reg_array_18_15_imag <= _zz_97;
      end
      if(_zz_21)begin
        img_reg_array_19_15_imag <= _zz_97;
      end
      if(_zz_22)begin
        img_reg_array_20_15_imag <= _zz_97;
      end
      if(_zz_23)begin
        img_reg_array_21_15_imag <= _zz_97;
      end
      if(_zz_24)begin
        img_reg_array_22_15_imag <= _zz_97;
      end
      if(_zz_25)begin
        img_reg_array_23_15_imag <= _zz_97;
      end
      if(_zz_26)begin
        img_reg_array_24_15_imag <= _zz_97;
      end
      if(_zz_27)begin
        img_reg_array_25_15_imag <= _zz_97;
      end
      if(_zz_28)begin
        img_reg_array_26_15_imag <= _zz_97;
      end
      if(_zz_29)begin
        img_reg_array_27_15_imag <= _zz_97;
      end
      if(_zz_30)begin
        img_reg_array_28_15_imag <= _zz_97;
      end
      if(_zz_31)begin
        img_reg_array_29_15_imag <= _zz_97;
      end
      if(_zz_32)begin
        img_reg_array_30_15_imag <= _zz_97;
      end
      if(_zz_33)begin
        img_reg_array_31_15_imag <= _zz_97;
      end
      if(_zz_34)begin
        img_reg_array_32_15_imag <= _zz_97;
      end
      if(_zz_35)begin
        img_reg_array_33_15_imag <= _zz_97;
      end
      if(_zz_36)begin
        img_reg_array_34_15_imag <= _zz_97;
      end
      if(_zz_37)begin
        img_reg_array_35_15_imag <= _zz_97;
      end
      if(_zz_38)begin
        img_reg_array_36_15_imag <= _zz_97;
      end
      if(_zz_39)begin
        img_reg_array_37_15_imag <= _zz_97;
      end
      if(_zz_40)begin
        img_reg_array_38_15_imag <= _zz_97;
      end
      if(_zz_41)begin
        img_reg_array_39_15_imag <= _zz_97;
      end
      if(_zz_42)begin
        img_reg_array_40_15_imag <= _zz_97;
      end
      if(_zz_43)begin
        img_reg_array_41_15_imag <= _zz_97;
      end
      if(_zz_44)begin
        img_reg_array_42_15_imag <= _zz_97;
      end
      if(_zz_45)begin
        img_reg_array_43_15_imag <= _zz_97;
      end
      if(_zz_46)begin
        img_reg_array_44_15_imag <= _zz_97;
      end
      if(_zz_47)begin
        img_reg_array_45_15_imag <= _zz_97;
      end
      if(_zz_48)begin
        img_reg_array_46_15_imag <= _zz_97;
      end
      if(_zz_49)begin
        img_reg_array_47_15_imag <= _zz_97;
      end
      if(_zz_50)begin
        img_reg_array_48_15_imag <= _zz_97;
      end
      if(_zz_51)begin
        img_reg_array_49_15_imag <= _zz_97;
      end
      if(_zz_52)begin
        img_reg_array_50_15_imag <= _zz_97;
      end
      if(_zz_53)begin
        img_reg_array_51_15_imag <= _zz_97;
      end
      if(_zz_54)begin
        img_reg_array_52_15_imag <= _zz_97;
      end
      if(_zz_55)begin
        img_reg_array_53_15_imag <= _zz_97;
      end
      if(_zz_56)begin
        img_reg_array_54_15_imag <= _zz_97;
      end
      if(_zz_57)begin
        img_reg_array_55_15_imag <= _zz_97;
      end
      if(_zz_58)begin
        img_reg_array_56_15_imag <= _zz_97;
      end
      if(_zz_59)begin
        img_reg_array_57_15_imag <= _zz_97;
      end
      if(_zz_60)begin
        img_reg_array_58_15_imag <= _zz_97;
      end
      if(_zz_61)begin
        img_reg_array_59_15_imag <= _zz_97;
      end
      if(_zz_62)begin
        img_reg_array_60_15_imag <= _zz_97;
      end
      if(_zz_63)begin
        img_reg_array_61_15_imag <= _zz_97;
      end
      if(_zz_64)begin
        img_reg_array_62_15_imag <= _zz_97;
      end
      if(_zz_65)begin
        img_reg_array_63_15_imag <= _zz_97;
      end
      if(_zz_2)begin
        img_reg_array_0_16_real <= _zz_98;
      end
      if(_zz_3)begin
        img_reg_array_1_16_real <= _zz_98;
      end
      if(_zz_4)begin
        img_reg_array_2_16_real <= _zz_98;
      end
      if(_zz_5)begin
        img_reg_array_3_16_real <= _zz_98;
      end
      if(_zz_6)begin
        img_reg_array_4_16_real <= _zz_98;
      end
      if(_zz_7)begin
        img_reg_array_5_16_real <= _zz_98;
      end
      if(_zz_8)begin
        img_reg_array_6_16_real <= _zz_98;
      end
      if(_zz_9)begin
        img_reg_array_7_16_real <= _zz_98;
      end
      if(_zz_10)begin
        img_reg_array_8_16_real <= _zz_98;
      end
      if(_zz_11)begin
        img_reg_array_9_16_real <= _zz_98;
      end
      if(_zz_12)begin
        img_reg_array_10_16_real <= _zz_98;
      end
      if(_zz_13)begin
        img_reg_array_11_16_real <= _zz_98;
      end
      if(_zz_14)begin
        img_reg_array_12_16_real <= _zz_98;
      end
      if(_zz_15)begin
        img_reg_array_13_16_real <= _zz_98;
      end
      if(_zz_16)begin
        img_reg_array_14_16_real <= _zz_98;
      end
      if(_zz_17)begin
        img_reg_array_15_16_real <= _zz_98;
      end
      if(_zz_18)begin
        img_reg_array_16_16_real <= _zz_98;
      end
      if(_zz_19)begin
        img_reg_array_17_16_real <= _zz_98;
      end
      if(_zz_20)begin
        img_reg_array_18_16_real <= _zz_98;
      end
      if(_zz_21)begin
        img_reg_array_19_16_real <= _zz_98;
      end
      if(_zz_22)begin
        img_reg_array_20_16_real <= _zz_98;
      end
      if(_zz_23)begin
        img_reg_array_21_16_real <= _zz_98;
      end
      if(_zz_24)begin
        img_reg_array_22_16_real <= _zz_98;
      end
      if(_zz_25)begin
        img_reg_array_23_16_real <= _zz_98;
      end
      if(_zz_26)begin
        img_reg_array_24_16_real <= _zz_98;
      end
      if(_zz_27)begin
        img_reg_array_25_16_real <= _zz_98;
      end
      if(_zz_28)begin
        img_reg_array_26_16_real <= _zz_98;
      end
      if(_zz_29)begin
        img_reg_array_27_16_real <= _zz_98;
      end
      if(_zz_30)begin
        img_reg_array_28_16_real <= _zz_98;
      end
      if(_zz_31)begin
        img_reg_array_29_16_real <= _zz_98;
      end
      if(_zz_32)begin
        img_reg_array_30_16_real <= _zz_98;
      end
      if(_zz_33)begin
        img_reg_array_31_16_real <= _zz_98;
      end
      if(_zz_34)begin
        img_reg_array_32_16_real <= _zz_98;
      end
      if(_zz_35)begin
        img_reg_array_33_16_real <= _zz_98;
      end
      if(_zz_36)begin
        img_reg_array_34_16_real <= _zz_98;
      end
      if(_zz_37)begin
        img_reg_array_35_16_real <= _zz_98;
      end
      if(_zz_38)begin
        img_reg_array_36_16_real <= _zz_98;
      end
      if(_zz_39)begin
        img_reg_array_37_16_real <= _zz_98;
      end
      if(_zz_40)begin
        img_reg_array_38_16_real <= _zz_98;
      end
      if(_zz_41)begin
        img_reg_array_39_16_real <= _zz_98;
      end
      if(_zz_42)begin
        img_reg_array_40_16_real <= _zz_98;
      end
      if(_zz_43)begin
        img_reg_array_41_16_real <= _zz_98;
      end
      if(_zz_44)begin
        img_reg_array_42_16_real <= _zz_98;
      end
      if(_zz_45)begin
        img_reg_array_43_16_real <= _zz_98;
      end
      if(_zz_46)begin
        img_reg_array_44_16_real <= _zz_98;
      end
      if(_zz_47)begin
        img_reg_array_45_16_real <= _zz_98;
      end
      if(_zz_48)begin
        img_reg_array_46_16_real <= _zz_98;
      end
      if(_zz_49)begin
        img_reg_array_47_16_real <= _zz_98;
      end
      if(_zz_50)begin
        img_reg_array_48_16_real <= _zz_98;
      end
      if(_zz_51)begin
        img_reg_array_49_16_real <= _zz_98;
      end
      if(_zz_52)begin
        img_reg_array_50_16_real <= _zz_98;
      end
      if(_zz_53)begin
        img_reg_array_51_16_real <= _zz_98;
      end
      if(_zz_54)begin
        img_reg_array_52_16_real <= _zz_98;
      end
      if(_zz_55)begin
        img_reg_array_53_16_real <= _zz_98;
      end
      if(_zz_56)begin
        img_reg_array_54_16_real <= _zz_98;
      end
      if(_zz_57)begin
        img_reg_array_55_16_real <= _zz_98;
      end
      if(_zz_58)begin
        img_reg_array_56_16_real <= _zz_98;
      end
      if(_zz_59)begin
        img_reg_array_57_16_real <= _zz_98;
      end
      if(_zz_60)begin
        img_reg_array_58_16_real <= _zz_98;
      end
      if(_zz_61)begin
        img_reg_array_59_16_real <= _zz_98;
      end
      if(_zz_62)begin
        img_reg_array_60_16_real <= _zz_98;
      end
      if(_zz_63)begin
        img_reg_array_61_16_real <= _zz_98;
      end
      if(_zz_64)begin
        img_reg_array_62_16_real <= _zz_98;
      end
      if(_zz_65)begin
        img_reg_array_63_16_real <= _zz_98;
      end
      if(_zz_2)begin
        img_reg_array_0_16_imag <= _zz_99;
      end
      if(_zz_3)begin
        img_reg_array_1_16_imag <= _zz_99;
      end
      if(_zz_4)begin
        img_reg_array_2_16_imag <= _zz_99;
      end
      if(_zz_5)begin
        img_reg_array_3_16_imag <= _zz_99;
      end
      if(_zz_6)begin
        img_reg_array_4_16_imag <= _zz_99;
      end
      if(_zz_7)begin
        img_reg_array_5_16_imag <= _zz_99;
      end
      if(_zz_8)begin
        img_reg_array_6_16_imag <= _zz_99;
      end
      if(_zz_9)begin
        img_reg_array_7_16_imag <= _zz_99;
      end
      if(_zz_10)begin
        img_reg_array_8_16_imag <= _zz_99;
      end
      if(_zz_11)begin
        img_reg_array_9_16_imag <= _zz_99;
      end
      if(_zz_12)begin
        img_reg_array_10_16_imag <= _zz_99;
      end
      if(_zz_13)begin
        img_reg_array_11_16_imag <= _zz_99;
      end
      if(_zz_14)begin
        img_reg_array_12_16_imag <= _zz_99;
      end
      if(_zz_15)begin
        img_reg_array_13_16_imag <= _zz_99;
      end
      if(_zz_16)begin
        img_reg_array_14_16_imag <= _zz_99;
      end
      if(_zz_17)begin
        img_reg_array_15_16_imag <= _zz_99;
      end
      if(_zz_18)begin
        img_reg_array_16_16_imag <= _zz_99;
      end
      if(_zz_19)begin
        img_reg_array_17_16_imag <= _zz_99;
      end
      if(_zz_20)begin
        img_reg_array_18_16_imag <= _zz_99;
      end
      if(_zz_21)begin
        img_reg_array_19_16_imag <= _zz_99;
      end
      if(_zz_22)begin
        img_reg_array_20_16_imag <= _zz_99;
      end
      if(_zz_23)begin
        img_reg_array_21_16_imag <= _zz_99;
      end
      if(_zz_24)begin
        img_reg_array_22_16_imag <= _zz_99;
      end
      if(_zz_25)begin
        img_reg_array_23_16_imag <= _zz_99;
      end
      if(_zz_26)begin
        img_reg_array_24_16_imag <= _zz_99;
      end
      if(_zz_27)begin
        img_reg_array_25_16_imag <= _zz_99;
      end
      if(_zz_28)begin
        img_reg_array_26_16_imag <= _zz_99;
      end
      if(_zz_29)begin
        img_reg_array_27_16_imag <= _zz_99;
      end
      if(_zz_30)begin
        img_reg_array_28_16_imag <= _zz_99;
      end
      if(_zz_31)begin
        img_reg_array_29_16_imag <= _zz_99;
      end
      if(_zz_32)begin
        img_reg_array_30_16_imag <= _zz_99;
      end
      if(_zz_33)begin
        img_reg_array_31_16_imag <= _zz_99;
      end
      if(_zz_34)begin
        img_reg_array_32_16_imag <= _zz_99;
      end
      if(_zz_35)begin
        img_reg_array_33_16_imag <= _zz_99;
      end
      if(_zz_36)begin
        img_reg_array_34_16_imag <= _zz_99;
      end
      if(_zz_37)begin
        img_reg_array_35_16_imag <= _zz_99;
      end
      if(_zz_38)begin
        img_reg_array_36_16_imag <= _zz_99;
      end
      if(_zz_39)begin
        img_reg_array_37_16_imag <= _zz_99;
      end
      if(_zz_40)begin
        img_reg_array_38_16_imag <= _zz_99;
      end
      if(_zz_41)begin
        img_reg_array_39_16_imag <= _zz_99;
      end
      if(_zz_42)begin
        img_reg_array_40_16_imag <= _zz_99;
      end
      if(_zz_43)begin
        img_reg_array_41_16_imag <= _zz_99;
      end
      if(_zz_44)begin
        img_reg_array_42_16_imag <= _zz_99;
      end
      if(_zz_45)begin
        img_reg_array_43_16_imag <= _zz_99;
      end
      if(_zz_46)begin
        img_reg_array_44_16_imag <= _zz_99;
      end
      if(_zz_47)begin
        img_reg_array_45_16_imag <= _zz_99;
      end
      if(_zz_48)begin
        img_reg_array_46_16_imag <= _zz_99;
      end
      if(_zz_49)begin
        img_reg_array_47_16_imag <= _zz_99;
      end
      if(_zz_50)begin
        img_reg_array_48_16_imag <= _zz_99;
      end
      if(_zz_51)begin
        img_reg_array_49_16_imag <= _zz_99;
      end
      if(_zz_52)begin
        img_reg_array_50_16_imag <= _zz_99;
      end
      if(_zz_53)begin
        img_reg_array_51_16_imag <= _zz_99;
      end
      if(_zz_54)begin
        img_reg_array_52_16_imag <= _zz_99;
      end
      if(_zz_55)begin
        img_reg_array_53_16_imag <= _zz_99;
      end
      if(_zz_56)begin
        img_reg_array_54_16_imag <= _zz_99;
      end
      if(_zz_57)begin
        img_reg_array_55_16_imag <= _zz_99;
      end
      if(_zz_58)begin
        img_reg_array_56_16_imag <= _zz_99;
      end
      if(_zz_59)begin
        img_reg_array_57_16_imag <= _zz_99;
      end
      if(_zz_60)begin
        img_reg_array_58_16_imag <= _zz_99;
      end
      if(_zz_61)begin
        img_reg_array_59_16_imag <= _zz_99;
      end
      if(_zz_62)begin
        img_reg_array_60_16_imag <= _zz_99;
      end
      if(_zz_63)begin
        img_reg_array_61_16_imag <= _zz_99;
      end
      if(_zz_64)begin
        img_reg_array_62_16_imag <= _zz_99;
      end
      if(_zz_65)begin
        img_reg_array_63_16_imag <= _zz_99;
      end
      if(_zz_2)begin
        img_reg_array_0_17_real <= _zz_100;
      end
      if(_zz_3)begin
        img_reg_array_1_17_real <= _zz_100;
      end
      if(_zz_4)begin
        img_reg_array_2_17_real <= _zz_100;
      end
      if(_zz_5)begin
        img_reg_array_3_17_real <= _zz_100;
      end
      if(_zz_6)begin
        img_reg_array_4_17_real <= _zz_100;
      end
      if(_zz_7)begin
        img_reg_array_5_17_real <= _zz_100;
      end
      if(_zz_8)begin
        img_reg_array_6_17_real <= _zz_100;
      end
      if(_zz_9)begin
        img_reg_array_7_17_real <= _zz_100;
      end
      if(_zz_10)begin
        img_reg_array_8_17_real <= _zz_100;
      end
      if(_zz_11)begin
        img_reg_array_9_17_real <= _zz_100;
      end
      if(_zz_12)begin
        img_reg_array_10_17_real <= _zz_100;
      end
      if(_zz_13)begin
        img_reg_array_11_17_real <= _zz_100;
      end
      if(_zz_14)begin
        img_reg_array_12_17_real <= _zz_100;
      end
      if(_zz_15)begin
        img_reg_array_13_17_real <= _zz_100;
      end
      if(_zz_16)begin
        img_reg_array_14_17_real <= _zz_100;
      end
      if(_zz_17)begin
        img_reg_array_15_17_real <= _zz_100;
      end
      if(_zz_18)begin
        img_reg_array_16_17_real <= _zz_100;
      end
      if(_zz_19)begin
        img_reg_array_17_17_real <= _zz_100;
      end
      if(_zz_20)begin
        img_reg_array_18_17_real <= _zz_100;
      end
      if(_zz_21)begin
        img_reg_array_19_17_real <= _zz_100;
      end
      if(_zz_22)begin
        img_reg_array_20_17_real <= _zz_100;
      end
      if(_zz_23)begin
        img_reg_array_21_17_real <= _zz_100;
      end
      if(_zz_24)begin
        img_reg_array_22_17_real <= _zz_100;
      end
      if(_zz_25)begin
        img_reg_array_23_17_real <= _zz_100;
      end
      if(_zz_26)begin
        img_reg_array_24_17_real <= _zz_100;
      end
      if(_zz_27)begin
        img_reg_array_25_17_real <= _zz_100;
      end
      if(_zz_28)begin
        img_reg_array_26_17_real <= _zz_100;
      end
      if(_zz_29)begin
        img_reg_array_27_17_real <= _zz_100;
      end
      if(_zz_30)begin
        img_reg_array_28_17_real <= _zz_100;
      end
      if(_zz_31)begin
        img_reg_array_29_17_real <= _zz_100;
      end
      if(_zz_32)begin
        img_reg_array_30_17_real <= _zz_100;
      end
      if(_zz_33)begin
        img_reg_array_31_17_real <= _zz_100;
      end
      if(_zz_34)begin
        img_reg_array_32_17_real <= _zz_100;
      end
      if(_zz_35)begin
        img_reg_array_33_17_real <= _zz_100;
      end
      if(_zz_36)begin
        img_reg_array_34_17_real <= _zz_100;
      end
      if(_zz_37)begin
        img_reg_array_35_17_real <= _zz_100;
      end
      if(_zz_38)begin
        img_reg_array_36_17_real <= _zz_100;
      end
      if(_zz_39)begin
        img_reg_array_37_17_real <= _zz_100;
      end
      if(_zz_40)begin
        img_reg_array_38_17_real <= _zz_100;
      end
      if(_zz_41)begin
        img_reg_array_39_17_real <= _zz_100;
      end
      if(_zz_42)begin
        img_reg_array_40_17_real <= _zz_100;
      end
      if(_zz_43)begin
        img_reg_array_41_17_real <= _zz_100;
      end
      if(_zz_44)begin
        img_reg_array_42_17_real <= _zz_100;
      end
      if(_zz_45)begin
        img_reg_array_43_17_real <= _zz_100;
      end
      if(_zz_46)begin
        img_reg_array_44_17_real <= _zz_100;
      end
      if(_zz_47)begin
        img_reg_array_45_17_real <= _zz_100;
      end
      if(_zz_48)begin
        img_reg_array_46_17_real <= _zz_100;
      end
      if(_zz_49)begin
        img_reg_array_47_17_real <= _zz_100;
      end
      if(_zz_50)begin
        img_reg_array_48_17_real <= _zz_100;
      end
      if(_zz_51)begin
        img_reg_array_49_17_real <= _zz_100;
      end
      if(_zz_52)begin
        img_reg_array_50_17_real <= _zz_100;
      end
      if(_zz_53)begin
        img_reg_array_51_17_real <= _zz_100;
      end
      if(_zz_54)begin
        img_reg_array_52_17_real <= _zz_100;
      end
      if(_zz_55)begin
        img_reg_array_53_17_real <= _zz_100;
      end
      if(_zz_56)begin
        img_reg_array_54_17_real <= _zz_100;
      end
      if(_zz_57)begin
        img_reg_array_55_17_real <= _zz_100;
      end
      if(_zz_58)begin
        img_reg_array_56_17_real <= _zz_100;
      end
      if(_zz_59)begin
        img_reg_array_57_17_real <= _zz_100;
      end
      if(_zz_60)begin
        img_reg_array_58_17_real <= _zz_100;
      end
      if(_zz_61)begin
        img_reg_array_59_17_real <= _zz_100;
      end
      if(_zz_62)begin
        img_reg_array_60_17_real <= _zz_100;
      end
      if(_zz_63)begin
        img_reg_array_61_17_real <= _zz_100;
      end
      if(_zz_64)begin
        img_reg_array_62_17_real <= _zz_100;
      end
      if(_zz_65)begin
        img_reg_array_63_17_real <= _zz_100;
      end
      if(_zz_2)begin
        img_reg_array_0_17_imag <= _zz_101;
      end
      if(_zz_3)begin
        img_reg_array_1_17_imag <= _zz_101;
      end
      if(_zz_4)begin
        img_reg_array_2_17_imag <= _zz_101;
      end
      if(_zz_5)begin
        img_reg_array_3_17_imag <= _zz_101;
      end
      if(_zz_6)begin
        img_reg_array_4_17_imag <= _zz_101;
      end
      if(_zz_7)begin
        img_reg_array_5_17_imag <= _zz_101;
      end
      if(_zz_8)begin
        img_reg_array_6_17_imag <= _zz_101;
      end
      if(_zz_9)begin
        img_reg_array_7_17_imag <= _zz_101;
      end
      if(_zz_10)begin
        img_reg_array_8_17_imag <= _zz_101;
      end
      if(_zz_11)begin
        img_reg_array_9_17_imag <= _zz_101;
      end
      if(_zz_12)begin
        img_reg_array_10_17_imag <= _zz_101;
      end
      if(_zz_13)begin
        img_reg_array_11_17_imag <= _zz_101;
      end
      if(_zz_14)begin
        img_reg_array_12_17_imag <= _zz_101;
      end
      if(_zz_15)begin
        img_reg_array_13_17_imag <= _zz_101;
      end
      if(_zz_16)begin
        img_reg_array_14_17_imag <= _zz_101;
      end
      if(_zz_17)begin
        img_reg_array_15_17_imag <= _zz_101;
      end
      if(_zz_18)begin
        img_reg_array_16_17_imag <= _zz_101;
      end
      if(_zz_19)begin
        img_reg_array_17_17_imag <= _zz_101;
      end
      if(_zz_20)begin
        img_reg_array_18_17_imag <= _zz_101;
      end
      if(_zz_21)begin
        img_reg_array_19_17_imag <= _zz_101;
      end
      if(_zz_22)begin
        img_reg_array_20_17_imag <= _zz_101;
      end
      if(_zz_23)begin
        img_reg_array_21_17_imag <= _zz_101;
      end
      if(_zz_24)begin
        img_reg_array_22_17_imag <= _zz_101;
      end
      if(_zz_25)begin
        img_reg_array_23_17_imag <= _zz_101;
      end
      if(_zz_26)begin
        img_reg_array_24_17_imag <= _zz_101;
      end
      if(_zz_27)begin
        img_reg_array_25_17_imag <= _zz_101;
      end
      if(_zz_28)begin
        img_reg_array_26_17_imag <= _zz_101;
      end
      if(_zz_29)begin
        img_reg_array_27_17_imag <= _zz_101;
      end
      if(_zz_30)begin
        img_reg_array_28_17_imag <= _zz_101;
      end
      if(_zz_31)begin
        img_reg_array_29_17_imag <= _zz_101;
      end
      if(_zz_32)begin
        img_reg_array_30_17_imag <= _zz_101;
      end
      if(_zz_33)begin
        img_reg_array_31_17_imag <= _zz_101;
      end
      if(_zz_34)begin
        img_reg_array_32_17_imag <= _zz_101;
      end
      if(_zz_35)begin
        img_reg_array_33_17_imag <= _zz_101;
      end
      if(_zz_36)begin
        img_reg_array_34_17_imag <= _zz_101;
      end
      if(_zz_37)begin
        img_reg_array_35_17_imag <= _zz_101;
      end
      if(_zz_38)begin
        img_reg_array_36_17_imag <= _zz_101;
      end
      if(_zz_39)begin
        img_reg_array_37_17_imag <= _zz_101;
      end
      if(_zz_40)begin
        img_reg_array_38_17_imag <= _zz_101;
      end
      if(_zz_41)begin
        img_reg_array_39_17_imag <= _zz_101;
      end
      if(_zz_42)begin
        img_reg_array_40_17_imag <= _zz_101;
      end
      if(_zz_43)begin
        img_reg_array_41_17_imag <= _zz_101;
      end
      if(_zz_44)begin
        img_reg_array_42_17_imag <= _zz_101;
      end
      if(_zz_45)begin
        img_reg_array_43_17_imag <= _zz_101;
      end
      if(_zz_46)begin
        img_reg_array_44_17_imag <= _zz_101;
      end
      if(_zz_47)begin
        img_reg_array_45_17_imag <= _zz_101;
      end
      if(_zz_48)begin
        img_reg_array_46_17_imag <= _zz_101;
      end
      if(_zz_49)begin
        img_reg_array_47_17_imag <= _zz_101;
      end
      if(_zz_50)begin
        img_reg_array_48_17_imag <= _zz_101;
      end
      if(_zz_51)begin
        img_reg_array_49_17_imag <= _zz_101;
      end
      if(_zz_52)begin
        img_reg_array_50_17_imag <= _zz_101;
      end
      if(_zz_53)begin
        img_reg_array_51_17_imag <= _zz_101;
      end
      if(_zz_54)begin
        img_reg_array_52_17_imag <= _zz_101;
      end
      if(_zz_55)begin
        img_reg_array_53_17_imag <= _zz_101;
      end
      if(_zz_56)begin
        img_reg_array_54_17_imag <= _zz_101;
      end
      if(_zz_57)begin
        img_reg_array_55_17_imag <= _zz_101;
      end
      if(_zz_58)begin
        img_reg_array_56_17_imag <= _zz_101;
      end
      if(_zz_59)begin
        img_reg_array_57_17_imag <= _zz_101;
      end
      if(_zz_60)begin
        img_reg_array_58_17_imag <= _zz_101;
      end
      if(_zz_61)begin
        img_reg_array_59_17_imag <= _zz_101;
      end
      if(_zz_62)begin
        img_reg_array_60_17_imag <= _zz_101;
      end
      if(_zz_63)begin
        img_reg_array_61_17_imag <= _zz_101;
      end
      if(_zz_64)begin
        img_reg_array_62_17_imag <= _zz_101;
      end
      if(_zz_65)begin
        img_reg_array_63_17_imag <= _zz_101;
      end
      if(_zz_2)begin
        img_reg_array_0_18_real <= _zz_102;
      end
      if(_zz_3)begin
        img_reg_array_1_18_real <= _zz_102;
      end
      if(_zz_4)begin
        img_reg_array_2_18_real <= _zz_102;
      end
      if(_zz_5)begin
        img_reg_array_3_18_real <= _zz_102;
      end
      if(_zz_6)begin
        img_reg_array_4_18_real <= _zz_102;
      end
      if(_zz_7)begin
        img_reg_array_5_18_real <= _zz_102;
      end
      if(_zz_8)begin
        img_reg_array_6_18_real <= _zz_102;
      end
      if(_zz_9)begin
        img_reg_array_7_18_real <= _zz_102;
      end
      if(_zz_10)begin
        img_reg_array_8_18_real <= _zz_102;
      end
      if(_zz_11)begin
        img_reg_array_9_18_real <= _zz_102;
      end
      if(_zz_12)begin
        img_reg_array_10_18_real <= _zz_102;
      end
      if(_zz_13)begin
        img_reg_array_11_18_real <= _zz_102;
      end
      if(_zz_14)begin
        img_reg_array_12_18_real <= _zz_102;
      end
      if(_zz_15)begin
        img_reg_array_13_18_real <= _zz_102;
      end
      if(_zz_16)begin
        img_reg_array_14_18_real <= _zz_102;
      end
      if(_zz_17)begin
        img_reg_array_15_18_real <= _zz_102;
      end
      if(_zz_18)begin
        img_reg_array_16_18_real <= _zz_102;
      end
      if(_zz_19)begin
        img_reg_array_17_18_real <= _zz_102;
      end
      if(_zz_20)begin
        img_reg_array_18_18_real <= _zz_102;
      end
      if(_zz_21)begin
        img_reg_array_19_18_real <= _zz_102;
      end
      if(_zz_22)begin
        img_reg_array_20_18_real <= _zz_102;
      end
      if(_zz_23)begin
        img_reg_array_21_18_real <= _zz_102;
      end
      if(_zz_24)begin
        img_reg_array_22_18_real <= _zz_102;
      end
      if(_zz_25)begin
        img_reg_array_23_18_real <= _zz_102;
      end
      if(_zz_26)begin
        img_reg_array_24_18_real <= _zz_102;
      end
      if(_zz_27)begin
        img_reg_array_25_18_real <= _zz_102;
      end
      if(_zz_28)begin
        img_reg_array_26_18_real <= _zz_102;
      end
      if(_zz_29)begin
        img_reg_array_27_18_real <= _zz_102;
      end
      if(_zz_30)begin
        img_reg_array_28_18_real <= _zz_102;
      end
      if(_zz_31)begin
        img_reg_array_29_18_real <= _zz_102;
      end
      if(_zz_32)begin
        img_reg_array_30_18_real <= _zz_102;
      end
      if(_zz_33)begin
        img_reg_array_31_18_real <= _zz_102;
      end
      if(_zz_34)begin
        img_reg_array_32_18_real <= _zz_102;
      end
      if(_zz_35)begin
        img_reg_array_33_18_real <= _zz_102;
      end
      if(_zz_36)begin
        img_reg_array_34_18_real <= _zz_102;
      end
      if(_zz_37)begin
        img_reg_array_35_18_real <= _zz_102;
      end
      if(_zz_38)begin
        img_reg_array_36_18_real <= _zz_102;
      end
      if(_zz_39)begin
        img_reg_array_37_18_real <= _zz_102;
      end
      if(_zz_40)begin
        img_reg_array_38_18_real <= _zz_102;
      end
      if(_zz_41)begin
        img_reg_array_39_18_real <= _zz_102;
      end
      if(_zz_42)begin
        img_reg_array_40_18_real <= _zz_102;
      end
      if(_zz_43)begin
        img_reg_array_41_18_real <= _zz_102;
      end
      if(_zz_44)begin
        img_reg_array_42_18_real <= _zz_102;
      end
      if(_zz_45)begin
        img_reg_array_43_18_real <= _zz_102;
      end
      if(_zz_46)begin
        img_reg_array_44_18_real <= _zz_102;
      end
      if(_zz_47)begin
        img_reg_array_45_18_real <= _zz_102;
      end
      if(_zz_48)begin
        img_reg_array_46_18_real <= _zz_102;
      end
      if(_zz_49)begin
        img_reg_array_47_18_real <= _zz_102;
      end
      if(_zz_50)begin
        img_reg_array_48_18_real <= _zz_102;
      end
      if(_zz_51)begin
        img_reg_array_49_18_real <= _zz_102;
      end
      if(_zz_52)begin
        img_reg_array_50_18_real <= _zz_102;
      end
      if(_zz_53)begin
        img_reg_array_51_18_real <= _zz_102;
      end
      if(_zz_54)begin
        img_reg_array_52_18_real <= _zz_102;
      end
      if(_zz_55)begin
        img_reg_array_53_18_real <= _zz_102;
      end
      if(_zz_56)begin
        img_reg_array_54_18_real <= _zz_102;
      end
      if(_zz_57)begin
        img_reg_array_55_18_real <= _zz_102;
      end
      if(_zz_58)begin
        img_reg_array_56_18_real <= _zz_102;
      end
      if(_zz_59)begin
        img_reg_array_57_18_real <= _zz_102;
      end
      if(_zz_60)begin
        img_reg_array_58_18_real <= _zz_102;
      end
      if(_zz_61)begin
        img_reg_array_59_18_real <= _zz_102;
      end
      if(_zz_62)begin
        img_reg_array_60_18_real <= _zz_102;
      end
      if(_zz_63)begin
        img_reg_array_61_18_real <= _zz_102;
      end
      if(_zz_64)begin
        img_reg_array_62_18_real <= _zz_102;
      end
      if(_zz_65)begin
        img_reg_array_63_18_real <= _zz_102;
      end
      if(_zz_2)begin
        img_reg_array_0_18_imag <= _zz_103;
      end
      if(_zz_3)begin
        img_reg_array_1_18_imag <= _zz_103;
      end
      if(_zz_4)begin
        img_reg_array_2_18_imag <= _zz_103;
      end
      if(_zz_5)begin
        img_reg_array_3_18_imag <= _zz_103;
      end
      if(_zz_6)begin
        img_reg_array_4_18_imag <= _zz_103;
      end
      if(_zz_7)begin
        img_reg_array_5_18_imag <= _zz_103;
      end
      if(_zz_8)begin
        img_reg_array_6_18_imag <= _zz_103;
      end
      if(_zz_9)begin
        img_reg_array_7_18_imag <= _zz_103;
      end
      if(_zz_10)begin
        img_reg_array_8_18_imag <= _zz_103;
      end
      if(_zz_11)begin
        img_reg_array_9_18_imag <= _zz_103;
      end
      if(_zz_12)begin
        img_reg_array_10_18_imag <= _zz_103;
      end
      if(_zz_13)begin
        img_reg_array_11_18_imag <= _zz_103;
      end
      if(_zz_14)begin
        img_reg_array_12_18_imag <= _zz_103;
      end
      if(_zz_15)begin
        img_reg_array_13_18_imag <= _zz_103;
      end
      if(_zz_16)begin
        img_reg_array_14_18_imag <= _zz_103;
      end
      if(_zz_17)begin
        img_reg_array_15_18_imag <= _zz_103;
      end
      if(_zz_18)begin
        img_reg_array_16_18_imag <= _zz_103;
      end
      if(_zz_19)begin
        img_reg_array_17_18_imag <= _zz_103;
      end
      if(_zz_20)begin
        img_reg_array_18_18_imag <= _zz_103;
      end
      if(_zz_21)begin
        img_reg_array_19_18_imag <= _zz_103;
      end
      if(_zz_22)begin
        img_reg_array_20_18_imag <= _zz_103;
      end
      if(_zz_23)begin
        img_reg_array_21_18_imag <= _zz_103;
      end
      if(_zz_24)begin
        img_reg_array_22_18_imag <= _zz_103;
      end
      if(_zz_25)begin
        img_reg_array_23_18_imag <= _zz_103;
      end
      if(_zz_26)begin
        img_reg_array_24_18_imag <= _zz_103;
      end
      if(_zz_27)begin
        img_reg_array_25_18_imag <= _zz_103;
      end
      if(_zz_28)begin
        img_reg_array_26_18_imag <= _zz_103;
      end
      if(_zz_29)begin
        img_reg_array_27_18_imag <= _zz_103;
      end
      if(_zz_30)begin
        img_reg_array_28_18_imag <= _zz_103;
      end
      if(_zz_31)begin
        img_reg_array_29_18_imag <= _zz_103;
      end
      if(_zz_32)begin
        img_reg_array_30_18_imag <= _zz_103;
      end
      if(_zz_33)begin
        img_reg_array_31_18_imag <= _zz_103;
      end
      if(_zz_34)begin
        img_reg_array_32_18_imag <= _zz_103;
      end
      if(_zz_35)begin
        img_reg_array_33_18_imag <= _zz_103;
      end
      if(_zz_36)begin
        img_reg_array_34_18_imag <= _zz_103;
      end
      if(_zz_37)begin
        img_reg_array_35_18_imag <= _zz_103;
      end
      if(_zz_38)begin
        img_reg_array_36_18_imag <= _zz_103;
      end
      if(_zz_39)begin
        img_reg_array_37_18_imag <= _zz_103;
      end
      if(_zz_40)begin
        img_reg_array_38_18_imag <= _zz_103;
      end
      if(_zz_41)begin
        img_reg_array_39_18_imag <= _zz_103;
      end
      if(_zz_42)begin
        img_reg_array_40_18_imag <= _zz_103;
      end
      if(_zz_43)begin
        img_reg_array_41_18_imag <= _zz_103;
      end
      if(_zz_44)begin
        img_reg_array_42_18_imag <= _zz_103;
      end
      if(_zz_45)begin
        img_reg_array_43_18_imag <= _zz_103;
      end
      if(_zz_46)begin
        img_reg_array_44_18_imag <= _zz_103;
      end
      if(_zz_47)begin
        img_reg_array_45_18_imag <= _zz_103;
      end
      if(_zz_48)begin
        img_reg_array_46_18_imag <= _zz_103;
      end
      if(_zz_49)begin
        img_reg_array_47_18_imag <= _zz_103;
      end
      if(_zz_50)begin
        img_reg_array_48_18_imag <= _zz_103;
      end
      if(_zz_51)begin
        img_reg_array_49_18_imag <= _zz_103;
      end
      if(_zz_52)begin
        img_reg_array_50_18_imag <= _zz_103;
      end
      if(_zz_53)begin
        img_reg_array_51_18_imag <= _zz_103;
      end
      if(_zz_54)begin
        img_reg_array_52_18_imag <= _zz_103;
      end
      if(_zz_55)begin
        img_reg_array_53_18_imag <= _zz_103;
      end
      if(_zz_56)begin
        img_reg_array_54_18_imag <= _zz_103;
      end
      if(_zz_57)begin
        img_reg_array_55_18_imag <= _zz_103;
      end
      if(_zz_58)begin
        img_reg_array_56_18_imag <= _zz_103;
      end
      if(_zz_59)begin
        img_reg_array_57_18_imag <= _zz_103;
      end
      if(_zz_60)begin
        img_reg_array_58_18_imag <= _zz_103;
      end
      if(_zz_61)begin
        img_reg_array_59_18_imag <= _zz_103;
      end
      if(_zz_62)begin
        img_reg_array_60_18_imag <= _zz_103;
      end
      if(_zz_63)begin
        img_reg_array_61_18_imag <= _zz_103;
      end
      if(_zz_64)begin
        img_reg_array_62_18_imag <= _zz_103;
      end
      if(_zz_65)begin
        img_reg_array_63_18_imag <= _zz_103;
      end
      if(_zz_2)begin
        img_reg_array_0_19_real <= _zz_104;
      end
      if(_zz_3)begin
        img_reg_array_1_19_real <= _zz_104;
      end
      if(_zz_4)begin
        img_reg_array_2_19_real <= _zz_104;
      end
      if(_zz_5)begin
        img_reg_array_3_19_real <= _zz_104;
      end
      if(_zz_6)begin
        img_reg_array_4_19_real <= _zz_104;
      end
      if(_zz_7)begin
        img_reg_array_5_19_real <= _zz_104;
      end
      if(_zz_8)begin
        img_reg_array_6_19_real <= _zz_104;
      end
      if(_zz_9)begin
        img_reg_array_7_19_real <= _zz_104;
      end
      if(_zz_10)begin
        img_reg_array_8_19_real <= _zz_104;
      end
      if(_zz_11)begin
        img_reg_array_9_19_real <= _zz_104;
      end
      if(_zz_12)begin
        img_reg_array_10_19_real <= _zz_104;
      end
      if(_zz_13)begin
        img_reg_array_11_19_real <= _zz_104;
      end
      if(_zz_14)begin
        img_reg_array_12_19_real <= _zz_104;
      end
      if(_zz_15)begin
        img_reg_array_13_19_real <= _zz_104;
      end
      if(_zz_16)begin
        img_reg_array_14_19_real <= _zz_104;
      end
      if(_zz_17)begin
        img_reg_array_15_19_real <= _zz_104;
      end
      if(_zz_18)begin
        img_reg_array_16_19_real <= _zz_104;
      end
      if(_zz_19)begin
        img_reg_array_17_19_real <= _zz_104;
      end
      if(_zz_20)begin
        img_reg_array_18_19_real <= _zz_104;
      end
      if(_zz_21)begin
        img_reg_array_19_19_real <= _zz_104;
      end
      if(_zz_22)begin
        img_reg_array_20_19_real <= _zz_104;
      end
      if(_zz_23)begin
        img_reg_array_21_19_real <= _zz_104;
      end
      if(_zz_24)begin
        img_reg_array_22_19_real <= _zz_104;
      end
      if(_zz_25)begin
        img_reg_array_23_19_real <= _zz_104;
      end
      if(_zz_26)begin
        img_reg_array_24_19_real <= _zz_104;
      end
      if(_zz_27)begin
        img_reg_array_25_19_real <= _zz_104;
      end
      if(_zz_28)begin
        img_reg_array_26_19_real <= _zz_104;
      end
      if(_zz_29)begin
        img_reg_array_27_19_real <= _zz_104;
      end
      if(_zz_30)begin
        img_reg_array_28_19_real <= _zz_104;
      end
      if(_zz_31)begin
        img_reg_array_29_19_real <= _zz_104;
      end
      if(_zz_32)begin
        img_reg_array_30_19_real <= _zz_104;
      end
      if(_zz_33)begin
        img_reg_array_31_19_real <= _zz_104;
      end
      if(_zz_34)begin
        img_reg_array_32_19_real <= _zz_104;
      end
      if(_zz_35)begin
        img_reg_array_33_19_real <= _zz_104;
      end
      if(_zz_36)begin
        img_reg_array_34_19_real <= _zz_104;
      end
      if(_zz_37)begin
        img_reg_array_35_19_real <= _zz_104;
      end
      if(_zz_38)begin
        img_reg_array_36_19_real <= _zz_104;
      end
      if(_zz_39)begin
        img_reg_array_37_19_real <= _zz_104;
      end
      if(_zz_40)begin
        img_reg_array_38_19_real <= _zz_104;
      end
      if(_zz_41)begin
        img_reg_array_39_19_real <= _zz_104;
      end
      if(_zz_42)begin
        img_reg_array_40_19_real <= _zz_104;
      end
      if(_zz_43)begin
        img_reg_array_41_19_real <= _zz_104;
      end
      if(_zz_44)begin
        img_reg_array_42_19_real <= _zz_104;
      end
      if(_zz_45)begin
        img_reg_array_43_19_real <= _zz_104;
      end
      if(_zz_46)begin
        img_reg_array_44_19_real <= _zz_104;
      end
      if(_zz_47)begin
        img_reg_array_45_19_real <= _zz_104;
      end
      if(_zz_48)begin
        img_reg_array_46_19_real <= _zz_104;
      end
      if(_zz_49)begin
        img_reg_array_47_19_real <= _zz_104;
      end
      if(_zz_50)begin
        img_reg_array_48_19_real <= _zz_104;
      end
      if(_zz_51)begin
        img_reg_array_49_19_real <= _zz_104;
      end
      if(_zz_52)begin
        img_reg_array_50_19_real <= _zz_104;
      end
      if(_zz_53)begin
        img_reg_array_51_19_real <= _zz_104;
      end
      if(_zz_54)begin
        img_reg_array_52_19_real <= _zz_104;
      end
      if(_zz_55)begin
        img_reg_array_53_19_real <= _zz_104;
      end
      if(_zz_56)begin
        img_reg_array_54_19_real <= _zz_104;
      end
      if(_zz_57)begin
        img_reg_array_55_19_real <= _zz_104;
      end
      if(_zz_58)begin
        img_reg_array_56_19_real <= _zz_104;
      end
      if(_zz_59)begin
        img_reg_array_57_19_real <= _zz_104;
      end
      if(_zz_60)begin
        img_reg_array_58_19_real <= _zz_104;
      end
      if(_zz_61)begin
        img_reg_array_59_19_real <= _zz_104;
      end
      if(_zz_62)begin
        img_reg_array_60_19_real <= _zz_104;
      end
      if(_zz_63)begin
        img_reg_array_61_19_real <= _zz_104;
      end
      if(_zz_64)begin
        img_reg_array_62_19_real <= _zz_104;
      end
      if(_zz_65)begin
        img_reg_array_63_19_real <= _zz_104;
      end
      if(_zz_2)begin
        img_reg_array_0_19_imag <= _zz_105;
      end
      if(_zz_3)begin
        img_reg_array_1_19_imag <= _zz_105;
      end
      if(_zz_4)begin
        img_reg_array_2_19_imag <= _zz_105;
      end
      if(_zz_5)begin
        img_reg_array_3_19_imag <= _zz_105;
      end
      if(_zz_6)begin
        img_reg_array_4_19_imag <= _zz_105;
      end
      if(_zz_7)begin
        img_reg_array_5_19_imag <= _zz_105;
      end
      if(_zz_8)begin
        img_reg_array_6_19_imag <= _zz_105;
      end
      if(_zz_9)begin
        img_reg_array_7_19_imag <= _zz_105;
      end
      if(_zz_10)begin
        img_reg_array_8_19_imag <= _zz_105;
      end
      if(_zz_11)begin
        img_reg_array_9_19_imag <= _zz_105;
      end
      if(_zz_12)begin
        img_reg_array_10_19_imag <= _zz_105;
      end
      if(_zz_13)begin
        img_reg_array_11_19_imag <= _zz_105;
      end
      if(_zz_14)begin
        img_reg_array_12_19_imag <= _zz_105;
      end
      if(_zz_15)begin
        img_reg_array_13_19_imag <= _zz_105;
      end
      if(_zz_16)begin
        img_reg_array_14_19_imag <= _zz_105;
      end
      if(_zz_17)begin
        img_reg_array_15_19_imag <= _zz_105;
      end
      if(_zz_18)begin
        img_reg_array_16_19_imag <= _zz_105;
      end
      if(_zz_19)begin
        img_reg_array_17_19_imag <= _zz_105;
      end
      if(_zz_20)begin
        img_reg_array_18_19_imag <= _zz_105;
      end
      if(_zz_21)begin
        img_reg_array_19_19_imag <= _zz_105;
      end
      if(_zz_22)begin
        img_reg_array_20_19_imag <= _zz_105;
      end
      if(_zz_23)begin
        img_reg_array_21_19_imag <= _zz_105;
      end
      if(_zz_24)begin
        img_reg_array_22_19_imag <= _zz_105;
      end
      if(_zz_25)begin
        img_reg_array_23_19_imag <= _zz_105;
      end
      if(_zz_26)begin
        img_reg_array_24_19_imag <= _zz_105;
      end
      if(_zz_27)begin
        img_reg_array_25_19_imag <= _zz_105;
      end
      if(_zz_28)begin
        img_reg_array_26_19_imag <= _zz_105;
      end
      if(_zz_29)begin
        img_reg_array_27_19_imag <= _zz_105;
      end
      if(_zz_30)begin
        img_reg_array_28_19_imag <= _zz_105;
      end
      if(_zz_31)begin
        img_reg_array_29_19_imag <= _zz_105;
      end
      if(_zz_32)begin
        img_reg_array_30_19_imag <= _zz_105;
      end
      if(_zz_33)begin
        img_reg_array_31_19_imag <= _zz_105;
      end
      if(_zz_34)begin
        img_reg_array_32_19_imag <= _zz_105;
      end
      if(_zz_35)begin
        img_reg_array_33_19_imag <= _zz_105;
      end
      if(_zz_36)begin
        img_reg_array_34_19_imag <= _zz_105;
      end
      if(_zz_37)begin
        img_reg_array_35_19_imag <= _zz_105;
      end
      if(_zz_38)begin
        img_reg_array_36_19_imag <= _zz_105;
      end
      if(_zz_39)begin
        img_reg_array_37_19_imag <= _zz_105;
      end
      if(_zz_40)begin
        img_reg_array_38_19_imag <= _zz_105;
      end
      if(_zz_41)begin
        img_reg_array_39_19_imag <= _zz_105;
      end
      if(_zz_42)begin
        img_reg_array_40_19_imag <= _zz_105;
      end
      if(_zz_43)begin
        img_reg_array_41_19_imag <= _zz_105;
      end
      if(_zz_44)begin
        img_reg_array_42_19_imag <= _zz_105;
      end
      if(_zz_45)begin
        img_reg_array_43_19_imag <= _zz_105;
      end
      if(_zz_46)begin
        img_reg_array_44_19_imag <= _zz_105;
      end
      if(_zz_47)begin
        img_reg_array_45_19_imag <= _zz_105;
      end
      if(_zz_48)begin
        img_reg_array_46_19_imag <= _zz_105;
      end
      if(_zz_49)begin
        img_reg_array_47_19_imag <= _zz_105;
      end
      if(_zz_50)begin
        img_reg_array_48_19_imag <= _zz_105;
      end
      if(_zz_51)begin
        img_reg_array_49_19_imag <= _zz_105;
      end
      if(_zz_52)begin
        img_reg_array_50_19_imag <= _zz_105;
      end
      if(_zz_53)begin
        img_reg_array_51_19_imag <= _zz_105;
      end
      if(_zz_54)begin
        img_reg_array_52_19_imag <= _zz_105;
      end
      if(_zz_55)begin
        img_reg_array_53_19_imag <= _zz_105;
      end
      if(_zz_56)begin
        img_reg_array_54_19_imag <= _zz_105;
      end
      if(_zz_57)begin
        img_reg_array_55_19_imag <= _zz_105;
      end
      if(_zz_58)begin
        img_reg_array_56_19_imag <= _zz_105;
      end
      if(_zz_59)begin
        img_reg_array_57_19_imag <= _zz_105;
      end
      if(_zz_60)begin
        img_reg_array_58_19_imag <= _zz_105;
      end
      if(_zz_61)begin
        img_reg_array_59_19_imag <= _zz_105;
      end
      if(_zz_62)begin
        img_reg_array_60_19_imag <= _zz_105;
      end
      if(_zz_63)begin
        img_reg_array_61_19_imag <= _zz_105;
      end
      if(_zz_64)begin
        img_reg_array_62_19_imag <= _zz_105;
      end
      if(_zz_65)begin
        img_reg_array_63_19_imag <= _zz_105;
      end
      if(_zz_2)begin
        img_reg_array_0_20_real <= _zz_106;
      end
      if(_zz_3)begin
        img_reg_array_1_20_real <= _zz_106;
      end
      if(_zz_4)begin
        img_reg_array_2_20_real <= _zz_106;
      end
      if(_zz_5)begin
        img_reg_array_3_20_real <= _zz_106;
      end
      if(_zz_6)begin
        img_reg_array_4_20_real <= _zz_106;
      end
      if(_zz_7)begin
        img_reg_array_5_20_real <= _zz_106;
      end
      if(_zz_8)begin
        img_reg_array_6_20_real <= _zz_106;
      end
      if(_zz_9)begin
        img_reg_array_7_20_real <= _zz_106;
      end
      if(_zz_10)begin
        img_reg_array_8_20_real <= _zz_106;
      end
      if(_zz_11)begin
        img_reg_array_9_20_real <= _zz_106;
      end
      if(_zz_12)begin
        img_reg_array_10_20_real <= _zz_106;
      end
      if(_zz_13)begin
        img_reg_array_11_20_real <= _zz_106;
      end
      if(_zz_14)begin
        img_reg_array_12_20_real <= _zz_106;
      end
      if(_zz_15)begin
        img_reg_array_13_20_real <= _zz_106;
      end
      if(_zz_16)begin
        img_reg_array_14_20_real <= _zz_106;
      end
      if(_zz_17)begin
        img_reg_array_15_20_real <= _zz_106;
      end
      if(_zz_18)begin
        img_reg_array_16_20_real <= _zz_106;
      end
      if(_zz_19)begin
        img_reg_array_17_20_real <= _zz_106;
      end
      if(_zz_20)begin
        img_reg_array_18_20_real <= _zz_106;
      end
      if(_zz_21)begin
        img_reg_array_19_20_real <= _zz_106;
      end
      if(_zz_22)begin
        img_reg_array_20_20_real <= _zz_106;
      end
      if(_zz_23)begin
        img_reg_array_21_20_real <= _zz_106;
      end
      if(_zz_24)begin
        img_reg_array_22_20_real <= _zz_106;
      end
      if(_zz_25)begin
        img_reg_array_23_20_real <= _zz_106;
      end
      if(_zz_26)begin
        img_reg_array_24_20_real <= _zz_106;
      end
      if(_zz_27)begin
        img_reg_array_25_20_real <= _zz_106;
      end
      if(_zz_28)begin
        img_reg_array_26_20_real <= _zz_106;
      end
      if(_zz_29)begin
        img_reg_array_27_20_real <= _zz_106;
      end
      if(_zz_30)begin
        img_reg_array_28_20_real <= _zz_106;
      end
      if(_zz_31)begin
        img_reg_array_29_20_real <= _zz_106;
      end
      if(_zz_32)begin
        img_reg_array_30_20_real <= _zz_106;
      end
      if(_zz_33)begin
        img_reg_array_31_20_real <= _zz_106;
      end
      if(_zz_34)begin
        img_reg_array_32_20_real <= _zz_106;
      end
      if(_zz_35)begin
        img_reg_array_33_20_real <= _zz_106;
      end
      if(_zz_36)begin
        img_reg_array_34_20_real <= _zz_106;
      end
      if(_zz_37)begin
        img_reg_array_35_20_real <= _zz_106;
      end
      if(_zz_38)begin
        img_reg_array_36_20_real <= _zz_106;
      end
      if(_zz_39)begin
        img_reg_array_37_20_real <= _zz_106;
      end
      if(_zz_40)begin
        img_reg_array_38_20_real <= _zz_106;
      end
      if(_zz_41)begin
        img_reg_array_39_20_real <= _zz_106;
      end
      if(_zz_42)begin
        img_reg_array_40_20_real <= _zz_106;
      end
      if(_zz_43)begin
        img_reg_array_41_20_real <= _zz_106;
      end
      if(_zz_44)begin
        img_reg_array_42_20_real <= _zz_106;
      end
      if(_zz_45)begin
        img_reg_array_43_20_real <= _zz_106;
      end
      if(_zz_46)begin
        img_reg_array_44_20_real <= _zz_106;
      end
      if(_zz_47)begin
        img_reg_array_45_20_real <= _zz_106;
      end
      if(_zz_48)begin
        img_reg_array_46_20_real <= _zz_106;
      end
      if(_zz_49)begin
        img_reg_array_47_20_real <= _zz_106;
      end
      if(_zz_50)begin
        img_reg_array_48_20_real <= _zz_106;
      end
      if(_zz_51)begin
        img_reg_array_49_20_real <= _zz_106;
      end
      if(_zz_52)begin
        img_reg_array_50_20_real <= _zz_106;
      end
      if(_zz_53)begin
        img_reg_array_51_20_real <= _zz_106;
      end
      if(_zz_54)begin
        img_reg_array_52_20_real <= _zz_106;
      end
      if(_zz_55)begin
        img_reg_array_53_20_real <= _zz_106;
      end
      if(_zz_56)begin
        img_reg_array_54_20_real <= _zz_106;
      end
      if(_zz_57)begin
        img_reg_array_55_20_real <= _zz_106;
      end
      if(_zz_58)begin
        img_reg_array_56_20_real <= _zz_106;
      end
      if(_zz_59)begin
        img_reg_array_57_20_real <= _zz_106;
      end
      if(_zz_60)begin
        img_reg_array_58_20_real <= _zz_106;
      end
      if(_zz_61)begin
        img_reg_array_59_20_real <= _zz_106;
      end
      if(_zz_62)begin
        img_reg_array_60_20_real <= _zz_106;
      end
      if(_zz_63)begin
        img_reg_array_61_20_real <= _zz_106;
      end
      if(_zz_64)begin
        img_reg_array_62_20_real <= _zz_106;
      end
      if(_zz_65)begin
        img_reg_array_63_20_real <= _zz_106;
      end
      if(_zz_2)begin
        img_reg_array_0_20_imag <= _zz_107;
      end
      if(_zz_3)begin
        img_reg_array_1_20_imag <= _zz_107;
      end
      if(_zz_4)begin
        img_reg_array_2_20_imag <= _zz_107;
      end
      if(_zz_5)begin
        img_reg_array_3_20_imag <= _zz_107;
      end
      if(_zz_6)begin
        img_reg_array_4_20_imag <= _zz_107;
      end
      if(_zz_7)begin
        img_reg_array_5_20_imag <= _zz_107;
      end
      if(_zz_8)begin
        img_reg_array_6_20_imag <= _zz_107;
      end
      if(_zz_9)begin
        img_reg_array_7_20_imag <= _zz_107;
      end
      if(_zz_10)begin
        img_reg_array_8_20_imag <= _zz_107;
      end
      if(_zz_11)begin
        img_reg_array_9_20_imag <= _zz_107;
      end
      if(_zz_12)begin
        img_reg_array_10_20_imag <= _zz_107;
      end
      if(_zz_13)begin
        img_reg_array_11_20_imag <= _zz_107;
      end
      if(_zz_14)begin
        img_reg_array_12_20_imag <= _zz_107;
      end
      if(_zz_15)begin
        img_reg_array_13_20_imag <= _zz_107;
      end
      if(_zz_16)begin
        img_reg_array_14_20_imag <= _zz_107;
      end
      if(_zz_17)begin
        img_reg_array_15_20_imag <= _zz_107;
      end
      if(_zz_18)begin
        img_reg_array_16_20_imag <= _zz_107;
      end
      if(_zz_19)begin
        img_reg_array_17_20_imag <= _zz_107;
      end
      if(_zz_20)begin
        img_reg_array_18_20_imag <= _zz_107;
      end
      if(_zz_21)begin
        img_reg_array_19_20_imag <= _zz_107;
      end
      if(_zz_22)begin
        img_reg_array_20_20_imag <= _zz_107;
      end
      if(_zz_23)begin
        img_reg_array_21_20_imag <= _zz_107;
      end
      if(_zz_24)begin
        img_reg_array_22_20_imag <= _zz_107;
      end
      if(_zz_25)begin
        img_reg_array_23_20_imag <= _zz_107;
      end
      if(_zz_26)begin
        img_reg_array_24_20_imag <= _zz_107;
      end
      if(_zz_27)begin
        img_reg_array_25_20_imag <= _zz_107;
      end
      if(_zz_28)begin
        img_reg_array_26_20_imag <= _zz_107;
      end
      if(_zz_29)begin
        img_reg_array_27_20_imag <= _zz_107;
      end
      if(_zz_30)begin
        img_reg_array_28_20_imag <= _zz_107;
      end
      if(_zz_31)begin
        img_reg_array_29_20_imag <= _zz_107;
      end
      if(_zz_32)begin
        img_reg_array_30_20_imag <= _zz_107;
      end
      if(_zz_33)begin
        img_reg_array_31_20_imag <= _zz_107;
      end
      if(_zz_34)begin
        img_reg_array_32_20_imag <= _zz_107;
      end
      if(_zz_35)begin
        img_reg_array_33_20_imag <= _zz_107;
      end
      if(_zz_36)begin
        img_reg_array_34_20_imag <= _zz_107;
      end
      if(_zz_37)begin
        img_reg_array_35_20_imag <= _zz_107;
      end
      if(_zz_38)begin
        img_reg_array_36_20_imag <= _zz_107;
      end
      if(_zz_39)begin
        img_reg_array_37_20_imag <= _zz_107;
      end
      if(_zz_40)begin
        img_reg_array_38_20_imag <= _zz_107;
      end
      if(_zz_41)begin
        img_reg_array_39_20_imag <= _zz_107;
      end
      if(_zz_42)begin
        img_reg_array_40_20_imag <= _zz_107;
      end
      if(_zz_43)begin
        img_reg_array_41_20_imag <= _zz_107;
      end
      if(_zz_44)begin
        img_reg_array_42_20_imag <= _zz_107;
      end
      if(_zz_45)begin
        img_reg_array_43_20_imag <= _zz_107;
      end
      if(_zz_46)begin
        img_reg_array_44_20_imag <= _zz_107;
      end
      if(_zz_47)begin
        img_reg_array_45_20_imag <= _zz_107;
      end
      if(_zz_48)begin
        img_reg_array_46_20_imag <= _zz_107;
      end
      if(_zz_49)begin
        img_reg_array_47_20_imag <= _zz_107;
      end
      if(_zz_50)begin
        img_reg_array_48_20_imag <= _zz_107;
      end
      if(_zz_51)begin
        img_reg_array_49_20_imag <= _zz_107;
      end
      if(_zz_52)begin
        img_reg_array_50_20_imag <= _zz_107;
      end
      if(_zz_53)begin
        img_reg_array_51_20_imag <= _zz_107;
      end
      if(_zz_54)begin
        img_reg_array_52_20_imag <= _zz_107;
      end
      if(_zz_55)begin
        img_reg_array_53_20_imag <= _zz_107;
      end
      if(_zz_56)begin
        img_reg_array_54_20_imag <= _zz_107;
      end
      if(_zz_57)begin
        img_reg_array_55_20_imag <= _zz_107;
      end
      if(_zz_58)begin
        img_reg_array_56_20_imag <= _zz_107;
      end
      if(_zz_59)begin
        img_reg_array_57_20_imag <= _zz_107;
      end
      if(_zz_60)begin
        img_reg_array_58_20_imag <= _zz_107;
      end
      if(_zz_61)begin
        img_reg_array_59_20_imag <= _zz_107;
      end
      if(_zz_62)begin
        img_reg_array_60_20_imag <= _zz_107;
      end
      if(_zz_63)begin
        img_reg_array_61_20_imag <= _zz_107;
      end
      if(_zz_64)begin
        img_reg_array_62_20_imag <= _zz_107;
      end
      if(_zz_65)begin
        img_reg_array_63_20_imag <= _zz_107;
      end
      if(_zz_2)begin
        img_reg_array_0_21_real <= _zz_108;
      end
      if(_zz_3)begin
        img_reg_array_1_21_real <= _zz_108;
      end
      if(_zz_4)begin
        img_reg_array_2_21_real <= _zz_108;
      end
      if(_zz_5)begin
        img_reg_array_3_21_real <= _zz_108;
      end
      if(_zz_6)begin
        img_reg_array_4_21_real <= _zz_108;
      end
      if(_zz_7)begin
        img_reg_array_5_21_real <= _zz_108;
      end
      if(_zz_8)begin
        img_reg_array_6_21_real <= _zz_108;
      end
      if(_zz_9)begin
        img_reg_array_7_21_real <= _zz_108;
      end
      if(_zz_10)begin
        img_reg_array_8_21_real <= _zz_108;
      end
      if(_zz_11)begin
        img_reg_array_9_21_real <= _zz_108;
      end
      if(_zz_12)begin
        img_reg_array_10_21_real <= _zz_108;
      end
      if(_zz_13)begin
        img_reg_array_11_21_real <= _zz_108;
      end
      if(_zz_14)begin
        img_reg_array_12_21_real <= _zz_108;
      end
      if(_zz_15)begin
        img_reg_array_13_21_real <= _zz_108;
      end
      if(_zz_16)begin
        img_reg_array_14_21_real <= _zz_108;
      end
      if(_zz_17)begin
        img_reg_array_15_21_real <= _zz_108;
      end
      if(_zz_18)begin
        img_reg_array_16_21_real <= _zz_108;
      end
      if(_zz_19)begin
        img_reg_array_17_21_real <= _zz_108;
      end
      if(_zz_20)begin
        img_reg_array_18_21_real <= _zz_108;
      end
      if(_zz_21)begin
        img_reg_array_19_21_real <= _zz_108;
      end
      if(_zz_22)begin
        img_reg_array_20_21_real <= _zz_108;
      end
      if(_zz_23)begin
        img_reg_array_21_21_real <= _zz_108;
      end
      if(_zz_24)begin
        img_reg_array_22_21_real <= _zz_108;
      end
      if(_zz_25)begin
        img_reg_array_23_21_real <= _zz_108;
      end
      if(_zz_26)begin
        img_reg_array_24_21_real <= _zz_108;
      end
      if(_zz_27)begin
        img_reg_array_25_21_real <= _zz_108;
      end
      if(_zz_28)begin
        img_reg_array_26_21_real <= _zz_108;
      end
      if(_zz_29)begin
        img_reg_array_27_21_real <= _zz_108;
      end
      if(_zz_30)begin
        img_reg_array_28_21_real <= _zz_108;
      end
      if(_zz_31)begin
        img_reg_array_29_21_real <= _zz_108;
      end
      if(_zz_32)begin
        img_reg_array_30_21_real <= _zz_108;
      end
      if(_zz_33)begin
        img_reg_array_31_21_real <= _zz_108;
      end
      if(_zz_34)begin
        img_reg_array_32_21_real <= _zz_108;
      end
      if(_zz_35)begin
        img_reg_array_33_21_real <= _zz_108;
      end
      if(_zz_36)begin
        img_reg_array_34_21_real <= _zz_108;
      end
      if(_zz_37)begin
        img_reg_array_35_21_real <= _zz_108;
      end
      if(_zz_38)begin
        img_reg_array_36_21_real <= _zz_108;
      end
      if(_zz_39)begin
        img_reg_array_37_21_real <= _zz_108;
      end
      if(_zz_40)begin
        img_reg_array_38_21_real <= _zz_108;
      end
      if(_zz_41)begin
        img_reg_array_39_21_real <= _zz_108;
      end
      if(_zz_42)begin
        img_reg_array_40_21_real <= _zz_108;
      end
      if(_zz_43)begin
        img_reg_array_41_21_real <= _zz_108;
      end
      if(_zz_44)begin
        img_reg_array_42_21_real <= _zz_108;
      end
      if(_zz_45)begin
        img_reg_array_43_21_real <= _zz_108;
      end
      if(_zz_46)begin
        img_reg_array_44_21_real <= _zz_108;
      end
      if(_zz_47)begin
        img_reg_array_45_21_real <= _zz_108;
      end
      if(_zz_48)begin
        img_reg_array_46_21_real <= _zz_108;
      end
      if(_zz_49)begin
        img_reg_array_47_21_real <= _zz_108;
      end
      if(_zz_50)begin
        img_reg_array_48_21_real <= _zz_108;
      end
      if(_zz_51)begin
        img_reg_array_49_21_real <= _zz_108;
      end
      if(_zz_52)begin
        img_reg_array_50_21_real <= _zz_108;
      end
      if(_zz_53)begin
        img_reg_array_51_21_real <= _zz_108;
      end
      if(_zz_54)begin
        img_reg_array_52_21_real <= _zz_108;
      end
      if(_zz_55)begin
        img_reg_array_53_21_real <= _zz_108;
      end
      if(_zz_56)begin
        img_reg_array_54_21_real <= _zz_108;
      end
      if(_zz_57)begin
        img_reg_array_55_21_real <= _zz_108;
      end
      if(_zz_58)begin
        img_reg_array_56_21_real <= _zz_108;
      end
      if(_zz_59)begin
        img_reg_array_57_21_real <= _zz_108;
      end
      if(_zz_60)begin
        img_reg_array_58_21_real <= _zz_108;
      end
      if(_zz_61)begin
        img_reg_array_59_21_real <= _zz_108;
      end
      if(_zz_62)begin
        img_reg_array_60_21_real <= _zz_108;
      end
      if(_zz_63)begin
        img_reg_array_61_21_real <= _zz_108;
      end
      if(_zz_64)begin
        img_reg_array_62_21_real <= _zz_108;
      end
      if(_zz_65)begin
        img_reg_array_63_21_real <= _zz_108;
      end
      if(_zz_2)begin
        img_reg_array_0_21_imag <= _zz_109;
      end
      if(_zz_3)begin
        img_reg_array_1_21_imag <= _zz_109;
      end
      if(_zz_4)begin
        img_reg_array_2_21_imag <= _zz_109;
      end
      if(_zz_5)begin
        img_reg_array_3_21_imag <= _zz_109;
      end
      if(_zz_6)begin
        img_reg_array_4_21_imag <= _zz_109;
      end
      if(_zz_7)begin
        img_reg_array_5_21_imag <= _zz_109;
      end
      if(_zz_8)begin
        img_reg_array_6_21_imag <= _zz_109;
      end
      if(_zz_9)begin
        img_reg_array_7_21_imag <= _zz_109;
      end
      if(_zz_10)begin
        img_reg_array_8_21_imag <= _zz_109;
      end
      if(_zz_11)begin
        img_reg_array_9_21_imag <= _zz_109;
      end
      if(_zz_12)begin
        img_reg_array_10_21_imag <= _zz_109;
      end
      if(_zz_13)begin
        img_reg_array_11_21_imag <= _zz_109;
      end
      if(_zz_14)begin
        img_reg_array_12_21_imag <= _zz_109;
      end
      if(_zz_15)begin
        img_reg_array_13_21_imag <= _zz_109;
      end
      if(_zz_16)begin
        img_reg_array_14_21_imag <= _zz_109;
      end
      if(_zz_17)begin
        img_reg_array_15_21_imag <= _zz_109;
      end
      if(_zz_18)begin
        img_reg_array_16_21_imag <= _zz_109;
      end
      if(_zz_19)begin
        img_reg_array_17_21_imag <= _zz_109;
      end
      if(_zz_20)begin
        img_reg_array_18_21_imag <= _zz_109;
      end
      if(_zz_21)begin
        img_reg_array_19_21_imag <= _zz_109;
      end
      if(_zz_22)begin
        img_reg_array_20_21_imag <= _zz_109;
      end
      if(_zz_23)begin
        img_reg_array_21_21_imag <= _zz_109;
      end
      if(_zz_24)begin
        img_reg_array_22_21_imag <= _zz_109;
      end
      if(_zz_25)begin
        img_reg_array_23_21_imag <= _zz_109;
      end
      if(_zz_26)begin
        img_reg_array_24_21_imag <= _zz_109;
      end
      if(_zz_27)begin
        img_reg_array_25_21_imag <= _zz_109;
      end
      if(_zz_28)begin
        img_reg_array_26_21_imag <= _zz_109;
      end
      if(_zz_29)begin
        img_reg_array_27_21_imag <= _zz_109;
      end
      if(_zz_30)begin
        img_reg_array_28_21_imag <= _zz_109;
      end
      if(_zz_31)begin
        img_reg_array_29_21_imag <= _zz_109;
      end
      if(_zz_32)begin
        img_reg_array_30_21_imag <= _zz_109;
      end
      if(_zz_33)begin
        img_reg_array_31_21_imag <= _zz_109;
      end
      if(_zz_34)begin
        img_reg_array_32_21_imag <= _zz_109;
      end
      if(_zz_35)begin
        img_reg_array_33_21_imag <= _zz_109;
      end
      if(_zz_36)begin
        img_reg_array_34_21_imag <= _zz_109;
      end
      if(_zz_37)begin
        img_reg_array_35_21_imag <= _zz_109;
      end
      if(_zz_38)begin
        img_reg_array_36_21_imag <= _zz_109;
      end
      if(_zz_39)begin
        img_reg_array_37_21_imag <= _zz_109;
      end
      if(_zz_40)begin
        img_reg_array_38_21_imag <= _zz_109;
      end
      if(_zz_41)begin
        img_reg_array_39_21_imag <= _zz_109;
      end
      if(_zz_42)begin
        img_reg_array_40_21_imag <= _zz_109;
      end
      if(_zz_43)begin
        img_reg_array_41_21_imag <= _zz_109;
      end
      if(_zz_44)begin
        img_reg_array_42_21_imag <= _zz_109;
      end
      if(_zz_45)begin
        img_reg_array_43_21_imag <= _zz_109;
      end
      if(_zz_46)begin
        img_reg_array_44_21_imag <= _zz_109;
      end
      if(_zz_47)begin
        img_reg_array_45_21_imag <= _zz_109;
      end
      if(_zz_48)begin
        img_reg_array_46_21_imag <= _zz_109;
      end
      if(_zz_49)begin
        img_reg_array_47_21_imag <= _zz_109;
      end
      if(_zz_50)begin
        img_reg_array_48_21_imag <= _zz_109;
      end
      if(_zz_51)begin
        img_reg_array_49_21_imag <= _zz_109;
      end
      if(_zz_52)begin
        img_reg_array_50_21_imag <= _zz_109;
      end
      if(_zz_53)begin
        img_reg_array_51_21_imag <= _zz_109;
      end
      if(_zz_54)begin
        img_reg_array_52_21_imag <= _zz_109;
      end
      if(_zz_55)begin
        img_reg_array_53_21_imag <= _zz_109;
      end
      if(_zz_56)begin
        img_reg_array_54_21_imag <= _zz_109;
      end
      if(_zz_57)begin
        img_reg_array_55_21_imag <= _zz_109;
      end
      if(_zz_58)begin
        img_reg_array_56_21_imag <= _zz_109;
      end
      if(_zz_59)begin
        img_reg_array_57_21_imag <= _zz_109;
      end
      if(_zz_60)begin
        img_reg_array_58_21_imag <= _zz_109;
      end
      if(_zz_61)begin
        img_reg_array_59_21_imag <= _zz_109;
      end
      if(_zz_62)begin
        img_reg_array_60_21_imag <= _zz_109;
      end
      if(_zz_63)begin
        img_reg_array_61_21_imag <= _zz_109;
      end
      if(_zz_64)begin
        img_reg_array_62_21_imag <= _zz_109;
      end
      if(_zz_65)begin
        img_reg_array_63_21_imag <= _zz_109;
      end
      if(_zz_2)begin
        img_reg_array_0_22_real <= _zz_110;
      end
      if(_zz_3)begin
        img_reg_array_1_22_real <= _zz_110;
      end
      if(_zz_4)begin
        img_reg_array_2_22_real <= _zz_110;
      end
      if(_zz_5)begin
        img_reg_array_3_22_real <= _zz_110;
      end
      if(_zz_6)begin
        img_reg_array_4_22_real <= _zz_110;
      end
      if(_zz_7)begin
        img_reg_array_5_22_real <= _zz_110;
      end
      if(_zz_8)begin
        img_reg_array_6_22_real <= _zz_110;
      end
      if(_zz_9)begin
        img_reg_array_7_22_real <= _zz_110;
      end
      if(_zz_10)begin
        img_reg_array_8_22_real <= _zz_110;
      end
      if(_zz_11)begin
        img_reg_array_9_22_real <= _zz_110;
      end
      if(_zz_12)begin
        img_reg_array_10_22_real <= _zz_110;
      end
      if(_zz_13)begin
        img_reg_array_11_22_real <= _zz_110;
      end
      if(_zz_14)begin
        img_reg_array_12_22_real <= _zz_110;
      end
      if(_zz_15)begin
        img_reg_array_13_22_real <= _zz_110;
      end
      if(_zz_16)begin
        img_reg_array_14_22_real <= _zz_110;
      end
      if(_zz_17)begin
        img_reg_array_15_22_real <= _zz_110;
      end
      if(_zz_18)begin
        img_reg_array_16_22_real <= _zz_110;
      end
      if(_zz_19)begin
        img_reg_array_17_22_real <= _zz_110;
      end
      if(_zz_20)begin
        img_reg_array_18_22_real <= _zz_110;
      end
      if(_zz_21)begin
        img_reg_array_19_22_real <= _zz_110;
      end
      if(_zz_22)begin
        img_reg_array_20_22_real <= _zz_110;
      end
      if(_zz_23)begin
        img_reg_array_21_22_real <= _zz_110;
      end
      if(_zz_24)begin
        img_reg_array_22_22_real <= _zz_110;
      end
      if(_zz_25)begin
        img_reg_array_23_22_real <= _zz_110;
      end
      if(_zz_26)begin
        img_reg_array_24_22_real <= _zz_110;
      end
      if(_zz_27)begin
        img_reg_array_25_22_real <= _zz_110;
      end
      if(_zz_28)begin
        img_reg_array_26_22_real <= _zz_110;
      end
      if(_zz_29)begin
        img_reg_array_27_22_real <= _zz_110;
      end
      if(_zz_30)begin
        img_reg_array_28_22_real <= _zz_110;
      end
      if(_zz_31)begin
        img_reg_array_29_22_real <= _zz_110;
      end
      if(_zz_32)begin
        img_reg_array_30_22_real <= _zz_110;
      end
      if(_zz_33)begin
        img_reg_array_31_22_real <= _zz_110;
      end
      if(_zz_34)begin
        img_reg_array_32_22_real <= _zz_110;
      end
      if(_zz_35)begin
        img_reg_array_33_22_real <= _zz_110;
      end
      if(_zz_36)begin
        img_reg_array_34_22_real <= _zz_110;
      end
      if(_zz_37)begin
        img_reg_array_35_22_real <= _zz_110;
      end
      if(_zz_38)begin
        img_reg_array_36_22_real <= _zz_110;
      end
      if(_zz_39)begin
        img_reg_array_37_22_real <= _zz_110;
      end
      if(_zz_40)begin
        img_reg_array_38_22_real <= _zz_110;
      end
      if(_zz_41)begin
        img_reg_array_39_22_real <= _zz_110;
      end
      if(_zz_42)begin
        img_reg_array_40_22_real <= _zz_110;
      end
      if(_zz_43)begin
        img_reg_array_41_22_real <= _zz_110;
      end
      if(_zz_44)begin
        img_reg_array_42_22_real <= _zz_110;
      end
      if(_zz_45)begin
        img_reg_array_43_22_real <= _zz_110;
      end
      if(_zz_46)begin
        img_reg_array_44_22_real <= _zz_110;
      end
      if(_zz_47)begin
        img_reg_array_45_22_real <= _zz_110;
      end
      if(_zz_48)begin
        img_reg_array_46_22_real <= _zz_110;
      end
      if(_zz_49)begin
        img_reg_array_47_22_real <= _zz_110;
      end
      if(_zz_50)begin
        img_reg_array_48_22_real <= _zz_110;
      end
      if(_zz_51)begin
        img_reg_array_49_22_real <= _zz_110;
      end
      if(_zz_52)begin
        img_reg_array_50_22_real <= _zz_110;
      end
      if(_zz_53)begin
        img_reg_array_51_22_real <= _zz_110;
      end
      if(_zz_54)begin
        img_reg_array_52_22_real <= _zz_110;
      end
      if(_zz_55)begin
        img_reg_array_53_22_real <= _zz_110;
      end
      if(_zz_56)begin
        img_reg_array_54_22_real <= _zz_110;
      end
      if(_zz_57)begin
        img_reg_array_55_22_real <= _zz_110;
      end
      if(_zz_58)begin
        img_reg_array_56_22_real <= _zz_110;
      end
      if(_zz_59)begin
        img_reg_array_57_22_real <= _zz_110;
      end
      if(_zz_60)begin
        img_reg_array_58_22_real <= _zz_110;
      end
      if(_zz_61)begin
        img_reg_array_59_22_real <= _zz_110;
      end
      if(_zz_62)begin
        img_reg_array_60_22_real <= _zz_110;
      end
      if(_zz_63)begin
        img_reg_array_61_22_real <= _zz_110;
      end
      if(_zz_64)begin
        img_reg_array_62_22_real <= _zz_110;
      end
      if(_zz_65)begin
        img_reg_array_63_22_real <= _zz_110;
      end
      if(_zz_2)begin
        img_reg_array_0_22_imag <= _zz_111;
      end
      if(_zz_3)begin
        img_reg_array_1_22_imag <= _zz_111;
      end
      if(_zz_4)begin
        img_reg_array_2_22_imag <= _zz_111;
      end
      if(_zz_5)begin
        img_reg_array_3_22_imag <= _zz_111;
      end
      if(_zz_6)begin
        img_reg_array_4_22_imag <= _zz_111;
      end
      if(_zz_7)begin
        img_reg_array_5_22_imag <= _zz_111;
      end
      if(_zz_8)begin
        img_reg_array_6_22_imag <= _zz_111;
      end
      if(_zz_9)begin
        img_reg_array_7_22_imag <= _zz_111;
      end
      if(_zz_10)begin
        img_reg_array_8_22_imag <= _zz_111;
      end
      if(_zz_11)begin
        img_reg_array_9_22_imag <= _zz_111;
      end
      if(_zz_12)begin
        img_reg_array_10_22_imag <= _zz_111;
      end
      if(_zz_13)begin
        img_reg_array_11_22_imag <= _zz_111;
      end
      if(_zz_14)begin
        img_reg_array_12_22_imag <= _zz_111;
      end
      if(_zz_15)begin
        img_reg_array_13_22_imag <= _zz_111;
      end
      if(_zz_16)begin
        img_reg_array_14_22_imag <= _zz_111;
      end
      if(_zz_17)begin
        img_reg_array_15_22_imag <= _zz_111;
      end
      if(_zz_18)begin
        img_reg_array_16_22_imag <= _zz_111;
      end
      if(_zz_19)begin
        img_reg_array_17_22_imag <= _zz_111;
      end
      if(_zz_20)begin
        img_reg_array_18_22_imag <= _zz_111;
      end
      if(_zz_21)begin
        img_reg_array_19_22_imag <= _zz_111;
      end
      if(_zz_22)begin
        img_reg_array_20_22_imag <= _zz_111;
      end
      if(_zz_23)begin
        img_reg_array_21_22_imag <= _zz_111;
      end
      if(_zz_24)begin
        img_reg_array_22_22_imag <= _zz_111;
      end
      if(_zz_25)begin
        img_reg_array_23_22_imag <= _zz_111;
      end
      if(_zz_26)begin
        img_reg_array_24_22_imag <= _zz_111;
      end
      if(_zz_27)begin
        img_reg_array_25_22_imag <= _zz_111;
      end
      if(_zz_28)begin
        img_reg_array_26_22_imag <= _zz_111;
      end
      if(_zz_29)begin
        img_reg_array_27_22_imag <= _zz_111;
      end
      if(_zz_30)begin
        img_reg_array_28_22_imag <= _zz_111;
      end
      if(_zz_31)begin
        img_reg_array_29_22_imag <= _zz_111;
      end
      if(_zz_32)begin
        img_reg_array_30_22_imag <= _zz_111;
      end
      if(_zz_33)begin
        img_reg_array_31_22_imag <= _zz_111;
      end
      if(_zz_34)begin
        img_reg_array_32_22_imag <= _zz_111;
      end
      if(_zz_35)begin
        img_reg_array_33_22_imag <= _zz_111;
      end
      if(_zz_36)begin
        img_reg_array_34_22_imag <= _zz_111;
      end
      if(_zz_37)begin
        img_reg_array_35_22_imag <= _zz_111;
      end
      if(_zz_38)begin
        img_reg_array_36_22_imag <= _zz_111;
      end
      if(_zz_39)begin
        img_reg_array_37_22_imag <= _zz_111;
      end
      if(_zz_40)begin
        img_reg_array_38_22_imag <= _zz_111;
      end
      if(_zz_41)begin
        img_reg_array_39_22_imag <= _zz_111;
      end
      if(_zz_42)begin
        img_reg_array_40_22_imag <= _zz_111;
      end
      if(_zz_43)begin
        img_reg_array_41_22_imag <= _zz_111;
      end
      if(_zz_44)begin
        img_reg_array_42_22_imag <= _zz_111;
      end
      if(_zz_45)begin
        img_reg_array_43_22_imag <= _zz_111;
      end
      if(_zz_46)begin
        img_reg_array_44_22_imag <= _zz_111;
      end
      if(_zz_47)begin
        img_reg_array_45_22_imag <= _zz_111;
      end
      if(_zz_48)begin
        img_reg_array_46_22_imag <= _zz_111;
      end
      if(_zz_49)begin
        img_reg_array_47_22_imag <= _zz_111;
      end
      if(_zz_50)begin
        img_reg_array_48_22_imag <= _zz_111;
      end
      if(_zz_51)begin
        img_reg_array_49_22_imag <= _zz_111;
      end
      if(_zz_52)begin
        img_reg_array_50_22_imag <= _zz_111;
      end
      if(_zz_53)begin
        img_reg_array_51_22_imag <= _zz_111;
      end
      if(_zz_54)begin
        img_reg_array_52_22_imag <= _zz_111;
      end
      if(_zz_55)begin
        img_reg_array_53_22_imag <= _zz_111;
      end
      if(_zz_56)begin
        img_reg_array_54_22_imag <= _zz_111;
      end
      if(_zz_57)begin
        img_reg_array_55_22_imag <= _zz_111;
      end
      if(_zz_58)begin
        img_reg_array_56_22_imag <= _zz_111;
      end
      if(_zz_59)begin
        img_reg_array_57_22_imag <= _zz_111;
      end
      if(_zz_60)begin
        img_reg_array_58_22_imag <= _zz_111;
      end
      if(_zz_61)begin
        img_reg_array_59_22_imag <= _zz_111;
      end
      if(_zz_62)begin
        img_reg_array_60_22_imag <= _zz_111;
      end
      if(_zz_63)begin
        img_reg_array_61_22_imag <= _zz_111;
      end
      if(_zz_64)begin
        img_reg_array_62_22_imag <= _zz_111;
      end
      if(_zz_65)begin
        img_reg_array_63_22_imag <= _zz_111;
      end
      if(_zz_2)begin
        img_reg_array_0_23_real <= _zz_112;
      end
      if(_zz_3)begin
        img_reg_array_1_23_real <= _zz_112;
      end
      if(_zz_4)begin
        img_reg_array_2_23_real <= _zz_112;
      end
      if(_zz_5)begin
        img_reg_array_3_23_real <= _zz_112;
      end
      if(_zz_6)begin
        img_reg_array_4_23_real <= _zz_112;
      end
      if(_zz_7)begin
        img_reg_array_5_23_real <= _zz_112;
      end
      if(_zz_8)begin
        img_reg_array_6_23_real <= _zz_112;
      end
      if(_zz_9)begin
        img_reg_array_7_23_real <= _zz_112;
      end
      if(_zz_10)begin
        img_reg_array_8_23_real <= _zz_112;
      end
      if(_zz_11)begin
        img_reg_array_9_23_real <= _zz_112;
      end
      if(_zz_12)begin
        img_reg_array_10_23_real <= _zz_112;
      end
      if(_zz_13)begin
        img_reg_array_11_23_real <= _zz_112;
      end
      if(_zz_14)begin
        img_reg_array_12_23_real <= _zz_112;
      end
      if(_zz_15)begin
        img_reg_array_13_23_real <= _zz_112;
      end
      if(_zz_16)begin
        img_reg_array_14_23_real <= _zz_112;
      end
      if(_zz_17)begin
        img_reg_array_15_23_real <= _zz_112;
      end
      if(_zz_18)begin
        img_reg_array_16_23_real <= _zz_112;
      end
      if(_zz_19)begin
        img_reg_array_17_23_real <= _zz_112;
      end
      if(_zz_20)begin
        img_reg_array_18_23_real <= _zz_112;
      end
      if(_zz_21)begin
        img_reg_array_19_23_real <= _zz_112;
      end
      if(_zz_22)begin
        img_reg_array_20_23_real <= _zz_112;
      end
      if(_zz_23)begin
        img_reg_array_21_23_real <= _zz_112;
      end
      if(_zz_24)begin
        img_reg_array_22_23_real <= _zz_112;
      end
      if(_zz_25)begin
        img_reg_array_23_23_real <= _zz_112;
      end
      if(_zz_26)begin
        img_reg_array_24_23_real <= _zz_112;
      end
      if(_zz_27)begin
        img_reg_array_25_23_real <= _zz_112;
      end
      if(_zz_28)begin
        img_reg_array_26_23_real <= _zz_112;
      end
      if(_zz_29)begin
        img_reg_array_27_23_real <= _zz_112;
      end
      if(_zz_30)begin
        img_reg_array_28_23_real <= _zz_112;
      end
      if(_zz_31)begin
        img_reg_array_29_23_real <= _zz_112;
      end
      if(_zz_32)begin
        img_reg_array_30_23_real <= _zz_112;
      end
      if(_zz_33)begin
        img_reg_array_31_23_real <= _zz_112;
      end
      if(_zz_34)begin
        img_reg_array_32_23_real <= _zz_112;
      end
      if(_zz_35)begin
        img_reg_array_33_23_real <= _zz_112;
      end
      if(_zz_36)begin
        img_reg_array_34_23_real <= _zz_112;
      end
      if(_zz_37)begin
        img_reg_array_35_23_real <= _zz_112;
      end
      if(_zz_38)begin
        img_reg_array_36_23_real <= _zz_112;
      end
      if(_zz_39)begin
        img_reg_array_37_23_real <= _zz_112;
      end
      if(_zz_40)begin
        img_reg_array_38_23_real <= _zz_112;
      end
      if(_zz_41)begin
        img_reg_array_39_23_real <= _zz_112;
      end
      if(_zz_42)begin
        img_reg_array_40_23_real <= _zz_112;
      end
      if(_zz_43)begin
        img_reg_array_41_23_real <= _zz_112;
      end
      if(_zz_44)begin
        img_reg_array_42_23_real <= _zz_112;
      end
      if(_zz_45)begin
        img_reg_array_43_23_real <= _zz_112;
      end
      if(_zz_46)begin
        img_reg_array_44_23_real <= _zz_112;
      end
      if(_zz_47)begin
        img_reg_array_45_23_real <= _zz_112;
      end
      if(_zz_48)begin
        img_reg_array_46_23_real <= _zz_112;
      end
      if(_zz_49)begin
        img_reg_array_47_23_real <= _zz_112;
      end
      if(_zz_50)begin
        img_reg_array_48_23_real <= _zz_112;
      end
      if(_zz_51)begin
        img_reg_array_49_23_real <= _zz_112;
      end
      if(_zz_52)begin
        img_reg_array_50_23_real <= _zz_112;
      end
      if(_zz_53)begin
        img_reg_array_51_23_real <= _zz_112;
      end
      if(_zz_54)begin
        img_reg_array_52_23_real <= _zz_112;
      end
      if(_zz_55)begin
        img_reg_array_53_23_real <= _zz_112;
      end
      if(_zz_56)begin
        img_reg_array_54_23_real <= _zz_112;
      end
      if(_zz_57)begin
        img_reg_array_55_23_real <= _zz_112;
      end
      if(_zz_58)begin
        img_reg_array_56_23_real <= _zz_112;
      end
      if(_zz_59)begin
        img_reg_array_57_23_real <= _zz_112;
      end
      if(_zz_60)begin
        img_reg_array_58_23_real <= _zz_112;
      end
      if(_zz_61)begin
        img_reg_array_59_23_real <= _zz_112;
      end
      if(_zz_62)begin
        img_reg_array_60_23_real <= _zz_112;
      end
      if(_zz_63)begin
        img_reg_array_61_23_real <= _zz_112;
      end
      if(_zz_64)begin
        img_reg_array_62_23_real <= _zz_112;
      end
      if(_zz_65)begin
        img_reg_array_63_23_real <= _zz_112;
      end
      if(_zz_2)begin
        img_reg_array_0_23_imag <= _zz_113;
      end
      if(_zz_3)begin
        img_reg_array_1_23_imag <= _zz_113;
      end
      if(_zz_4)begin
        img_reg_array_2_23_imag <= _zz_113;
      end
      if(_zz_5)begin
        img_reg_array_3_23_imag <= _zz_113;
      end
      if(_zz_6)begin
        img_reg_array_4_23_imag <= _zz_113;
      end
      if(_zz_7)begin
        img_reg_array_5_23_imag <= _zz_113;
      end
      if(_zz_8)begin
        img_reg_array_6_23_imag <= _zz_113;
      end
      if(_zz_9)begin
        img_reg_array_7_23_imag <= _zz_113;
      end
      if(_zz_10)begin
        img_reg_array_8_23_imag <= _zz_113;
      end
      if(_zz_11)begin
        img_reg_array_9_23_imag <= _zz_113;
      end
      if(_zz_12)begin
        img_reg_array_10_23_imag <= _zz_113;
      end
      if(_zz_13)begin
        img_reg_array_11_23_imag <= _zz_113;
      end
      if(_zz_14)begin
        img_reg_array_12_23_imag <= _zz_113;
      end
      if(_zz_15)begin
        img_reg_array_13_23_imag <= _zz_113;
      end
      if(_zz_16)begin
        img_reg_array_14_23_imag <= _zz_113;
      end
      if(_zz_17)begin
        img_reg_array_15_23_imag <= _zz_113;
      end
      if(_zz_18)begin
        img_reg_array_16_23_imag <= _zz_113;
      end
      if(_zz_19)begin
        img_reg_array_17_23_imag <= _zz_113;
      end
      if(_zz_20)begin
        img_reg_array_18_23_imag <= _zz_113;
      end
      if(_zz_21)begin
        img_reg_array_19_23_imag <= _zz_113;
      end
      if(_zz_22)begin
        img_reg_array_20_23_imag <= _zz_113;
      end
      if(_zz_23)begin
        img_reg_array_21_23_imag <= _zz_113;
      end
      if(_zz_24)begin
        img_reg_array_22_23_imag <= _zz_113;
      end
      if(_zz_25)begin
        img_reg_array_23_23_imag <= _zz_113;
      end
      if(_zz_26)begin
        img_reg_array_24_23_imag <= _zz_113;
      end
      if(_zz_27)begin
        img_reg_array_25_23_imag <= _zz_113;
      end
      if(_zz_28)begin
        img_reg_array_26_23_imag <= _zz_113;
      end
      if(_zz_29)begin
        img_reg_array_27_23_imag <= _zz_113;
      end
      if(_zz_30)begin
        img_reg_array_28_23_imag <= _zz_113;
      end
      if(_zz_31)begin
        img_reg_array_29_23_imag <= _zz_113;
      end
      if(_zz_32)begin
        img_reg_array_30_23_imag <= _zz_113;
      end
      if(_zz_33)begin
        img_reg_array_31_23_imag <= _zz_113;
      end
      if(_zz_34)begin
        img_reg_array_32_23_imag <= _zz_113;
      end
      if(_zz_35)begin
        img_reg_array_33_23_imag <= _zz_113;
      end
      if(_zz_36)begin
        img_reg_array_34_23_imag <= _zz_113;
      end
      if(_zz_37)begin
        img_reg_array_35_23_imag <= _zz_113;
      end
      if(_zz_38)begin
        img_reg_array_36_23_imag <= _zz_113;
      end
      if(_zz_39)begin
        img_reg_array_37_23_imag <= _zz_113;
      end
      if(_zz_40)begin
        img_reg_array_38_23_imag <= _zz_113;
      end
      if(_zz_41)begin
        img_reg_array_39_23_imag <= _zz_113;
      end
      if(_zz_42)begin
        img_reg_array_40_23_imag <= _zz_113;
      end
      if(_zz_43)begin
        img_reg_array_41_23_imag <= _zz_113;
      end
      if(_zz_44)begin
        img_reg_array_42_23_imag <= _zz_113;
      end
      if(_zz_45)begin
        img_reg_array_43_23_imag <= _zz_113;
      end
      if(_zz_46)begin
        img_reg_array_44_23_imag <= _zz_113;
      end
      if(_zz_47)begin
        img_reg_array_45_23_imag <= _zz_113;
      end
      if(_zz_48)begin
        img_reg_array_46_23_imag <= _zz_113;
      end
      if(_zz_49)begin
        img_reg_array_47_23_imag <= _zz_113;
      end
      if(_zz_50)begin
        img_reg_array_48_23_imag <= _zz_113;
      end
      if(_zz_51)begin
        img_reg_array_49_23_imag <= _zz_113;
      end
      if(_zz_52)begin
        img_reg_array_50_23_imag <= _zz_113;
      end
      if(_zz_53)begin
        img_reg_array_51_23_imag <= _zz_113;
      end
      if(_zz_54)begin
        img_reg_array_52_23_imag <= _zz_113;
      end
      if(_zz_55)begin
        img_reg_array_53_23_imag <= _zz_113;
      end
      if(_zz_56)begin
        img_reg_array_54_23_imag <= _zz_113;
      end
      if(_zz_57)begin
        img_reg_array_55_23_imag <= _zz_113;
      end
      if(_zz_58)begin
        img_reg_array_56_23_imag <= _zz_113;
      end
      if(_zz_59)begin
        img_reg_array_57_23_imag <= _zz_113;
      end
      if(_zz_60)begin
        img_reg_array_58_23_imag <= _zz_113;
      end
      if(_zz_61)begin
        img_reg_array_59_23_imag <= _zz_113;
      end
      if(_zz_62)begin
        img_reg_array_60_23_imag <= _zz_113;
      end
      if(_zz_63)begin
        img_reg_array_61_23_imag <= _zz_113;
      end
      if(_zz_64)begin
        img_reg_array_62_23_imag <= _zz_113;
      end
      if(_zz_65)begin
        img_reg_array_63_23_imag <= _zz_113;
      end
      if(_zz_2)begin
        img_reg_array_0_24_real <= _zz_114;
      end
      if(_zz_3)begin
        img_reg_array_1_24_real <= _zz_114;
      end
      if(_zz_4)begin
        img_reg_array_2_24_real <= _zz_114;
      end
      if(_zz_5)begin
        img_reg_array_3_24_real <= _zz_114;
      end
      if(_zz_6)begin
        img_reg_array_4_24_real <= _zz_114;
      end
      if(_zz_7)begin
        img_reg_array_5_24_real <= _zz_114;
      end
      if(_zz_8)begin
        img_reg_array_6_24_real <= _zz_114;
      end
      if(_zz_9)begin
        img_reg_array_7_24_real <= _zz_114;
      end
      if(_zz_10)begin
        img_reg_array_8_24_real <= _zz_114;
      end
      if(_zz_11)begin
        img_reg_array_9_24_real <= _zz_114;
      end
      if(_zz_12)begin
        img_reg_array_10_24_real <= _zz_114;
      end
      if(_zz_13)begin
        img_reg_array_11_24_real <= _zz_114;
      end
      if(_zz_14)begin
        img_reg_array_12_24_real <= _zz_114;
      end
      if(_zz_15)begin
        img_reg_array_13_24_real <= _zz_114;
      end
      if(_zz_16)begin
        img_reg_array_14_24_real <= _zz_114;
      end
      if(_zz_17)begin
        img_reg_array_15_24_real <= _zz_114;
      end
      if(_zz_18)begin
        img_reg_array_16_24_real <= _zz_114;
      end
      if(_zz_19)begin
        img_reg_array_17_24_real <= _zz_114;
      end
      if(_zz_20)begin
        img_reg_array_18_24_real <= _zz_114;
      end
      if(_zz_21)begin
        img_reg_array_19_24_real <= _zz_114;
      end
      if(_zz_22)begin
        img_reg_array_20_24_real <= _zz_114;
      end
      if(_zz_23)begin
        img_reg_array_21_24_real <= _zz_114;
      end
      if(_zz_24)begin
        img_reg_array_22_24_real <= _zz_114;
      end
      if(_zz_25)begin
        img_reg_array_23_24_real <= _zz_114;
      end
      if(_zz_26)begin
        img_reg_array_24_24_real <= _zz_114;
      end
      if(_zz_27)begin
        img_reg_array_25_24_real <= _zz_114;
      end
      if(_zz_28)begin
        img_reg_array_26_24_real <= _zz_114;
      end
      if(_zz_29)begin
        img_reg_array_27_24_real <= _zz_114;
      end
      if(_zz_30)begin
        img_reg_array_28_24_real <= _zz_114;
      end
      if(_zz_31)begin
        img_reg_array_29_24_real <= _zz_114;
      end
      if(_zz_32)begin
        img_reg_array_30_24_real <= _zz_114;
      end
      if(_zz_33)begin
        img_reg_array_31_24_real <= _zz_114;
      end
      if(_zz_34)begin
        img_reg_array_32_24_real <= _zz_114;
      end
      if(_zz_35)begin
        img_reg_array_33_24_real <= _zz_114;
      end
      if(_zz_36)begin
        img_reg_array_34_24_real <= _zz_114;
      end
      if(_zz_37)begin
        img_reg_array_35_24_real <= _zz_114;
      end
      if(_zz_38)begin
        img_reg_array_36_24_real <= _zz_114;
      end
      if(_zz_39)begin
        img_reg_array_37_24_real <= _zz_114;
      end
      if(_zz_40)begin
        img_reg_array_38_24_real <= _zz_114;
      end
      if(_zz_41)begin
        img_reg_array_39_24_real <= _zz_114;
      end
      if(_zz_42)begin
        img_reg_array_40_24_real <= _zz_114;
      end
      if(_zz_43)begin
        img_reg_array_41_24_real <= _zz_114;
      end
      if(_zz_44)begin
        img_reg_array_42_24_real <= _zz_114;
      end
      if(_zz_45)begin
        img_reg_array_43_24_real <= _zz_114;
      end
      if(_zz_46)begin
        img_reg_array_44_24_real <= _zz_114;
      end
      if(_zz_47)begin
        img_reg_array_45_24_real <= _zz_114;
      end
      if(_zz_48)begin
        img_reg_array_46_24_real <= _zz_114;
      end
      if(_zz_49)begin
        img_reg_array_47_24_real <= _zz_114;
      end
      if(_zz_50)begin
        img_reg_array_48_24_real <= _zz_114;
      end
      if(_zz_51)begin
        img_reg_array_49_24_real <= _zz_114;
      end
      if(_zz_52)begin
        img_reg_array_50_24_real <= _zz_114;
      end
      if(_zz_53)begin
        img_reg_array_51_24_real <= _zz_114;
      end
      if(_zz_54)begin
        img_reg_array_52_24_real <= _zz_114;
      end
      if(_zz_55)begin
        img_reg_array_53_24_real <= _zz_114;
      end
      if(_zz_56)begin
        img_reg_array_54_24_real <= _zz_114;
      end
      if(_zz_57)begin
        img_reg_array_55_24_real <= _zz_114;
      end
      if(_zz_58)begin
        img_reg_array_56_24_real <= _zz_114;
      end
      if(_zz_59)begin
        img_reg_array_57_24_real <= _zz_114;
      end
      if(_zz_60)begin
        img_reg_array_58_24_real <= _zz_114;
      end
      if(_zz_61)begin
        img_reg_array_59_24_real <= _zz_114;
      end
      if(_zz_62)begin
        img_reg_array_60_24_real <= _zz_114;
      end
      if(_zz_63)begin
        img_reg_array_61_24_real <= _zz_114;
      end
      if(_zz_64)begin
        img_reg_array_62_24_real <= _zz_114;
      end
      if(_zz_65)begin
        img_reg_array_63_24_real <= _zz_114;
      end
      if(_zz_2)begin
        img_reg_array_0_24_imag <= _zz_115;
      end
      if(_zz_3)begin
        img_reg_array_1_24_imag <= _zz_115;
      end
      if(_zz_4)begin
        img_reg_array_2_24_imag <= _zz_115;
      end
      if(_zz_5)begin
        img_reg_array_3_24_imag <= _zz_115;
      end
      if(_zz_6)begin
        img_reg_array_4_24_imag <= _zz_115;
      end
      if(_zz_7)begin
        img_reg_array_5_24_imag <= _zz_115;
      end
      if(_zz_8)begin
        img_reg_array_6_24_imag <= _zz_115;
      end
      if(_zz_9)begin
        img_reg_array_7_24_imag <= _zz_115;
      end
      if(_zz_10)begin
        img_reg_array_8_24_imag <= _zz_115;
      end
      if(_zz_11)begin
        img_reg_array_9_24_imag <= _zz_115;
      end
      if(_zz_12)begin
        img_reg_array_10_24_imag <= _zz_115;
      end
      if(_zz_13)begin
        img_reg_array_11_24_imag <= _zz_115;
      end
      if(_zz_14)begin
        img_reg_array_12_24_imag <= _zz_115;
      end
      if(_zz_15)begin
        img_reg_array_13_24_imag <= _zz_115;
      end
      if(_zz_16)begin
        img_reg_array_14_24_imag <= _zz_115;
      end
      if(_zz_17)begin
        img_reg_array_15_24_imag <= _zz_115;
      end
      if(_zz_18)begin
        img_reg_array_16_24_imag <= _zz_115;
      end
      if(_zz_19)begin
        img_reg_array_17_24_imag <= _zz_115;
      end
      if(_zz_20)begin
        img_reg_array_18_24_imag <= _zz_115;
      end
      if(_zz_21)begin
        img_reg_array_19_24_imag <= _zz_115;
      end
      if(_zz_22)begin
        img_reg_array_20_24_imag <= _zz_115;
      end
      if(_zz_23)begin
        img_reg_array_21_24_imag <= _zz_115;
      end
      if(_zz_24)begin
        img_reg_array_22_24_imag <= _zz_115;
      end
      if(_zz_25)begin
        img_reg_array_23_24_imag <= _zz_115;
      end
      if(_zz_26)begin
        img_reg_array_24_24_imag <= _zz_115;
      end
      if(_zz_27)begin
        img_reg_array_25_24_imag <= _zz_115;
      end
      if(_zz_28)begin
        img_reg_array_26_24_imag <= _zz_115;
      end
      if(_zz_29)begin
        img_reg_array_27_24_imag <= _zz_115;
      end
      if(_zz_30)begin
        img_reg_array_28_24_imag <= _zz_115;
      end
      if(_zz_31)begin
        img_reg_array_29_24_imag <= _zz_115;
      end
      if(_zz_32)begin
        img_reg_array_30_24_imag <= _zz_115;
      end
      if(_zz_33)begin
        img_reg_array_31_24_imag <= _zz_115;
      end
      if(_zz_34)begin
        img_reg_array_32_24_imag <= _zz_115;
      end
      if(_zz_35)begin
        img_reg_array_33_24_imag <= _zz_115;
      end
      if(_zz_36)begin
        img_reg_array_34_24_imag <= _zz_115;
      end
      if(_zz_37)begin
        img_reg_array_35_24_imag <= _zz_115;
      end
      if(_zz_38)begin
        img_reg_array_36_24_imag <= _zz_115;
      end
      if(_zz_39)begin
        img_reg_array_37_24_imag <= _zz_115;
      end
      if(_zz_40)begin
        img_reg_array_38_24_imag <= _zz_115;
      end
      if(_zz_41)begin
        img_reg_array_39_24_imag <= _zz_115;
      end
      if(_zz_42)begin
        img_reg_array_40_24_imag <= _zz_115;
      end
      if(_zz_43)begin
        img_reg_array_41_24_imag <= _zz_115;
      end
      if(_zz_44)begin
        img_reg_array_42_24_imag <= _zz_115;
      end
      if(_zz_45)begin
        img_reg_array_43_24_imag <= _zz_115;
      end
      if(_zz_46)begin
        img_reg_array_44_24_imag <= _zz_115;
      end
      if(_zz_47)begin
        img_reg_array_45_24_imag <= _zz_115;
      end
      if(_zz_48)begin
        img_reg_array_46_24_imag <= _zz_115;
      end
      if(_zz_49)begin
        img_reg_array_47_24_imag <= _zz_115;
      end
      if(_zz_50)begin
        img_reg_array_48_24_imag <= _zz_115;
      end
      if(_zz_51)begin
        img_reg_array_49_24_imag <= _zz_115;
      end
      if(_zz_52)begin
        img_reg_array_50_24_imag <= _zz_115;
      end
      if(_zz_53)begin
        img_reg_array_51_24_imag <= _zz_115;
      end
      if(_zz_54)begin
        img_reg_array_52_24_imag <= _zz_115;
      end
      if(_zz_55)begin
        img_reg_array_53_24_imag <= _zz_115;
      end
      if(_zz_56)begin
        img_reg_array_54_24_imag <= _zz_115;
      end
      if(_zz_57)begin
        img_reg_array_55_24_imag <= _zz_115;
      end
      if(_zz_58)begin
        img_reg_array_56_24_imag <= _zz_115;
      end
      if(_zz_59)begin
        img_reg_array_57_24_imag <= _zz_115;
      end
      if(_zz_60)begin
        img_reg_array_58_24_imag <= _zz_115;
      end
      if(_zz_61)begin
        img_reg_array_59_24_imag <= _zz_115;
      end
      if(_zz_62)begin
        img_reg_array_60_24_imag <= _zz_115;
      end
      if(_zz_63)begin
        img_reg_array_61_24_imag <= _zz_115;
      end
      if(_zz_64)begin
        img_reg_array_62_24_imag <= _zz_115;
      end
      if(_zz_65)begin
        img_reg_array_63_24_imag <= _zz_115;
      end
      if(_zz_2)begin
        img_reg_array_0_25_real <= _zz_116;
      end
      if(_zz_3)begin
        img_reg_array_1_25_real <= _zz_116;
      end
      if(_zz_4)begin
        img_reg_array_2_25_real <= _zz_116;
      end
      if(_zz_5)begin
        img_reg_array_3_25_real <= _zz_116;
      end
      if(_zz_6)begin
        img_reg_array_4_25_real <= _zz_116;
      end
      if(_zz_7)begin
        img_reg_array_5_25_real <= _zz_116;
      end
      if(_zz_8)begin
        img_reg_array_6_25_real <= _zz_116;
      end
      if(_zz_9)begin
        img_reg_array_7_25_real <= _zz_116;
      end
      if(_zz_10)begin
        img_reg_array_8_25_real <= _zz_116;
      end
      if(_zz_11)begin
        img_reg_array_9_25_real <= _zz_116;
      end
      if(_zz_12)begin
        img_reg_array_10_25_real <= _zz_116;
      end
      if(_zz_13)begin
        img_reg_array_11_25_real <= _zz_116;
      end
      if(_zz_14)begin
        img_reg_array_12_25_real <= _zz_116;
      end
      if(_zz_15)begin
        img_reg_array_13_25_real <= _zz_116;
      end
      if(_zz_16)begin
        img_reg_array_14_25_real <= _zz_116;
      end
      if(_zz_17)begin
        img_reg_array_15_25_real <= _zz_116;
      end
      if(_zz_18)begin
        img_reg_array_16_25_real <= _zz_116;
      end
      if(_zz_19)begin
        img_reg_array_17_25_real <= _zz_116;
      end
      if(_zz_20)begin
        img_reg_array_18_25_real <= _zz_116;
      end
      if(_zz_21)begin
        img_reg_array_19_25_real <= _zz_116;
      end
      if(_zz_22)begin
        img_reg_array_20_25_real <= _zz_116;
      end
      if(_zz_23)begin
        img_reg_array_21_25_real <= _zz_116;
      end
      if(_zz_24)begin
        img_reg_array_22_25_real <= _zz_116;
      end
      if(_zz_25)begin
        img_reg_array_23_25_real <= _zz_116;
      end
      if(_zz_26)begin
        img_reg_array_24_25_real <= _zz_116;
      end
      if(_zz_27)begin
        img_reg_array_25_25_real <= _zz_116;
      end
      if(_zz_28)begin
        img_reg_array_26_25_real <= _zz_116;
      end
      if(_zz_29)begin
        img_reg_array_27_25_real <= _zz_116;
      end
      if(_zz_30)begin
        img_reg_array_28_25_real <= _zz_116;
      end
      if(_zz_31)begin
        img_reg_array_29_25_real <= _zz_116;
      end
      if(_zz_32)begin
        img_reg_array_30_25_real <= _zz_116;
      end
      if(_zz_33)begin
        img_reg_array_31_25_real <= _zz_116;
      end
      if(_zz_34)begin
        img_reg_array_32_25_real <= _zz_116;
      end
      if(_zz_35)begin
        img_reg_array_33_25_real <= _zz_116;
      end
      if(_zz_36)begin
        img_reg_array_34_25_real <= _zz_116;
      end
      if(_zz_37)begin
        img_reg_array_35_25_real <= _zz_116;
      end
      if(_zz_38)begin
        img_reg_array_36_25_real <= _zz_116;
      end
      if(_zz_39)begin
        img_reg_array_37_25_real <= _zz_116;
      end
      if(_zz_40)begin
        img_reg_array_38_25_real <= _zz_116;
      end
      if(_zz_41)begin
        img_reg_array_39_25_real <= _zz_116;
      end
      if(_zz_42)begin
        img_reg_array_40_25_real <= _zz_116;
      end
      if(_zz_43)begin
        img_reg_array_41_25_real <= _zz_116;
      end
      if(_zz_44)begin
        img_reg_array_42_25_real <= _zz_116;
      end
      if(_zz_45)begin
        img_reg_array_43_25_real <= _zz_116;
      end
      if(_zz_46)begin
        img_reg_array_44_25_real <= _zz_116;
      end
      if(_zz_47)begin
        img_reg_array_45_25_real <= _zz_116;
      end
      if(_zz_48)begin
        img_reg_array_46_25_real <= _zz_116;
      end
      if(_zz_49)begin
        img_reg_array_47_25_real <= _zz_116;
      end
      if(_zz_50)begin
        img_reg_array_48_25_real <= _zz_116;
      end
      if(_zz_51)begin
        img_reg_array_49_25_real <= _zz_116;
      end
      if(_zz_52)begin
        img_reg_array_50_25_real <= _zz_116;
      end
      if(_zz_53)begin
        img_reg_array_51_25_real <= _zz_116;
      end
      if(_zz_54)begin
        img_reg_array_52_25_real <= _zz_116;
      end
      if(_zz_55)begin
        img_reg_array_53_25_real <= _zz_116;
      end
      if(_zz_56)begin
        img_reg_array_54_25_real <= _zz_116;
      end
      if(_zz_57)begin
        img_reg_array_55_25_real <= _zz_116;
      end
      if(_zz_58)begin
        img_reg_array_56_25_real <= _zz_116;
      end
      if(_zz_59)begin
        img_reg_array_57_25_real <= _zz_116;
      end
      if(_zz_60)begin
        img_reg_array_58_25_real <= _zz_116;
      end
      if(_zz_61)begin
        img_reg_array_59_25_real <= _zz_116;
      end
      if(_zz_62)begin
        img_reg_array_60_25_real <= _zz_116;
      end
      if(_zz_63)begin
        img_reg_array_61_25_real <= _zz_116;
      end
      if(_zz_64)begin
        img_reg_array_62_25_real <= _zz_116;
      end
      if(_zz_65)begin
        img_reg_array_63_25_real <= _zz_116;
      end
      if(_zz_2)begin
        img_reg_array_0_25_imag <= _zz_117;
      end
      if(_zz_3)begin
        img_reg_array_1_25_imag <= _zz_117;
      end
      if(_zz_4)begin
        img_reg_array_2_25_imag <= _zz_117;
      end
      if(_zz_5)begin
        img_reg_array_3_25_imag <= _zz_117;
      end
      if(_zz_6)begin
        img_reg_array_4_25_imag <= _zz_117;
      end
      if(_zz_7)begin
        img_reg_array_5_25_imag <= _zz_117;
      end
      if(_zz_8)begin
        img_reg_array_6_25_imag <= _zz_117;
      end
      if(_zz_9)begin
        img_reg_array_7_25_imag <= _zz_117;
      end
      if(_zz_10)begin
        img_reg_array_8_25_imag <= _zz_117;
      end
      if(_zz_11)begin
        img_reg_array_9_25_imag <= _zz_117;
      end
      if(_zz_12)begin
        img_reg_array_10_25_imag <= _zz_117;
      end
      if(_zz_13)begin
        img_reg_array_11_25_imag <= _zz_117;
      end
      if(_zz_14)begin
        img_reg_array_12_25_imag <= _zz_117;
      end
      if(_zz_15)begin
        img_reg_array_13_25_imag <= _zz_117;
      end
      if(_zz_16)begin
        img_reg_array_14_25_imag <= _zz_117;
      end
      if(_zz_17)begin
        img_reg_array_15_25_imag <= _zz_117;
      end
      if(_zz_18)begin
        img_reg_array_16_25_imag <= _zz_117;
      end
      if(_zz_19)begin
        img_reg_array_17_25_imag <= _zz_117;
      end
      if(_zz_20)begin
        img_reg_array_18_25_imag <= _zz_117;
      end
      if(_zz_21)begin
        img_reg_array_19_25_imag <= _zz_117;
      end
      if(_zz_22)begin
        img_reg_array_20_25_imag <= _zz_117;
      end
      if(_zz_23)begin
        img_reg_array_21_25_imag <= _zz_117;
      end
      if(_zz_24)begin
        img_reg_array_22_25_imag <= _zz_117;
      end
      if(_zz_25)begin
        img_reg_array_23_25_imag <= _zz_117;
      end
      if(_zz_26)begin
        img_reg_array_24_25_imag <= _zz_117;
      end
      if(_zz_27)begin
        img_reg_array_25_25_imag <= _zz_117;
      end
      if(_zz_28)begin
        img_reg_array_26_25_imag <= _zz_117;
      end
      if(_zz_29)begin
        img_reg_array_27_25_imag <= _zz_117;
      end
      if(_zz_30)begin
        img_reg_array_28_25_imag <= _zz_117;
      end
      if(_zz_31)begin
        img_reg_array_29_25_imag <= _zz_117;
      end
      if(_zz_32)begin
        img_reg_array_30_25_imag <= _zz_117;
      end
      if(_zz_33)begin
        img_reg_array_31_25_imag <= _zz_117;
      end
      if(_zz_34)begin
        img_reg_array_32_25_imag <= _zz_117;
      end
      if(_zz_35)begin
        img_reg_array_33_25_imag <= _zz_117;
      end
      if(_zz_36)begin
        img_reg_array_34_25_imag <= _zz_117;
      end
      if(_zz_37)begin
        img_reg_array_35_25_imag <= _zz_117;
      end
      if(_zz_38)begin
        img_reg_array_36_25_imag <= _zz_117;
      end
      if(_zz_39)begin
        img_reg_array_37_25_imag <= _zz_117;
      end
      if(_zz_40)begin
        img_reg_array_38_25_imag <= _zz_117;
      end
      if(_zz_41)begin
        img_reg_array_39_25_imag <= _zz_117;
      end
      if(_zz_42)begin
        img_reg_array_40_25_imag <= _zz_117;
      end
      if(_zz_43)begin
        img_reg_array_41_25_imag <= _zz_117;
      end
      if(_zz_44)begin
        img_reg_array_42_25_imag <= _zz_117;
      end
      if(_zz_45)begin
        img_reg_array_43_25_imag <= _zz_117;
      end
      if(_zz_46)begin
        img_reg_array_44_25_imag <= _zz_117;
      end
      if(_zz_47)begin
        img_reg_array_45_25_imag <= _zz_117;
      end
      if(_zz_48)begin
        img_reg_array_46_25_imag <= _zz_117;
      end
      if(_zz_49)begin
        img_reg_array_47_25_imag <= _zz_117;
      end
      if(_zz_50)begin
        img_reg_array_48_25_imag <= _zz_117;
      end
      if(_zz_51)begin
        img_reg_array_49_25_imag <= _zz_117;
      end
      if(_zz_52)begin
        img_reg_array_50_25_imag <= _zz_117;
      end
      if(_zz_53)begin
        img_reg_array_51_25_imag <= _zz_117;
      end
      if(_zz_54)begin
        img_reg_array_52_25_imag <= _zz_117;
      end
      if(_zz_55)begin
        img_reg_array_53_25_imag <= _zz_117;
      end
      if(_zz_56)begin
        img_reg_array_54_25_imag <= _zz_117;
      end
      if(_zz_57)begin
        img_reg_array_55_25_imag <= _zz_117;
      end
      if(_zz_58)begin
        img_reg_array_56_25_imag <= _zz_117;
      end
      if(_zz_59)begin
        img_reg_array_57_25_imag <= _zz_117;
      end
      if(_zz_60)begin
        img_reg_array_58_25_imag <= _zz_117;
      end
      if(_zz_61)begin
        img_reg_array_59_25_imag <= _zz_117;
      end
      if(_zz_62)begin
        img_reg_array_60_25_imag <= _zz_117;
      end
      if(_zz_63)begin
        img_reg_array_61_25_imag <= _zz_117;
      end
      if(_zz_64)begin
        img_reg_array_62_25_imag <= _zz_117;
      end
      if(_zz_65)begin
        img_reg_array_63_25_imag <= _zz_117;
      end
      if(_zz_2)begin
        img_reg_array_0_26_real <= _zz_118;
      end
      if(_zz_3)begin
        img_reg_array_1_26_real <= _zz_118;
      end
      if(_zz_4)begin
        img_reg_array_2_26_real <= _zz_118;
      end
      if(_zz_5)begin
        img_reg_array_3_26_real <= _zz_118;
      end
      if(_zz_6)begin
        img_reg_array_4_26_real <= _zz_118;
      end
      if(_zz_7)begin
        img_reg_array_5_26_real <= _zz_118;
      end
      if(_zz_8)begin
        img_reg_array_6_26_real <= _zz_118;
      end
      if(_zz_9)begin
        img_reg_array_7_26_real <= _zz_118;
      end
      if(_zz_10)begin
        img_reg_array_8_26_real <= _zz_118;
      end
      if(_zz_11)begin
        img_reg_array_9_26_real <= _zz_118;
      end
      if(_zz_12)begin
        img_reg_array_10_26_real <= _zz_118;
      end
      if(_zz_13)begin
        img_reg_array_11_26_real <= _zz_118;
      end
      if(_zz_14)begin
        img_reg_array_12_26_real <= _zz_118;
      end
      if(_zz_15)begin
        img_reg_array_13_26_real <= _zz_118;
      end
      if(_zz_16)begin
        img_reg_array_14_26_real <= _zz_118;
      end
      if(_zz_17)begin
        img_reg_array_15_26_real <= _zz_118;
      end
      if(_zz_18)begin
        img_reg_array_16_26_real <= _zz_118;
      end
      if(_zz_19)begin
        img_reg_array_17_26_real <= _zz_118;
      end
      if(_zz_20)begin
        img_reg_array_18_26_real <= _zz_118;
      end
      if(_zz_21)begin
        img_reg_array_19_26_real <= _zz_118;
      end
      if(_zz_22)begin
        img_reg_array_20_26_real <= _zz_118;
      end
      if(_zz_23)begin
        img_reg_array_21_26_real <= _zz_118;
      end
      if(_zz_24)begin
        img_reg_array_22_26_real <= _zz_118;
      end
      if(_zz_25)begin
        img_reg_array_23_26_real <= _zz_118;
      end
      if(_zz_26)begin
        img_reg_array_24_26_real <= _zz_118;
      end
      if(_zz_27)begin
        img_reg_array_25_26_real <= _zz_118;
      end
      if(_zz_28)begin
        img_reg_array_26_26_real <= _zz_118;
      end
      if(_zz_29)begin
        img_reg_array_27_26_real <= _zz_118;
      end
      if(_zz_30)begin
        img_reg_array_28_26_real <= _zz_118;
      end
      if(_zz_31)begin
        img_reg_array_29_26_real <= _zz_118;
      end
      if(_zz_32)begin
        img_reg_array_30_26_real <= _zz_118;
      end
      if(_zz_33)begin
        img_reg_array_31_26_real <= _zz_118;
      end
      if(_zz_34)begin
        img_reg_array_32_26_real <= _zz_118;
      end
      if(_zz_35)begin
        img_reg_array_33_26_real <= _zz_118;
      end
      if(_zz_36)begin
        img_reg_array_34_26_real <= _zz_118;
      end
      if(_zz_37)begin
        img_reg_array_35_26_real <= _zz_118;
      end
      if(_zz_38)begin
        img_reg_array_36_26_real <= _zz_118;
      end
      if(_zz_39)begin
        img_reg_array_37_26_real <= _zz_118;
      end
      if(_zz_40)begin
        img_reg_array_38_26_real <= _zz_118;
      end
      if(_zz_41)begin
        img_reg_array_39_26_real <= _zz_118;
      end
      if(_zz_42)begin
        img_reg_array_40_26_real <= _zz_118;
      end
      if(_zz_43)begin
        img_reg_array_41_26_real <= _zz_118;
      end
      if(_zz_44)begin
        img_reg_array_42_26_real <= _zz_118;
      end
      if(_zz_45)begin
        img_reg_array_43_26_real <= _zz_118;
      end
      if(_zz_46)begin
        img_reg_array_44_26_real <= _zz_118;
      end
      if(_zz_47)begin
        img_reg_array_45_26_real <= _zz_118;
      end
      if(_zz_48)begin
        img_reg_array_46_26_real <= _zz_118;
      end
      if(_zz_49)begin
        img_reg_array_47_26_real <= _zz_118;
      end
      if(_zz_50)begin
        img_reg_array_48_26_real <= _zz_118;
      end
      if(_zz_51)begin
        img_reg_array_49_26_real <= _zz_118;
      end
      if(_zz_52)begin
        img_reg_array_50_26_real <= _zz_118;
      end
      if(_zz_53)begin
        img_reg_array_51_26_real <= _zz_118;
      end
      if(_zz_54)begin
        img_reg_array_52_26_real <= _zz_118;
      end
      if(_zz_55)begin
        img_reg_array_53_26_real <= _zz_118;
      end
      if(_zz_56)begin
        img_reg_array_54_26_real <= _zz_118;
      end
      if(_zz_57)begin
        img_reg_array_55_26_real <= _zz_118;
      end
      if(_zz_58)begin
        img_reg_array_56_26_real <= _zz_118;
      end
      if(_zz_59)begin
        img_reg_array_57_26_real <= _zz_118;
      end
      if(_zz_60)begin
        img_reg_array_58_26_real <= _zz_118;
      end
      if(_zz_61)begin
        img_reg_array_59_26_real <= _zz_118;
      end
      if(_zz_62)begin
        img_reg_array_60_26_real <= _zz_118;
      end
      if(_zz_63)begin
        img_reg_array_61_26_real <= _zz_118;
      end
      if(_zz_64)begin
        img_reg_array_62_26_real <= _zz_118;
      end
      if(_zz_65)begin
        img_reg_array_63_26_real <= _zz_118;
      end
      if(_zz_2)begin
        img_reg_array_0_26_imag <= _zz_119;
      end
      if(_zz_3)begin
        img_reg_array_1_26_imag <= _zz_119;
      end
      if(_zz_4)begin
        img_reg_array_2_26_imag <= _zz_119;
      end
      if(_zz_5)begin
        img_reg_array_3_26_imag <= _zz_119;
      end
      if(_zz_6)begin
        img_reg_array_4_26_imag <= _zz_119;
      end
      if(_zz_7)begin
        img_reg_array_5_26_imag <= _zz_119;
      end
      if(_zz_8)begin
        img_reg_array_6_26_imag <= _zz_119;
      end
      if(_zz_9)begin
        img_reg_array_7_26_imag <= _zz_119;
      end
      if(_zz_10)begin
        img_reg_array_8_26_imag <= _zz_119;
      end
      if(_zz_11)begin
        img_reg_array_9_26_imag <= _zz_119;
      end
      if(_zz_12)begin
        img_reg_array_10_26_imag <= _zz_119;
      end
      if(_zz_13)begin
        img_reg_array_11_26_imag <= _zz_119;
      end
      if(_zz_14)begin
        img_reg_array_12_26_imag <= _zz_119;
      end
      if(_zz_15)begin
        img_reg_array_13_26_imag <= _zz_119;
      end
      if(_zz_16)begin
        img_reg_array_14_26_imag <= _zz_119;
      end
      if(_zz_17)begin
        img_reg_array_15_26_imag <= _zz_119;
      end
      if(_zz_18)begin
        img_reg_array_16_26_imag <= _zz_119;
      end
      if(_zz_19)begin
        img_reg_array_17_26_imag <= _zz_119;
      end
      if(_zz_20)begin
        img_reg_array_18_26_imag <= _zz_119;
      end
      if(_zz_21)begin
        img_reg_array_19_26_imag <= _zz_119;
      end
      if(_zz_22)begin
        img_reg_array_20_26_imag <= _zz_119;
      end
      if(_zz_23)begin
        img_reg_array_21_26_imag <= _zz_119;
      end
      if(_zz_24)begin
        img_reg_array_22_26_imag <= _zz_119;
      end
      if(_zz_25)begin
        img_reg_array_23_26_imag <= _zz_119;
      end
      if(_zz_26)begin
        img_reg_array_24_26_imag <= _zz_119;
      end
      if(_zz_27)begin
        img_reg_array_25_26_imag <= _zz_119;
      end
      if(_zz_28)begin
        img_reg_array_26_26_imag <= _zz_119;
      end
      if(_zz_29)begin
        img_reg_array_27_26_imag <= _zz_119;
      end
      if(_zz_30)begin
        img_reg_array_28_26_imag <= _zz_119;
      end
      if(_zz_31)begin
        img_reg_array_29_26_imag <= _zz_119;
      end
      if(_zz_32)begin
        img_reg_array_30_26_imag <= _zz_119;
      end
      if(_zz_33)begin
        img_reg_array_31_26_imag <= _zz_119;
      end
      if(_zz_34)begin
        img_reg_array_32_26_imag <= _zz_119;
      end
      if(_zz_35)begin
        img_reg_array_33_26_imag <= _zz_119;
      end
      if(_zz_36)begin
        img_reg_array_34_26_imag <= _zz_119;
      end
      if(_zz_37)begin
        img_reg_array_35_26_imag <= _zz_119;
      end
      if(_zz_38)begin
        img_reg_array_36_26_imag <= _zz_119;
      end
      if(_zz_39)begin
        img_reg_array_37_26_imag <= _zz_119;
      end
      if(_zz_40)begin
        img_reg_array_38_26_imag <= _zz_119;
      end
      if(_zz_41)begin
        img_reg_array_39_26_imag <= _zz_119;
      end
      if(_zz_42)begin
        img_reg_array_40_26_imag <= _zz_119;
      end
      if(_zz_43)begin
        img_reg_array_41_26_imag <= _zz_119;
      end
      if(_zz_44)begin
        img_reg_array_42_26_imag <= _zz_119;
      end
      if(_zz_45)begin
        img_reg_array_43_26_imag <= _zz_119;
      end
      if(_zz_46)begin
        img_reg_array_44_26_imag <= _zz_119;
      end
      if(_zz_47)begin
        img_reg_array_45_26_imag <= _zz_119;
      end
      if(_zz_48)begin
        img_reg_array_46_26_imag <= _zz_119;
      end
      if(_zz_49)begin
        img_reg_array_47_26_imag <= _zz_119;
      end
      if(_zz_50)begin
        img_reg_array_48_26_imag <= _zz_119;
      end
      if(_zz_51)begin
        img_reg_array_49_26_imag <= _zz_119;
      end
      if(_zz_52)begin
        img_reg_array_50_26_imag <= _zz_119;
      end
      if(_zz_53)begin
        img_reg_array_51_26_imag <= _zz_119;
      end
      if(_zz_54)begin
        img_reg_array_52_26_imag <= _zz_119;
      end
      if(_zz_55)begin
        img_reg_array_53_26_imag <= _zz_119;
      end
      if(_zz_56)begin
        img_reg_array_54_26_imag <= _zz_119;
      end
      if(_zz_57)begin
        img_reg_array_55_26_imag <= _zz_119;
      end
      if(_zz_58)begin
        img_reg_array_56_26_imag <= _zz_119;
      end
      if(_zz_59)begin
        img_reg_array_57_26_imag <= _zz_119;
      end
      if(_zz_60)begin
        img_reg_array_58_26_imag <= _zz_119;
      end
      if(_zz_61)begin
        img_reg_array_59_26_imag <= _zz_119;
      end
      if(_zz_62)begin
        img_reg_array_60_26_imag <= _zz_119;
      end
      if(_zz_63)begin
        img_reg_array_61_26_imag <= _zz_119;
      end
      if(_zz_64)begin
        img_reg_array_62_26_imag <= _zz_119;
      end
      if(_zz_65)begin
        img_reg_array_63_26_imag <= _zz_119;
      end
      if(_zz_2)begin
        img_reg_array_0_27_real <= _zz_120;
      end
      if(_zz_3)begin
        img_reg_array_1_27_real <= _zz_120;
      end
      if(_zz_4)begin
        img_reg_array_2_27_real <= _zz_120;
      end
      if(_zz_5)begin
        img_reg_array_3_27_real <= _zz_120;
      end
      if(_zz_6)begin
        img_reg_array_4_27_real <= _zz_120;
      end
      if(_zz_7)begin
        img_reg_array_5_27_real <= _zz_120;
      end
      if(_zz_8)begin
        img_reg_array_6_27_real <= _zz_120;
      end
      if(_zz_9)begin
        img_reg_array_7_27_real <= _zz_120;
      end
      if(_zz_10)begin
        img_reg_array_8_27_real <= _zz_120;
      end
      if(_zz_11)begin
        img_reg_array_9_27_real <= _zz_120;
      end
      if(_zz_12)begin
        img_reg_array_10_27_real <= _zz_120;
      end
      if(_zz_13)begin
        img_reg_array_11_27_real <= _zz_120;
      end
      if(_zz_14)begin
        img_reg_array_12_27_real <= _zz_120;
      end
      if(_zz_15)begin
        img_reg_array_13_27_real <= _zz_120;
      end
      if(_zz_16)begin
        img_reg_array_14_27_real <= _zz_120;
      end
      if(_zz_17)begin
        img_reg_array_15_27_real <= _zz_120;
      end
      if(_zz_18)begin
        img_reg_array_16_27_real <= _zz_120;
      end
      if(_zz_19)begin
        img_reg_array_17_27_real <= _zz_120;
      end
      if(_zz_20)begin
        img_reg_array_18_27_real <= _zz_120;
      end
      if(_zz_21)begin
        img_reg_array_19_27_real <= _zz_120;
      end
      if(_zz_22)begin
        img_reg_array_20_27_real <= _zz_120;
      end
      if(_zz_23)begin
        img_reg_array_21_27_real <= _zz_120;
      end
      if(_zz_24)begin
        img_reg_array_22_27_real <= _zz_120;
      end
      if(_zz_25)begin
        img_reg_array_23_27_real <= _zz_120;
      end
      if(_zz_26)begin
        img_reg_array_24_27_real <= _zz_120;
      end
      if(_zz_27)begin
        img_reg_array_25_27_real <= _zz_120;
      end
      if(_zz_28)begin
        img_reg_array_26_27_real <= _zz_120;
      end
      if(_zz_29)begin
        img_reg_array_27_27_real <= _zz_120;
      end
      if(_zz_30)begin
        img_reg_array_28_27_real <= _zz_120;
      end
      if(_zz_31)begin
        img_reg_array_29_27_real <= _zz_120;
      end
      if(_zz_32)begin
        img_reg_array_30_27_real <= _zz_120;
      end
      if(_zz_33)begin
        img_reg_array_31_27_real <= _zz_120;
      end
      if(_zz_34)begin
        img_reg_array_32_27_real <= _zz_120;
      end
      if(_zz_35)begin
        img_reg_array_33_27_real <= _zz_120;
      end
      if(_zz_36)begin
        img_reg_array_34_27_real <= _zz_120;
      end
      if(_zz_37)begin
        img_reg_array_35_27_real <= _zz_120;
      end
      if(_zz_38)begin
        img_reg_array_36_27_real <= _zz_120;
      end
      if(_zz_39)begin
        img_reg_array_37_27_real <= _zz_120;
      end
      if(_zz_40)begin
        img_reg_array_38_27_real <= _zz_120;
      end
      if(_zz_41)begin
        img_reg_array_39_27_real <= _zz_120;
      end
      if(_zz_42)begin
        img_reg_array_40_27_real <= _zz_120;
      end
      if(_zz_43)begin
        img_reg_array_41_27_real <= _zz_120;
      end
      if(_zz_44)begin
        img_reg_array_42_27_real <= _zz_120;
      end
      if(_zz_45)begin
        img_reg_array_43_27_real <= _zz_120;
      end
      if(_zz_46)begin
        img_reg_array_44_27_real <= _zz_120;
      end
      if(_zz_47)begin
        img_reg_array_45_27_real <= _zz_120;
      end
      if(_zz_48)begin
        img_reg_array_46_27_real <= _zz_120;
      end
      if(_zz_49)begin
        img_reg_array_47_27_real <= _zz_120;
      end
      if(_zz_50)begin
        img_reg_array_48_27_real <= _zz_120;
      end
      if(_zz_51)begin
        img_reg_array_49_27_real <= _zz_120;
      end
      if(_zz_52)begin
        img_reg_array_50_27_real <= _zz_120;
      end
      if(_zz_53)begin
        img_reg_array_51_27_real <= _zz_120;
      end
      if(_zz_54)begin
        img_reg_array_52_27_real <= _zz_120;
      end
      if(_zz_55)begin
        img_reg_array_53_27_real <= _zz_120;
      end
      if(_zz_56)begin
        img_reg_array_54_27_real <= _zz_120;
      end
      if(_zz_57)begin
        img_reg_array_55_27_real <= _zz_120;
      end
      if(_zz_58)begin
        img_reg_array_56_27_real <= _zz_120;
      end
      if(_zz_59)begin
        img_reg_array_57_27_real <= _zz_120;
      end
      if(_zz_60)begin
        img_reg_array_58_27_real <= _zz_120;
      end
      if(_zz_61)begin
        img_reg_array_59_27_real <= _zz_120;
      end
      if(_zz_62)begin
        img_reg_array_60_27_real <= _zz_120;
      end
      if(_zz_63)begin
        img_reg_array_61_27_real <= _zz_120;
      end
      if(_zz_64)begin
        img_reg_array_62_27_real <= _zz_120;
      end
      if(_zz_65)begin
        img_reg_array_63_27_real <= _zz_120;
      end
      if(_zz_2)begin
        img_reg_array_0_27_imag <= _zz_121;
      end
      if(_zz_3)begin
        img_reg_array_1_27_imag <= _zz_121;
      end
      if(_zz_4)begin
        img_reg_array_2_27_imag <= _zz_121;
      end
      if(_zz_5)begin
        img_reg_array_3_27_imag <= _zz_121;
      end
      if(_zz_6)begin
        img_reg_array_4_27_imag <= _zz_121;
      end
      if(_zz_7)begin
        img_reg_array_5_27_imag <= _zz_121;
      end
      if(_zz_8)begin
        img_reg_array_6_27_imag <= _zz_121;
      end
      if(_zz_9)begin
        img_reg_array_7_27_imag <= _zz_121;
      end
      if(_zz_10)begin
        img_reg_array_8_27_imag <= _zz_121;
      end
      if(_zz_11)begin
        img_reg_array_9_27_imag <= _zz_121;
      end
      if(_zz_12)begin
        img_reg_array_10_27_imag <= _zz_121;
      end
      if(_zz_13)begin
        img_reg_array_11_27_imag <= _zz_121;
      end
      if(_zz_14)begin
        img_reg_array_12_27_imag <= _zz_121;
      end
      if(_zz_15)begin
        img_reg_array_13_27_imag <= _zz_121;
      end
      if(_zz_16)begin
        img_reg_array_14_27_imag <= _zz_121;
      end
      if(_zz_17)begin
        img_reg_array_15_27_imag <= _zz_121;
      end
      if(_zz_18)begin
        img_reg_array_16_27_imag <= _zz_121;
      end
      if(_zz_19)begin
        img_reg_array_17_27_imag <= _zz_121;
      end
      if(_zz_20)begin
        img_reg_array_18_27_imag <= _zz_121;
      end
      if(_zz_21)begin
        img_reg_array_19_27_imag <= _zz_121;
      end
      if(_zz_22)begin
        img_reg_array_20_27_imag <= _zz_121;
      end
      if(_zz_23)begin
        img_reg_array_21_27_imag <= _zz_121;
      end
      if(_zz_24)begin
        img_reg_array_22_27_imag <= _zz_121;
      end
      if(_zz_25)begin
        img_reg_array_23_27_imag <= _zz_121;
      end
      if(_zz_26)begin
        img_reg_array_24_27_imag <= _zz_121;
      end
      if(_zz_27)begin
        img_reg_array_25_27_imag <= _zz_121;
      end
      if(_zz_28)begin
        img_reg_array_26_27_imag <= _zz_121;
      end
      if(_zz_29)begin
        img_reg_array_27_27_imag <= _zz_121;
      end
      if(_zz_30)begin
        img_reg_array_28_27_imag <= _zz_121;
      end
      if(_zz_31)begin
        img_reg_array_29_27_imag <= _zz_121;
      end
      if(_zz_32)begin
        img_reg_array_30_27_imag <= _zz_121;
      end
      if(_zz_33)begin
        img_reg_array_31_27_imag <= _zz_121;
      end
      if(_zz_34)begin
        img_reg_array_32_27_imag <= _zz_121;
      end
      if(_zz_35)begin
        img_reg_array_33_27_imag <= _zz_121;
      end
      if(_zz_36)begin
        img_reg_array_34_27_imag <= _zz_121;
      end
      if(_zz_37)begin
        img_reg_array_35_27_imag <= _zz_121;
      end
      if(_zz_38)begin
        img_reg_array_36_27_imag <= _zz_121;
      end
      if(_zz_39)begin
        img_reg_array_37_27_imag <= _zz_121;
      end
      if(_zz_40)begin
        img_reg_array_38_27_imag <= _zz_121;
      end
      if(_zz_41)begin
        img_reg_array_39_27_imag <= _zz_121;
      end
      if(_zz_42)begin
        img_reg_array_40_27_imag <= _zz_121;
      end
      if(_zz_43)begin
        img_reg_array_41_27_imag <= _zz_121;
      end
      if(_zz_44)begin
        img_reg_array_42_27_imag <= _zz_121;
      end
      if(_zz_45)begin
        img_reg_array_43_27_imag <= _zz_121;
      end
      if(_zz_46)begin
        img_reg_array_44_27_imag <= _zz_121;
      end
      if(_zz_47)begin
        img_reg_array_45_27_imag <= _zz_121;
      end
      if(_zz_48)begin
        img_reg_array_46_27_imag <= _zz_121;
      end
      if(_zz_49)begin
        img_reg_array_47_27_imag <= _zz_121;
      end
      if(_zz_50)begin
        img_reg_array_48_27_imag <= _zz_121;
      end
      if(_zz_51)begin
        img_reg_array_49_27_imag <= _zz_121;
      end
      if(_zz_52)begin
        img_reg_array_50_27_imag <= _zz_121;
      end
      if(_zz_53)begin
        img_reg_array_51_27_imag <= _zz_121;
      end
      if(_zz_54)begin
        img_reg_array_52_27_imag <= _zz_121;
      end
      if(_zz_55)begin
        img_reg_array_53_27_imag <= _zz_121;
      end
      if(_zz_56)begin
        img_reg_array_54_27_imag <= _zz_121;
      end
      if(_zz_57)begin
        img_reg_array_55_27_imag <= _zz_121;
      end
      if(_zz_58)begin
        img_reg_array_56_27_imag <= _zz_121;
      end
      if(_zz_59)begin
        img_reg_array_57_27_imag <= _zz_121;
      end
      if(_zz_60)begin
        img_reg_array_58_27_imag <= _zz_121;
      end
      if(_zz_61)begin
        img_reg_array_59_27_imag <= _zz_121;
      end
      if(_zz_62)begin
        img_reg_array_60_27_imag <= _zz_121;
      end
      if(_zz_63)begin
        img_reg_array_61_27_imag <= _zz_121;
      end
      if(_zz_64)begin
        img_reg_array_62_27_imag <= _zz_121;
      end
      if(_zz_65)begin
        img_reg_array_63_27_imag <= _zz_121;
      end
      if(_zz_2)begin
        img_reg_array_0_28_real <= _zz_122;
      end
      if(_zz_3)begin
        img_reg_array_1_28_real <= _zz_122;
      end
      if(_zz_4)begin
        img_reg_array_2_28_real <= _zz_122;
      end
      if(_zz_5)begin
        img_reg_array_3_28_real <= _zz_122;
      end
      if(_zz_6)begin
        img_reg_array_4_28_real <= _zz_122;
      end
      if(_zz_7)begin
        img_reg_array_5_28_real <= _zz_122;
      end
      if(_zz_8)begin
        img_reg_array_6_28_real <= _zz_122;
      end
      if(_zz_9)begin
        img_reg_array_7_28_real <= _zz_122;
      end
      if(_zz_10)begin
        img_reg_array_8_28_real <= _zz_122;
      end
      if(_zz_11)begin
        img_reg_array_9_28_real <= _zz_122;
      end
      if(_zz_12)begin
        img_reg_array_10_28_real <= _zz_122;
      end
      if(_zz_13)begin
        img_reg_array_11_28_real <= _zz_122;
      end
      if(_zz_14)begin
        img_reg_array_12_28_real <= _zz_122;
      end
      if(_zz_15)begin
        img_reg_array_13_28_real <= _zz_122;
      end
      if(_zz_16)begin
        img_reg_array_14_28_real <= _zz_122;
      end
      if(_zz_17)begin
        img_reg_array_15_28_real <= _zz_122;
      end
      if(_zz_18)begin
        img_reg_array_16_28_real <= _zz_122;
      end
      if(_zz_19)begin
        img_reg_array_17_28_real <= _zz_122;
      end
      if(_zz_20)begin
        img_reg_array_18_28_real <= _zz_122;
      end
      if(_zz_21)begin
        img_reg_array_19_28_real <= _zz_122;
      end
      if(_zz_22)begin
        img_reg_array_20_28_real <= _zz_122;
      end
      if(_zz_23)begin
        img_reg_array_21_28_real <= _zz_122;
      end
      if(_zz_24)begin
        img_reg_array_22_28_real <= _zz_122;
      end
      if(_zz_25)begin
        img_reg_array_23_28_real <= _zz_122;
      end
      if(_zz_26)begin
        img_reg_array_24_28_real <= _zz_122;
      end
      if(_zz_27)begin
        img_reg_array_25_28_real <= _zz_122;
      end
      if(_zz_28)begin
        img_reg_array_26_28_real <= _zz_122;
      end
      if(_zz_29)begin
        img_reg_array_27_28_real <= _zz_122;
      end
      if(_zz_30)begin
        img_reg_array_28_28_real <= _zz_122;
      end
      if(_zz_31)begin
        img_reg_array_29_28_real <= _zz_122;
      end
      if(_zz_32)begin
        img_reg_array_30_28_real <= _zz_122;
      end
      if(_zz_33)begin
        img_reg_array_31_28_real <= _zz_122;
      end
      if(_zz_34)begin
        img_reg_array_32_28_real <= _zz_122;
      end
      if(_zz_35)begin
        img_reg_array_33_28_real <= _zz_122;
      end
      if(_zz_36)begin
        img_reg_array_34_28_real <= _zz_122;
      end
      if(_zz_37)begin
        img_reg_array_35_28_real <= _zz_122;
      end
      if(_zz_38)begin
        img_reg_array_36_28_real <= _zz_122;
      end
      if(_zz_39)begin
        img_reg_array_37_28_real <= _zz_122;
      end
      if(_zz_40)begin
        img_reg_array_38_28_real <= _zz_122;
      end
      if(_zz_41)begin
        img_reg_array_39_28_real <= _zz_122;
      end
      if(_zz_42)begin
        img_reg_array_40_28_real <= _zz_122;
      end
      if(_zz_43)begin
        img_reg_array_41_28_real <= _zz_122;
      end
      if(_zz_44)begin
        img_reg_array_42_28_real <= _zz_122;
      end
      if(_zz_45)begin
        img_reg_array_43_28_real <= _zz_122;
      end
      if(_zz_46)begin
        img_reg_array_44_28_real <= _zz_122;
      end
      if(_zz_47)begin
        img_reg_array_45_28_real <= _zz_122;
      end
      if(_zz_48)begin
        img_reg_array_46_28_real <= _zz_122;
      end
      if(_zz_49)begin
        img_reg_array_47_28_real <= _zz_122;
      end
      if(_zz_50)begin
        img_reg_array_48_28_real <= _zz_122;
      end
      if(_zz_51)begin
        img_reg_array_49_28_real <= _zz_122;
      end
      if(_zz_52)begin
        img_reg_array_50_28_real <= _zz_122;
      end
      if(_zz_53)begin
        img_reg_array_51_28_real <= _zz_122;
      end
      if(_zz_54)begin
        img_reg_array_52_28_real <= _zz_122;
      end
      if(_zz_55)begin
        img_reg_array_53_28_real <= _zz_122;
      end
      if(_zz_56)begin
        img_reg_array_54_28_real <= _zz_122;
      end
      if(_zz_57)begin
        img_reg_array_55_28_real <= _zz_122;
      end
      if(_zz_58)begin
        img_reg_array_56_28_real <= _zz_122;
      end
      if(_zz_59)begin
        img_reg_array_57_28_real <= _zz_122;
      end
      if(_zz_60)begin
        img_reg_array_58_28_real <= _zz_122;
      end
      if(_zz_61)begin
        img_reg_array_59_28_real <= _zz_122;
      end
      if(_zz_62)begin
        img_reg_array_60_28_real <= _zz_122;
      end
      if(_zz_63)begin
        img_reg_array_61_28_real <= _zz_122;
      end
      if(_zz_64)begin
        img_reg_array_62_28_real <= _zz_122;
      end
      if(_zz_65)begin
        img_reg_array_63_28_real <= _zz_122;
      end
      if(_zz_2)begin
        img_reg_array_0_28_imag <= _zz_123;
      end
      if(_zz_3)begin
        img_reg_array_1_28_imag <= _zz_123;
      end
      if(_zz_4)begin
        img_reg_array_2_28_imag <= _zz_123;
      end
      if(_zz_5)begin
        img_reg_array_3_28_imag <= _zz_123;
      end
      if(_zz_6)begin
        img_reg_array_4_28_imag <= _zz_123;
      end
      if(_zz_7)begin
        img_reg_array_5_28_imag <= _zz_123;
      end
      if(_zz_8)begin
        img_reg_array_6_28_imag <= _zz_123;
      end
      if(_zz_9)begin
        img_reg_array_7_28_imag <= _zz_123;
      end
      if(_zz_10)begin
        img_reg_array_8_28_imag <= _zz_123;
      end
      if(_zz_11)begin
        img_reg_array_9_28_imag <= _zz_123;
      end
      if(_zz_12)begin
        img_reg_array_10_28_imag <= _zz_123;
      end
      if(_zz_13)begin
        img_reg_array_11_28_imag <= _zz_123;
      end
      if(_zz_14)begin
        img_reg_array_12_28_imag <= _zz_123;
      end
      if(_zz_15)begin
        img_reg_array_13_28_imag <= _zz_123;
      end
      if(_zz_16)begin
        img_reg_array_14_28_imag <= _zz_123;
      end
      if(_zz_17)begin
        img_reg_array_15_28_imag <= _zz_123;
      end
      if(_zz_18)begin
        img_reg_array_16_28_imag <= _zz_123;
      end
      if(_zz_19)begin
        img_reg_array_17_28_imag <= _zz_123;
      end
      if(_zz_20)begin
        img_reg_array_18_28_imag <= _zz_123;
      end
      if(_zz_21)begin
        img_reg_array_19_28_imag <= _zz_123;
      end
      if(_zz_22)begin
        img_reg_array_20_28_imag <= _zz_123;
      end
      if(_zz_23)begin
        img_reg_array_21_28_imag <= _zz_123;
      end
      if(_zz_24)begin
        img_reg_array_22_28_imag <= _zz_123;
      end
      if(_zz_25)begin
        img_reg_array_23_28_imag <= _zz_123;
      end
      if(_zz_26)begin
        img_reg_array_24_28_imag <= _zz_123;
      end
      if(_zz_27)begin
        img_reg_array_25_28_imag <= _zz_123;
      end
      if(_zz_28)begin
        img_reg_array_26_28_imag <= _zz_123;
      end
      if(_zz_29)begin
        img_reg_array_27_28_imag <= _zz_123;
      end
      if(_zz_30)begin
        img_reg_array_28_28_imag <= _zz_123;
      end
      if(_zz_31)begin
        img_reg_array_29_28_imag <= _zz_123;
      end
      if(_zz_32)begin
        img_reg_array_30_28_imag <= _zz_123;
      end
      if(_zz_33)begin
        img_reg_array_31_28_imag <= _zz_123;
      end
      if(_zz_34)begin
        img_reg_array_32_28_imag <= _zz_123;
      end
      if(_zz_35)begin
        img_reg_array_33_28_imag <= _zz_123;
      end
      if(_zz_36)begin
        img_reg_array_34_28_imag <= _zz_123;
      end
      if(_zz_37)begin
        img_reg_array_35_28_imag <= _zz_123;
      end
      if(_zz_38)begin
        img_reg_array_36_28_imag <= _zz_123;
      end
      if(_zz_39)begin
        img_reg_array_37_28_imag <= _zz_123;
      end
      if(_zz_40)begin
        img_reg_array_38_28_imag <= _zz_123;
      end
      if(_zz_41)begin
        img_reg_array_39_28_imag <= _zz_123;
      end
      if(_zz_42)begin
        img_reg_array_40_28_imag <= _zz_123;
      end
      if(_zz_43)begin
        img_reg_array_41_28_imag <= _zz_123;
      end
      if(_zz_44)begin
        img_reg_array_42_28_imag <= _zz_123;
      end
      if(_zz_45)begin
        img_reg_array_43_28_imag <= _zz_123;
      end
      if(_zz_46)begin
        img_reg_array_44_28_imag <= _zz_123;
      end
      if(_zz_47)begin
        img_reg_array_45_28_imag <= _zz_123;
      end
      if(_zz_48)begin
        img_reg_array_46_28_imag <= _zz_123;
      end
      if(_zz_49)begin
        img_reg_array_47_28_imag <= _zz_123;
      end
      if(_zz_50)begin
        img_reg_array_48_28_imag <= _zz_123;
      end
      if(_zz_51)begin
        img_reg_array_49_28_imag <= _zz_123;
      end
      if(_zz_52)begin
        img_reg_array_50_28_imag <= _zz_123;
      end
      if(_zz_53)begin
        img_reg_array_51_28_imag <= _zz_123;
      end
      if(_zz_54)begin
        img_reg_array_52_28_imag <= _zz_123;
      end
      if(_zz_55)begin
        img_reg_array_53_28_imag <= _zz_123;
      end
      if(_zz_56)begin
        img_reg_array_54_28_imag <= _zz_123;
      end
      if(_zz_57)begin
        img_reg_array_55_28_imag <= _zz_123;
      end
      if(_zz_58)begin
        img_reg_array_56_28_imag <= _zz_123;
      end
      if(_zz_59)begin
        img_reg_array_57_28_imag <= _zz_123;
      end
      if(_zz_60)begin
        img_reg_array_58_28_imag <= _zz_123;
      end
      if(_zz_61)begin
        img_reg_array_59_28_imag <= _zz_123;
      end
      if(_zz_62)begin
        img_reg_array_60_28_imag <= _zz_123;
      end
      if(_zz_63)begin
        img_reg_array_61_28_imag <= _zz_123;
      end
      if(_zz_64)begin
        img_reg_array_62_28_imag <= _zz_123;
      end
      if(_zz_65)begin
        img_reg_array_63_28_imag <= _zz_123;
      end
      if(_zz_2)begin
        img_reg_array_0_29_real <= _zz_124;
      end
      if(_zz_3)begin
        img_reg_array_1_29_real <= _zz_124;
      end
      if(_zz_4)begin
        img_reg_array_2_29_real <= _zz_124;
      end
      if(_zz_5)begin
        img_reg_array_3_29_real <= _zz_124;
      end
      if(_zz_6)begin
        img_reg_array_4_29_real <= _zz_124;
      end
      if(_zz_7)begin
        img_reg_array_5_29_real <= _zz_124;
      end
      if(_zz_8)begin
        img_reg_array_6_29_real <= _zz_124;
      end
      if(_zz_9)begin
        img_reg_array_7_29_real <= _zz_124;
      end
      if(_zz_10)begin
        img_reg_array_8_29_real <= _zz_124;
      end
      if(_zz_11)begin
        img_reg_array_9_29_real <= _zz_124;
      end
      if(_zz_12)begin
        img_reg_array_10_29_real <= _zz_124;
      end
      if(_zz_13)begin
        img_reg_array_11_29_real <= _zz_124;
      end
      if(_zz_14)begin
        img_reg_array_12_29_real <= _zz_124;
      end
      if(_zz_15)begin
        img_reg_array_13_29_real <= _zz_124;
      end
      if(_zz_16)begin
        img_reg_array_14_29_real <= _zz_124;
      end
      if(_zz_17)begin
        img_reg_array_15_29_real <= _zz_124;
      end
      if(_zz_18)begin
        img_reg_array_16_29_real <= _zz_124;
      end
      if(_zz_19)begin
        img_reg_array_17_29_real <= _zz_124;
      end
      if(_zz_20)begin
        img_reg_array_18_29_real <= _zz_124;
      end
      if(_zz_21)begin
        img_reg_array_19_29_real <= _zz_124;
      end
      if(_zz_22)begin
        img_reg_array_20_29_real <= _zz_124;
      end
      if(_zz_23)begin
        img_reg_array_21_29_real <= _zz_124;
      end
      if(_zz_24)begin
        img_reg_array_22_29_real <= _zz_124;
      end
      if(_zz_25)begin
        img_reg_array_23_29_real <= _zz_124;
      end
      if(_zz_26)begin
        img_reg_array_24_29_real <= _zz_124;
      end
      if(_zz_27)begin
        img_reg_array_25_29_real <= _zz_124;
      end
      if(_zz_28)begin
        img_reg_array_26_29_real <= _zz_124;
      end
      if(_zz_29)begin
        img_reg_array_27_29_real <= _zz_124;
      end
      if(_zz_30)begin
        img_reg_array_28_29_real <= _zz_124;
      end
      if(_zz_31)begin
        img_reg_array_29_29_real <= _zz_124;
      end
      if(_zz_32)begin
        img_reg_array_30_29_real <= _zz_124;
      end
      if(_zz_33)begin
        img_reg_array_31_29_real <= _zz_124;
      end
      if(_zz_34)begin
        img_reg_array_32_29_real <= _zz_124;
      end
      if(_zz_35)begin
        img_reg_array_33_29_real <= _zz_124;
      end
      if(_zz_36)begin
        img_reg_array_34_29_real <= _zz_124;
      end
      if(_zz_37)begin
        img_reg_array_35_29_real <= _zz_124;
      end
      if(_zz_38)begin
        img_reg_array_36_29_real <= _zz_124;
      end
      if(_zz_39)begin
        img_reg_array_37_29_real <= _zz_124;
      end
      if(_zz_40)begin
        img_reg_array_38_29_real <= _zz_124;
      end
      if(_zz_41)begin
        img_reg_array_39_29_real <= _zz_124;
      end
      if(_zz_42)begin
        img_reg_array_40_29_real <= _zz_124;
      end
      if(_zz_43)begin
        img_reg_array_41_29_real <= _zz_124;
      end
      if(_zz_44)begin
        img_reg_array_42_29_real <= _zz_124;
      end
      if(_zz_45)begin
        img_reg_array_43_29_real <= _zz_124;
      end
      if(_zz_46)begin
        img_reg_array_44_29_real <= _zz_124;
      end
      if(_zz_47)begin
        img_reg_array_45_29_real <= _zz_124;
      end
      if(_zz_48)begin
        img_reg_array_46_29_real <= _zz_124;
      end
      if(_zz_49)begin
        img_reg_array_47_29_real <= _zz_124;
      end
      if(_zz_50)begin
        img_reg_array_48_29_real <= _zz_124;
      end
      if(_zz_51)begin
        img_reg_array_49_29_real <= _zz_124;
      end
      if(_zz_52)begin
        img_reg_array_50_29_real <= _zz_124;
      end
      if(_zz_53)begin
        img_reg_array_51_29_real <= _zz_124;
      end
      if(_zz_54)begin
        img_reg_array_52_29_real <= _zz_124;
      end
      if(_zz_55)begin
        img_reg_array_53_29_real <= _zz_124;
      end
      if(_zz_56)begin
        img_reg_array_54_29_real <= _zz_124;
      end
      if(_zz_57)begin
        img_reg_array_55_29_real <= _zz_124;
      end
      if(_zz_58)begin
        img_reg_array_56_29_real <= _zz_124;
      end
      if(_zz_59)begin
        img_reg_array_57_29_real <= _zz_124;
      end
      if(_zz_60)begin
        img_reg_array_58_29_real <= _zz_124;
      end
      if(_zz_61)begin
        img_reg_array_59_29_real <= _zz_124;
      end
      if(_zz_62)begin
        img_reg_array_60_29_real <= _zz_124;
      end
      if(_zz_63)begin
        img_reg_array_61_29_real <= _zz_124;
      end
      if(_zz_64)begin
        img_reg_array_62_29_real <= _zz_124;
      end
      if(_zz_65)begin
        img_reg_array_63_29_real <= _zz_124;
      end
      if(_zz_2)begin
        img_reg_array_0_29_imag <= _zz_125;
      end
      if(_zz_3)begin
        img_reg_array_1_29_imag <= _zz_125;
      end
      if(_zz_4)begin
        img_reg_array_2_29_imag <= _zz_125;
      end
      if(_zz_5)begin
        img_reg_array_3_29_imag <= _zz_125;
      end
      if(_zz_6)begin
        img_reg_array_4_29_imag <= _zz_125;
      end
      if(_zz_7)begin
        img_reg_array_5_29_imag <= _zz_125;
      end
      if(_zz_8)begin
        img_reg_array_6_29_imag <= _zz_125;
      end
      if(_zz_9)begin
        img_reg_array_7_29_imag <= _zz_125;
      end
      if(_zz_10)begin
        img_reg_array_8_29_imag <= _zz_125;
      end
      if(_zz_11)begin
        img_reg_array_9_29_imag <= _zz_125;
      end
      if(_zz_12)begin
        img_reg_array_10_29_imag <= _zz_125;
      end
      if(_zz_13)begin
        img_reg_array_11_29_imag <= _zz_125;
      end
      if(_zz_14)begin
        img_reg_array_12_29_imag <= _zz_125;
      end
      if(_zz_15)begin
        img_reg_array_13_29_imag <= _zz_125;
      end
      if(_zz_16)begin
        img_reg_array_14_29_imag <= _zz_125;
      end
      if(_zz_17)begin
        img_reg_array_15_29_imag <= _zz_125;
      end
      if(_zz_18)begin
        img_reg_array_16_29_imag <= _zz_125;
      end
      if(_zz_19)begin
        img_reg_array_17_29_imag <= _zz_125;
      end
      if(_zz_20)begin
        img_reg_array_18_29_imag <= _zz_125;
      end
      if(_zz_21)begin
        img_reg_array_19_29_imag <= _zz_125;
      end
      if(_zz_22)begin
        img_reg_array_20_29_imag <= _zz_125;
      end
      if(_zz_23)begin
        img_reg_array_21_29_imag <= _zz_125;
      end
      if(_zz_24)begin
        img_reg_array_22_29_imag <= _zz_125;
      end
      if(_zz_25)begin
        img_reg_array_23_29_imag <= _zz_125;
      end
      if(_zz_26)begin
        img_reg_array_24_29_imag <= _zz_125;
      end
      if(_zz_27)begin
        img_reg_array_25_29_imag <= _zz_125;
      end
      if(_zz_28)begin
        img_reg_array_26_29_imag <= _zz_125;
      end
      if(_zz_29)begin
        img_reg_array_27_29_imag <= _zz_125;
      end
      if(_zz_30)begin
        img_reg_array_28_29_imag <= _zz_125;
      end
      if(_zz_31)begin
        img_reg_array_29_29_imag <= _zz_125;
      end
      if(_zz_32)begin
        img_reg_array_30_29_imag <= _zz_125;
      end
      if(_zz_33)begin
        img_reg_array_31_29_imag <= _zz_125;
      end
      if(_zz_34)begin
        img_reg_array_32_29_imag <= _zz_125;
      end
      if(_zz_35)begin
        img_reg_array_33_29_imag <= _zz_125;
      end
      if(_zz_36)begin
        img_reg_array_34_29_imag <= _zz_125;
      end
      if(_zz_37)begin
        img_reg_array_35_29_imag <= _zz_125;
      end
      if(_zz_38)begin
        img_reg_array_36_29_imag <= _zz_125;
      end
      if(_zz_39)begin
        img_reg_array_37_29_imag <= _zz_125;
      end
      if(_zz_40)begin
        img_reg_array_38_29_imag <= _zz_125;
      end
      if(_zz_41)begin
        img_reg_array_39_29_imag <= _zz_125;
      end
      if(_zz_42)begin
        img_reg_array_40_29_imag <= _zz_125;
      end
      if(_zz_43)begin
        img_reg_array_41_29_imag <= _zz_125;
      end
      if(_zz_44)begin
        img_reg_array_42_29_imag <= _zz_125;
      end
      if(_zz_45)begin
        img_reg_array_43_29_imag <= _zz_125;
      end
      if(_zz_46)begin
        img_reg_array_44_29_imag <= _zz_125;
      end
      if(_zz_47)begin
        img_reg_array_45_29_imag <= _zz_125;
      end
      if(_zz_48)begin
        img_reg_array_46_29_imag <= _zz_125;
      end
      if(_zz_49)begin
        img_reg_array_47_29_imag <= _zz_125;
      end
      if(_zz_50)begin
        img_reg_array_48_29_imag <= _zz_125;
      end
      if(_zz_51)begin
        img_reg_array_49_29_imag <= _zz_125;
      end
      if(_zz_52)begin
        img_reg_array_50_29_imag <= _zz_125;
      end
      if(_zz_53)begin
        img_reg_array_51_29_imag <= _zz_125;
      end
      if(_zz_54)begin
        img_reg_array_52_29_imag <= _zz_125;
      end
      if(_zz_55)begin
        img_reg_array_53_29_imag <= _zz_125;
      end
      if(_zz_56)begin
        img_reg_array_54_29_imag <= _zz_125;
      end
      if(_zz_57)begin
        img_reg_array_55_29_imag <= _zz_125;
      end
      if(_zz_58)begin
        img_reg_array_56_29_imag <= _zz_125;
      end
      if(_zz_59)begin
        img_reg_array_57_29_imag <= _zz_125;
      end
      if(_zz_60)begin
        img_reg_array_58_29_imag <= _zz_125;
      end
      if(_zz_61)begin
        img_reg_array_59_29_imag <= _zz_125;
      end
      if(_zz_62)begin
        img_reg_array_60_29_imag <= _zz_125;
      end
      if(_zz_63)begin
        img_reg_array_61_29_imag <= _zz_125;
      end
      if(_zz_64)begin
        img_reg_array_62_29_imag <= _zz_125;
      end
      if(_zz_65)begin
        img_reg_array_63_29_imag <= _zz_125;
      end
      if(_zz_2)begin
        img_reg_array_0_30_real <= _zz_126;
      end
      if(_zz_3)begin
        img_reg_array_1_30_real <= _zz_126;
      end
      if(_zz_4)begin
        img_reg_array_2_30_real <= _zz_126;
      end
      if(_zz_5)begin
        img_reg_array_3_30_real <= _zz_126;
      end
      if(_zz_6)begin
        img_reg_array_4_30_real <= _zz_126;
      end
      if(_zz_7)begin
        img_reg_array_5_30_real <= _zz_126;
      end
      if(_zz_8)begin
        img_reg_array_6_30_real <= _zz_126;
      end
      if(_zz_9)begin
        img_reg_array_7_30_real <= _zz_126;
      end
      if(_zz_10)begin
        img_reg_array_8_30_real <= _zz_126;
      end
      if(_zz_11)begin
        img_reg_array_9_30_real <= _zz_126;
      end
      if(_zz_12)begin
        img_reg_array_10_30_real <= _zz_126;
      end
      if(_zz_13)begin
        img_reg_array_11_30_real <= _zz_126;
      end
      if(_zz_14)begin
        img_reg_array_12_30_real <= _zz_126;
      end
      if(_zz_15)begin
        img_reg_array_13_30_real <= _zz_126;
      end
      if(_zz_16)begin
        img_reg_array_14_30_real <= _zz_126;
      end
      if(_zz_17)begin
        img_reg_array_15_30_real <= _zz_126;
      end
      if(_zz_18)begin
        img_reg_array_16_30_real <= _zz_126;
      end
      if(_zz_19)begin
        img_reg_array_17_30_real <= _zz_126;
      end
      if(_zz_20)begin
        img_reg_array_18_30_real <= _zz_126;
      end
      if(_zz_21)begin
        img_reg_array_19_30_real <= _zz_126;
      end
      if(_zz_22)begin
        img_reg_array_20_30_real <= _zz_126;
      end
      if(_zz_23)begin
        img_reg_array_21_30_real <= _zz_126;
      end
      if(_zz_24)begin
        img_reg_array_22_30_real <= _zz_126;
      end
      if(_zz_25)begin
        img_reg_array_23_30_real <= _zz_126;
      end
      if(_zz_26)begin
        img_reg_array_24_30_real <= _zz_126;
      end
      if(_zz_27)begin
        img_reg_array_25_30_real <= _zz_126;
      end
      if(_zz_28)begin
        img_reg_array_26_30_real <= _zz_126;
      end
      if(_zz_29)begin
        img_reg_array_27_30_real <= _zz_126;
      end
      if(_zz_30)begin
        img_reg_array_28_30_real <= _zz_126;
      end
      if(_zz_31)begin
        img_reg_array_29_30_real <= _zz_126;
      end
      if(_zz_32)begin
        img_reg_array_30_30_real <= _zz_126;
      end
      if(_zz_33)begin
        img_reg_array_31_30_real <= _zz_126;
      end
      if(_zz_34)begin
        img_reg_array_32_30_real <= _zz_126;
      end
      if(_zz_35)begin
        img_reg_array_33_30_real <= _zz_126;
      end
      if(_zz_36)begin
        img_reg_array_34_30_real <= _zz_126;
      end
      if(_zz_37)begin
        img_reg_array_35_30_real <= _zz_126;
      end
      if(_zz_38)begin
        img_reg_array_36_30_real <= _zz_126;
      end
      if(_zz_39)begin
        img_reg_array_37_30_real <= _zz_126;
      end
      if(_zz_40)begin
        img_reg_array_38_30_real <= _zz_126;
      end
      if(_zz_41)begin
        img_reg_array_39_30_real <= _zz_126;
      end
      if(_zz_42)begin
        img_reg_array_40_30_real <= _zz_126;
      end
      if(_zz_43)begin
        img_reg_array_41_30_real <= _zz_126;
      end
      if(_zz_44)begin
        img_reg_array_42_30_real <= _zz_126;
      end
      if(_zz_45)begin
        img_reg_array_43_30_real <= _zz_126;
      end
      if(_zz_46)begin
        img_reg_array_44_30_real <= _zz_126;
      end
      if(_zz_47)begin
        img_reg_array_45_30_real <= _zz_126;
      end
      if(_zz_48)begin
        img_reg_array_46_30_real <= _zz_126;
      end
      if(_zz_49)begin
        img_reg_array_47_30_real <= _zz_126;
      end
      if(_zz_50)begin
        img_reg_array_48_30_real <= _zz_126;
      end
      if(_zz_51)begin
        img_reg_array_49_30_real <= _zz_126;
      end
      if(_zz_52)begin
        img_reg_array_50_30_real <= _zz_126;
      end
      if(_zz_53)begin
        img_reg_array_51_30_real <= _zz_126;
      end
      if(_zz_54)begin
        img_reg_array_52_30_real <= _zz_126;
      end
      if(_zz_55)begin
        img_reg_array_53_30_real <= _zz_126;
      end
      if(_zz_56)begin
        img_reg_array_54_30_real <= _zz_126;
      end
      if(_zz_57)begin
        img_reg_array_55_30_real <= _zz_126;
      end
      if(_zz_58)begin
        img_reg_array_56_30_real <= _zz_126;
      end
      if(_zz_59)begin
        img_reg_array_57_30_real <= _zz_126;
      end
      if(_zz_60)begin
        img_reg_array_58_30_real <= _zz_126;
      end
      if(_zz_61)begin
        img_reg_array_59_30_real <= _zz_126;
      end
      if(_zz_62)begin
        img_reg_array_60_30_real <= _zz_126;
      end
      if(_zz_63)begin
        img_reg_array_61_30_real <= _zz_126;
      end
      if(_zz_64)begin
        img_reg_array_62_30_real <= _zz_126;
      end
      if(_zz_65)begin
        img_reg_array_63_30_real <= _zz_126;
      end
      if(_zz_2)begin
        img_reg_array_0_30_imag <= _zz_127;
      end
      if(_zz_3)begin
        img_reg_array_1_30_imag <= _zz_127;
      end
      if(_zz_4)begin
        img_reg_array_2_30_imag <= _zz_127;
      end
      if(_zz_5)begin
        img_reg_array_3_30_imag <= _zz_127;
      end
      if(_zz_6)begin
        img_reg_array_4_30_imag <= _zz_127;
      end
      if(_zz_7)begin
        img_reg_array_5_30_imag <= _zz_127;
      end
      if(_zz_8)begin
        img_reg_array_6_30_imag <= _zz_127;
      end
      if(_zz_9)begin
        img_reg_array_7_30_imag <= _zz_127;
      end
      if(_zz_10)begin
        img_reg_array_8_30_imag <= _zz_127;
      end
      if(_zz_11)begin
        img_reg_array_9_30_imag <= _zz_127;
      end
      if(_zz_12)begin
        img_reg_array_10_30_imag <= _zz_127;
      end
      if(_zz_13)begin
        img_reg_array_11_30_imag <= _zz_127;
      end
      if(_zz_14)begin
        img_reg_array_12_30_imag <= _zz_127;
      end
      if(_zz_15)begin
        img_reg_array_13_30_imag <= _zz_127;
      end
      if(_zz_16)begin
        img_reg_array_14_30_imag <= _zz_127;
      end
      if(_zz_17)begin
        img_reg_array_15_30_imag <= _zz_127;
      end
      if(_zz_18)begin
        img_reg_array_16_30_imag <= _zz_127;
      end
      if(_zz_19)begin
        img_reg_array_17_30_imag <= _zz_127;
      end
      if(_zz_20)begin
        img_reg_array_18_30_imag <= _zz_127;
      end
      if(_zz_21)begin
        img_reg_array_19_30_imag <= _zz_127;
      end
      if(_zz_22)begin
        img_reg_array_20_30_imag <= _zz_127;
      end
      if(_zz_23)begin
        img_reg_array_21_30_imag <= _zz_127;
      end
      if(_zz_24)begin
        img_reg_array_22_30_imag <= _zz_127;
      end
      if(_zz_25)begin
        img_reg_array_23_30_imag <= _zz_127;
      end
      if(_zz_26)begin
        img_reg_array_24_30_imag <= _zz_127;
      end
      if(_zz_27)begin
        img_reg_array_25_30_imag <= _zz_127;
      end
      if(_zz_28)begin
        img_reg_array_26_30_imag <= _zz_127;
      end
      if(_zz_29)begin
        img_reg_array_27_30_imag <= _zz_127;
      end
      if(_zz_30)begin
        img_reg_array_28_30_imag <= _zz_127;
      end
      if(_zz_31)begin
        img_reg_array_29_30_imag <= _zz_127;
      end
      if(_zz_32)begin
        img_reg_array_30_30_imag <= _zz_127;
      end
      if(_zz_33)begin
        img_reg_array_31_30_imag <= _zz_127;
      end
      if(_zz_34)begin
        img_reg_array_32_30_imag <= _zz_127;
      end
      if(_zz_35)begin
        img_reg_array_33_30_imag <= _zz_127;
      end
      if(_zz_36)begin
        img_reg_array_34_30_imag <= _zz_127;
      end
      if(_zz_37)begin
        img_reg_array_35_30_imag <= _zz_127;
      end
      if(_zz_38)begin
        img_reg_array_36_30_imag <= _zz_127;
      end
      if(_zz_39)begin
        img_reg_array_37_30_imag <= _zz_127;
      end
      if(_zz_40)begin
        img_reg_array_38_30_imag <= _zz_127;
      end
      if(_zz_41)begin
        img_reg_array_39_30_imag <= _zz_127;
      end
      if(_zz_42)begin
        img_reg_array_40_30_imag <= _zz_127;
      end
      if(_zz_43)begin
        img_reg_array_41_30_imag <= _zz_127;
      end
      if(_zz_44)begin
        img_reg_array_42_30_imag <= _zz_127;
      end
      if(_zz_45)begin
        img_reg_array_43_30_imag <= _zz_127;
      end
      if(_zz_46)begin
        img_reg_array_44_30_imag <= _zz_127;
      end
      if(_zz_47)begin
        img_reg_array_45_30_imag <= _zz_127;
      end
      if(_zz_48)begin
        img_reg_array_46_30_imag <= _zz_127;
      end
      if(_zz_49)begin
        img_reg_array_47_30_imag <= _zz_127;
      end
      if(_zz_50)begin
        img_reg_array_48_30_imag <= _zz_127;
      end
      if(_zz_51)begin
        img_reg_array_49_30_imag <= _zz_127;
      end
      if(_zz_52)begin
        img_reg_array_50_30_imag <= _zz_127;
      end
      if(_zz_53)begin
        img_reg_array_51_30_imag <= _zz_127;
      end
      if(_zz_54)begin
        img_reg_array_52_30_imag <= _zz_127;
      end
      if(_zz_55)begin
        img_reg_array_53_30_imag <= _zz_127;
      end
      if(_zz_56)begin
        img_reg_array_54_30_imag <= _zz_127;
      end
      if(_zz_57)begin
        img_reg_array_55_30_imag <= _zz_127;
      end
      if(_zz_58)begin
        img_reg_array_56_30_imag <= _zz_127;
      end
      if(_zz_59)begin
        img_reg_array_57_30_imag <= _zz_127;
      end
      if(_zz_60)begin
        img_reg_array_58_30_imag <= _zz_127;
      end
      if(_zz_61)begin
        img_reg_array_59_30_imag <= _zz_127;
      end
      if(_zz_62)begin
        img_reg_array_60_30_imag <= _zz_127;
      end
      if(_zz_63)begin
        img_reg_array_61_30_imag <= _zz_127;
      end
      if(_zz_64)begin
        img_reg_array_62_30_imag <= _zz_127;
      end
      if(_zz_65)begin
        img_reg_array_63_30_imag <= _zz_127;
      end
      if(_zz_2)begin
        img_reg_array_0_31_real <= _zz_128;
      end
      if(_zz_3)begin
        img_reg_array_1_31_real <= _zz_128;
      end
      if(_zz_4)begin
        img_reg_array_2_31_real <= _zz_128;
      end
      if(_zz_5)begin
        img_reg_array_3_31_real <= _zz_128;
      end
      if(_zz_6)begin
        img_reg_array_4_31_real <= _zz_128;
      end
      if(_zz_7)begin
        img_reg_array_5_31_real <= _zz_128;
      end
      if(_zz_8)begin
        img_reg_array_6_31_real <= _zz_128;
      end
      if(_zz_9)begin
        img_reg_array_7_31_real <= _zz_128;
      end
      if(_zz_10)begin
        img_reg_array_8_31_real <= _zz_128;
      end
      if(_zz_11)begin
        img_reg_array_9_31_real <= _zz_128;
      end
      if(_zz_12)begin
        img_reg_array_10_31_real <= _zz_128;
      end
      if(_zz_13)begin
        img_reg_array_11_31_real <= _zz_128;
      end
      if(_zz_14)begin
        img_reg_array_12_31_real <= _zz_128;
      end
      if(_zz_15)begin
        img_reg_array_13_31_real <= _zz_128;
      end
      if(_zz_16)begin
        img_reg_array_14_31_real <= _zz_128;
      end
      if(_zz_17)begin
        img_reg_array_15_31_real <= _zz_128;
      end
      if(_zz_18)begin
        img_reg_array_16_31_real <= _zz_128;
      end
      if(_zz_19)begin
        img_reg_array_17_31_real <= _zz_128;
      end
      if(_zz_20)begin
        img_reg_array_18_31_real <= _zz_128;
      end
      if(_zz_21)begin
        img_reg_array_19_31_real <= _zz_128;
      end
      if(_zz_22)begin
        img_reg_array_20_31_real <= _zz_128;
      end
      if(_zz_23)begin
        img_reg_array_21_31_real <= _zz_128;
      end
      if(_zz_24)begin
        img_reg_array_22_31_real <= _zz_128;
      end
      if(_zz_25)begin
        img_reg_array_23_31_real <= _zz_128;
      end
      if(_zz_26)begin
        img_reg_array_24_31_real <= _zz_128;
      end
      if(_zz_27)begin
        img_reg_array_25_31_real <= _zz_128;
      end
      if(_zz_28)begin
        img_reg_array_26_31_real <= _zz_128;
      end
      if(_zz_29)begin
        img_reg_array_27_31_real <= _zz_128;
      end
      if(_zz_30)begin
        img_reg_array_28_31_real <= _zz_128;
      end
      if(_zz_31)begin
        img_reg_array_29_31_real <= _zz_128;
      end
      if(_zz_32)begin
        img_reg_array_30_31_real <= _zz_128;
      end
      if(_zz_33)begin
        img_reg_array_31_31_real <= _zz_128;
      end
      if(_zz_34)begin
        img_reg_array_32_31_real <= _zz_128;
      end
      if(_zz_35)begin
        img_reg_array_33_31_real <= _zz_128;
      end
      if(_zz_36)begin
        img_reg_array_34_31_real <= _zz_128;
      end
      if(_zz_37)begin
        img_reg_array_35_31_real <= _zz_128;
      end
      if(_zz_38)begin
        img_reg_array_36_31_real <= _zz_128;
      end
      if(_zz_39)begin
        img_reg_array_37_31_real <= _zz_128;
      end
      if(_zz_40)begin
        img_reg_array_38_31_real <= _zz_128;
      end
      if(_zz_41)begin
        img_reg_array_39_31_real <= _zz_128;
      end
      if(_zz_42)begin
        img_reg_array_40_31_real <= _zz_128;
      end
      if(_zz_43)begin
        img_reg_array_41_31_real <= _zz_128;
      end
      if(_zz_44)begin
        img_reg_array_42_31_real <= _zz_128;
      end
      if(_zz_45)begin
        img_reg_array_43_31_real <= _zz_128;
      end
      if(_zz_46)begin
        img_reg_array_44_31_real <= _zz_128;
      end
      if(_zz_47)begin
        img_reg_array_45_31_real <= _zz_128;
      end
      if(_zz_48)begin
        img_reg_array_46_31_real <= _zz_128;
      end
      if(_zz_49)begin
        img_reg_array_47_31_real <= _zz_128;
      end
      if(_zz_50)begin
        img_reg_array_48_31_real <= _zz_128;
      end
      if(_zz_51)begin
        img_reg_array_49_31_real <= _zz_128;
      end
      if(_zz_52)begin
        img_reg_array_50_31_real <= _zz_128;
      end
      if(_zz_53)begin
        img_reg_array_51_31_real <= _zz_128;
      end
      if(_zz_54)begin
        img_reg_array_52_31_real <= _zz_128;
      end
      if(_zz_55)begin
        img_reg_array_53_31_real <= _zz_128;
      end
      if(_zz_56)begin
        img_reg_array_54_31_real <= _zz_128;
      end
      if(_zz_57)begin
        img_reg_array_55_31_real <= _zz_128;
      end
      if(_zz_58)begin
        img_reg_array_56_31_real <= _zz_128;
      end
      if(_zz_59)begin
        img_reg_array_57_31_real <= _zz_128;
      end
      if(_zz_60)begin
        img_reg_array_58_31_real <= _zz_128;
      end
      if(_zz_61)begin
        img_reg_array_59_31_real <= _zz_128;
      end
      if(_zz_62)begin
        img_reg_array_60_31_real <= _zz_128;
      end
      if(_zz_63)begin
        img_reg_array_61_31_real <= _zz_128;
      end
      if(_zz_64)begin
        img_reg_array_62_31_real <= _zz_128;
      end
      if(_zz_65)begin
        img_reg_array_63_31_real <= _zz_128;
      end
      if(_zz_2)begin
        img_reg_array_0_31_imag <= _zz_129;
      end
      if(_zz_3)begin
        img_reg_array_1_31_imag <= _zz_129;
      end
      if(_zz_4)begin
        img_reg_array_2_31_imag <= _zz_129;
      end
      if(_zz_5)begin
        img_reg_array_3_31_imag <= _zz_129;
      end
      if(_zz_6)begin
        img_reg_array_4_31_imag <= _zz_129;
      end
      if(_zz_7)begin
        img_reg_array_5_31_imag <= _zz_129;
      end
      if(_zz_8)begin
        img_reg_array_6_31_imag <= _zz_129;
      end
      if(_zz_9)begin
        img_reg_array_7_31_imag <= _zz_129;
      end
      if(_zz_10)begin
        img_reg_array_8_31_imag <= _zz_129;
      end
      if(_zz_11)begin
        img_reg_array_9_31_imag <= _zz_129;
      end
      if(_zz_12)begin
        img_reg_array_10_31_imag <= _zz_129;
      end
      if(_zz_13)begin
        img_reg_array_11_31_imag <= _zz_129;
      end
      if(_zz_14)begin
        img_reg_array_12_31_imag <= _zz_129;
      end
      if(_zz_15)begin
        img_reg_array_13_31_imag <= _zz_129;
      end
      if(_zz_16)begin
        img_reg_array_14_31_imag <= _zz_129;
      end
      if(_zz_17)begin
        img_reg_array_15_31_imag <= _zz_129;
      end
      if(_zz_18)begin
        img_reg_array_16_31_imag <= _zz_129;
      end
      if(_zz_19)begin
        img_reg_array_17_31_imag <= _zz_129;
      end
      if(_zz_20)begin
        img_reg_array_18_31_imag <= _zz_129;
      end
      if(_zz_21)begin
        img_reg_array_19_31_imag <= _zz_129;
      end
      if(_zz_22)begin
        img_reg_array_20_31_imag <= _zz_129;
      end
      if(_zz_23)begin
        img_reg_array_21_31_imag <= _zz_129;
      end
      if(_zz_24)begin
        img_reg_array_22_31_imag <= _zz_129;
      end
      if(_zz_25)begin
        img_reg_array_23_31_imag <= _zz_129;
      end
      if(_zz_26)begin
        img_reg_array_24_31_imag <= _zz_129;
      end
      if(_zz_27)begin
        img_reg_array_25_31_imag <= _zz_129;
      end
      if(_zz_28)begin
        img_reg_array_26_31_imag <= _zz_129;
      end
      if(_zz_29)begin
        img_reg_array_27_31_imag <= _zz_129;
      end
      if(_zz_30)begin
        img_reg_array_28_31_imag <= _zz_129;
      end
      if(_zz_31)begin
        img_reg_array_29_31_imag <= _zz_129;
      end
      if(_zz_32)begin
        img_reg_array_30_31_imag <= _zz_129;
      end
      if(_zz_33)begin
        img_reg_array_31_31_imag <= _zz_129;
      end
      if(_zz_34)begin
        img_reg_array_32_31_imag <= _zz_129;
      end
      if(_zz_35)begin
        img_reg_array_33_31_imag <= _zz_129;
      end
      if(_zz_36)begin
        img_reg_array_34_31_imag <= _zz_129;
      end
      if(_zz_37)begin
        img_reg_array_35_31_imag <= _zz_129;
      end
      if(_zz_38)begin
        img_reg_array_36_31_imag <= _zz_129;
      end
      if(_zz_39)begin
        img_reg_array_37_31_imag <= _zz_129;
      end
      if(_zz_40)begin
        img_reg_array_38_31_imag <= _zz_129;
      end
      if(_zz_41)begin
        img_reg_array_39_31_imag <= _zz_129;
      end
      if(_zz_42)begin
        img_reg_array_40_31_imag <= _zz_129;
      end
      if(_zz_43)begin
        img_reg_array_41_31_imag <= _zz_129;
      end
      if(_zz_44)begin
        img_reg_array_42_31_imag <= _zz_129;
      end
      if(_zz_45)begin
        img_reg_array_43_31_imag <= _zz_129;
      end
      if(_zz_46)begin
        img_reg_array_44_31_imag <= _zz_129;
      end
      if(_zz_47)begin
        img_reg_array_45_31_imag <= _zz_129;
      end
      if(_zz_48)begin
        img_reg_array_46_31_imag <= _zz_129;
      end
      if(_zz_49)begin
        img_reg_array_47_31_imag <= _zz_129;
      end
      if(_zz_50)begin
        img_reg_array_48_31_imag <= _zz_129;
      end
      if(_zz_51)begin
        img_reg_array_49_31_imag <= _zz_129;
      end
      if(_zz_52)begin
        img_reg_array_50_31_imag <= _zz_129;
      end
      if(_zz_53)begin
        img_reg_array_51_31_imag <= _zz_129;
      end
      if(_zz_54)begin
        img_reg_array_52_31_imag <= _zz_129;
      end
      if(_zz_55)begin
        img_reg_array_53_31_imag <= _zz_129;
      end
      if(_zz_56)begin
        img_reg_array_54_31_imag <= _zz_129;
      end
      if(_zz_57)begin
        img_reg_array_55_31_imag <= _zz_129;
      end
      if(_zz_58)begin
        img_reg_array_56_31_imag <= _zz_129;
      end
      if(_zz_59)begin
        img_reg_array_57_31_imag <= _zz_129;
      end
      if(_zz_60)begin
        img_reg_array_58_31_imag <= _zz_129;
      end
      if(_zz_61)begin
        img_reg_array_59_31_imag <= _zz_129;
      end
      if(_zz_62)begin
        img_reg_array_60_31_imag <= _zz_129;
      end
      if(_zz_63)begin
        img_reg_array_61_31_imag <= _zz_129;
      end
      if(_zz_64)begin
        img_reg_array_62_31_imag <= _zz_129;
      end
      if(_zz_65)begin
        img_reg_array_63_31_imag <= _zz_129;
      end
      if(_zz_2)begin
        img_reg_array_0_32_real <= _zz_130;
      end
      if(_zz_3)begin
        img_reg_array_1_32_real <= _zz_130;
      end
      if(_zz_4)begin
        img_reg_array_2_32_real <= _zz_130;
      end
      if(_zz_5)begin
        img_reg_array_3_32_real <= _zz_130;
      end
      if(_zz_6)begin
        img_reg_array_4_32_real <= _zz_130;
      end
      if(_zz_7)begin
        img_reg_array_5_32_real <= _zz_130;
      end
      if(_zz_8)begin
        img_reg_array_6_32_real <= _zz_130;
      end
      if(_zz_9)begin
        img_reg_array_7_32_real <= _zz_130;
      end
      if(_zz_10)begin
        img_reg_array_8_32_real <= _zz_130;
      end
      if(_zz_11)begin
        img_reg_array_9_32_real <= _zz_130;
      end
      if(_zz_12)begin
        img_reg_array_10_32_real <= _zz_130;
      end
      if(_zz_13)begin
        img_reg_array_11_32_real <= _zz_130;
      end
      if(_zz_14)begin
        img_reg_array_12_32_real <= _zz_130;
      end
      if(_zz_15)begin
        img_reg_array_13_32_real <= _zz_130;
      end
      if(_zz_16)begin
        img_reg_array_14_32_real <= _zz_130;
      end
      if(_zz_17)begin
        img_reg_array_15_32_real <= _zz_130;
      end
      if(_zz_18)begin
        img_reg_array_16_32_real <= _zz_130;
      end
      if(_zz_19)begin
        img_reg_array_17_32_real <= _zz_130;
      end
      if(_zz_20)begin
        img_reg_array_18_32_real <= _zz_130;
      end
      if(_zz_21)begin
        img_reg_array_19_32_real <= _zz_130;
      end
      if(_zz_22)begin
        img_reg_array_20_32_real <= _zz_130;
      end
      if(_zz_23)begin
        img_reg_array_21_32_real <= _zz_130;
      end
      if(_zz_24)begin
        img_reg_array_22_32_real <= _zz_130;
      end
      if(_zz_25)begin
        img_reg_array_23_32_real <= _zz_130;
      end
      if(_zz_26)begin
        img_reg_array_24_32_real <= _zz_130;
      end
      if(_zz_27)begin
        img_reg_array_25_32_real <= _zz_130;
      end
      if(_zz_28)begin
        img_reg_array_26_32_real <= _zz_130;
      end
      if(_zz_29)begin
        img_reg_array_27_32_real <= _zz_130;
      end
      if(_zz_30)begin
        img_reg_array_28_32_real <= _zz_130;
      end
      if(_zz_31)begin
        img_reg_array_29_32_real <= _zz_130;
      end
      if(_zz_32)begin
        img_reg_array_30_32_real <= _zz_130;
      end
      if(_zz_33)begin
        img_reg_array_31_32_real <= _zz_130;
      end
      if(_zz_34)begin
        img_reg_array_32_32_real <= _zz_130;
      end
      if(_zz_35)begin
        img_reg_array_33_32_real <= _zz_130;
      end
      if(_zz_36)begin
        img_reg_array_34_32_real <= _zz_130;
      end
      if(_zz_37)begin
        img_reg_array_35_32_real <= _zz_130;
      end
      if(_zz_38)begin
        img_reg_array_36_32_real <= _zz_130;
      end
      if(_zz_39)begin
        img_reg_array_37_32_real <= _zz_130;
      end
      if(_zz_40)begin
        img_reg_array_38_32_real <= _zz_130;
      end
      if(_zz_41)begin
        img_reg_array_39_32_real <= _zz_130;
      end
      if(_zz_42)begin
        img_reg_array_40_32_real <= _zz_130;
      end
      if(_zz_43)begin
        img_reg_array_41_32_real <= _zz_130;
      end
      if(_zz_44)begin
        img_reg_array_42_32_real <= _zz_130;
      end
      if(_zz_45)begin
        img_reg_array_43_32_real <= _zz_130;
      end
      if(_zz_46)begin
        img_reg_array_44_32_real <= _zz_130;
      end
      if(_zz_47)begin
        img_reg_array_45_32_real <= _zz_130;
      end
      if(_zz_48)begin
        img_reg_array_46_32_real <= _zz_130;
      end
      if(_zz_49)begin
        img_reg_array_47_32_real <= _zz_130;
      end
      if(_zz_50)begin
        img_reg_array_48_32_real <= _zz_130;
      end
      if(_zz_51)begin
        img_reg_array_49_32_real <= _zz_130;
      end
      if(_zz_52)begin
        img_reg_array_50_32_real <= _zz_130;
      end
      if(_zz_53)begin
        img_reg_array_51_32_real <= _zz_130;
      end
      if(_zz_54)begin
        img_reg_array_52_32_real <= _zz_130;
      end
      if(_zz_55)begin
        img_reg_array_53_32_real <= _zz_130;
      end
      if(_zz_56)begin
        img_reg_array_54_32_real <= _zz_130;
      end
      if(_zz_57)begin
        img_reg_array_55_32_real <= _zz_130;
      end
      if(_zz_58)begin
        img_reg_array_56_32_real <= _zz_130;
      end
      if(_zz_59)begin
        img_reg_array_57_32_real <= _zz_130;
      end
      if(_zz_60)begin
        img_reg_array_58_32_real <= _zz_130;
      end
      if(_zz_61)begin
        img_reg_array_59_32_real <= _zz_130;
      end
      if(_zz_62)begin
        img_reg_array_60_32_real <= _zz_130;
      end
      if(_zz_63)begin
        img_reg_array_61_32_real <= _zz_130;
      end
      if(_zz_64)begin
        img_reg_array_62_32_real <= _zz_130;
      end
      if(_zz_65)begin
        img_reg_array_63_32_real <= _zz_130;
      end
      if(_zz_2)begin
        img_reg_array_0_32_imag <= _zz_131;
      end
      if(_zz_3)begin
        img_reg_array_1_32_imag <= _zz_131;
      end
      if(_zz_4)begin
        img_reg_array_2_32_imag <= _zz_131;
      end
      if(_zz_5)begin
        img_reg_array_3_32_imag <= _zz_131;
      end
      if(_zz_6)begin
        img_reg_array_4_32_imag <= _zz_131;
      end
      if(_zz_7)begin
        img_reg_array_5_32_imag <= _zz_131;
      end
      if(_zz_8)begin
        img_reg_array_6_32_imag <= _zz_131;
      end
      if(_zz_9)begin
        img_reg_array_7_32_imag <= _zz_131;
      end
      if(_zz_10)begin
        img_reg_array_8_32_imag <= _zz_131;
      end
      if(_zz_11)begin
        img_reg_array_9_32_imag <= _zz_131;
      end
      if(_zz_12)begin
        img_reg_array_10_32_imag <= _zz_131;
      end
      if(_zz_13)begin
        img_reg_array_11_32_imag <= _zz_131;
      end
      if(_zz_14)begin
        img_reg_array_12_32_imag <= _zz_131;
      end
      if(_zz_15)begin
        img_reg_array_13_32_imag <= _zz_131;
      end
      if(_zz_16)begin
        img_reg_array_14_32_imag <= _zz_131;
      end
      if(_zz_17)begin
        img_reg_array_15_32_imag <= _zz_131;
      end
      if(_zz_18)begin
        img_reg_array_16_32_imag <= _zz_131;
      end
      if(_zz_19)begin
        img_reg_array_17_32_imag <= _zz_131;
      end
      if(_zz_20)begin
        img_reg_array_18_32_imag <= _zz_131;
      end
      if(_zz_21)begin
        img_reg_array_19_32_imag <= _zz_131;
      end
      if(_zz_22)begin
        img_reg_array_20_32_imag <= _zz_131;
      end
      if(_zz_23)begin
        img_reg_array_21_32_imag <= _zz_131;
      end
      if(_zz_24)begin
        img_reg_array_22_32_imag <= _zz_131;
      end
      if(_zz_25)begin
        img_reg_array_23_32_imag <= _zz_131;
      end
      if(_zz_26)begin
        img_reg_array_24_32_imag <= _zz_131;
      end
      if(_zz_27)begin
        img_reg_array_25_32_imag <= _zz_131;
      end
      if(_zz_28)begin
        img_reg_array_26_32_imag <= _zz_131;
      end
      if(_zz_29)begin
        img_reg_array_27_32_imag <= _zz_131;
      end
      if(_zz_30)begin
        img_reg_array_28_32_imag <= _zz_131;
      end
      if(_zz_31)begin
        img_reg_array_29_32_imag <= _zz_131;
      end
      if(_zz_32)begin
        img_reg_array_30_32_imag <= _zz_131;
      end
      if(_zz_33)begin
        img_reg_array_31_32_imag <= _zz_131;
      end
      if(_zz_34)begin
        img_reg_array_32_32_imag <= _zz_131;
      end
      if(_zz_35)begin
        img_reg_array_33_32_imag <= _zz_131;
      end
      if(_zz_36)begin
        img_reg_array_34_32_imag <= _zz_131;
      end
      if(_zz_37)begin
        img_reg_array_35_32_imag <= _zz_131;
      end
      if(_zz_38)begin
        img_reg_array_36_32_imag <= _zz_131;
      end
      if(_zz_39)begin
        img_reg_array_37_32_imag <= _zz_131;
      end
      if(_zz_40)begin
        img_reg_array_38_32_imag <= _zz_131;
      end
      if(_zz_41)begin
        img_reg_array_39_32_imag <= _zz_131;
      end
      if(_zz_42)begin
        img_reg_array_40_32_imag <= _zz_131;
      end
      if(_zz_43)begin
        img_reg_array_41_32_imag <= _zz_131;
      end
      if(_zz_44)begin
        img_reg_array_42_32_imag <= _zz_131;
      end
      if(_zz_45)begin
        img_reg_array_43_32_imag <= _zz_131;
      end
      if(_zz_46)begin
        img_reg_array_44_32_imag <= _zz_131;
      end
      if(_zz_47)begin
        img_reg_array_45_32_imag <= _zz_131;
      end
      if(_zz_48)begin
        img_reg_array_46_32_imag <= _zz_131;
      end
      if(_zz_49)begin
        img_reg_array_47_32_imag <= _zz_131;
      end
      if(_zz_50)begin
        img_reg_array_48_32_imag <= _zz_131;
      end
      if(_zz_51)begin
        img_reg_array_49_32_imag <= _zz_131;
      end
      if(_zz_52)begin
        img_reg_array_50_32_imag <= _zz_131;
      end
      if(_zz_53)begin
        img_reg_array_51_32_imag <= _zz_131;
      end
      if(_zz_54)begin
        img_reg_array_52_32_imag <= _zz_131;
      end
      if(_zz_55)begin
        img_reg_array_53_32_imag <= _zz_131;
      end
      if(_zz_56)begin
        img_reg_array_54_32_imag <= _zz_131;
      end
      if(_zz_57)begin
        img_reg_array_55_32_imag <= _zz_131;
      end
      if(_zz_58)begin
        img_reg_array_56_32_imag <= _zz_131;
      end
      if(_zz_59)begin
        img_reg_array_57_32_imag <= _zz_131;
      end
      if(_zz_60)begin
        img_reg_array_58_32_imag <= _zz_131;
      end
      if(_zz_61)begin
        img_reg_array_59_32_imag <= _zz_131;
      end
      if(_zz_62)begin
        img_reg_array_60_32_imag <= _zz_131;
      end
      if(_zz_63)begin
        img_reg_array_61_32_imag <= _zz_131;
      end
      if(_zz_64)begin
        img_reg_array_62_32_imag <= _zz_131;
      end
      if(_zz_65)begin
        img_reg_array_63_32_imag <= _zz_131;
      end
      if(_zz_2)begin
        img_reg_array_0_33_real <= _zz_132;
      end
      if(_zz_3)begin
        img_reg_array_1_33_real <= _zz_132;
      end
      if(_zz_4)begin
        img_reg_array_2_33_real <= _zz_132;
      end
      if(_zz_5)begin
        img_reg_array_3_33_real <= _zz_132;
      end
      if(_zz_6)begin
        img_reg_array_4_33_real <= _zz_132;
      end
      if(_zz_7)begin
        img_reg_array_5_33_real <= _zz_132;
      end
      if(_zz_8)begin
        img_reg_array_6_33_real <= _zz_132;
      end
      if(_zz_9)begin
        img_reg_array_7_33_real <= _zz_132;
      end
      if(_zz_10)begin
        img_reg_array_8_33_real <= _zz_132;
      end
      if(_zz_11)begin
        img_reg_array_9_33_real <= _zz_132;
      end
      if(_zz_12)begin
        img_reg_array_10_33_real <= _zz_132;
      end
      if(_zz_13)begin
        img_reg_array_11_33_real <= _zz_132;
      end
      if(_zz_14)begin
        img_reg_array_12_33_real <= _zz_132;
      end
      if(_zz_15)begin
        img_reg_array_13_33_real <= _zz_132;
      end
      if(_zz_16)begin
        img_reg_array_14_33_real <= _zz_132;
      end
      if(_zz_17)begin
        img_reg_array_15_33_real <= _zz_132;
      end
      if(_zz_18)begin
        img_reg_array_16_33_real <= _zz_132;
      end
      if(_zz_19)begin
        img_reg_array_17_33_real <= _zz_132;
      end
      if(_zz_20)begin
        img_reg_array_18_33_real <= _zz_132;
      end
      if(_zz_21)begin
        img_reg_array_19_33_real <= _zz_132;
      end
      if(_zz_22)begin
        img_reg_array_20_33_real <= _zz_132;
      end
      if(_zz_23)begin
        img_reg_array_21_33_real <= _zz_132;
      end
      if(_zz_24)begin
        img_reg_array_22_33_real <= _zz_132;
      end
      if(_zz_25)begin
        img_reg_array_23_33_real <= _zz_132;
      end
      if(_zz_26)begin
        img_reg_array_24_33_real <= _zz_132;
      end
      if(_zz_27)begin
        img_reg_array_25_33_real <= _zz_132;
      end
      if(_zz_28)begin
        img_reg_array_26_33_real <= _zz_132;
      end
      if(_zz_29)begin
        img_reg_array_27_33_real <= _zz_132;
      end
      if(_zz_30)begin
        img_reg_array_28_33_real <= _zz_132;
      end
      if(_zz_31)begin
        img_reg_array_29_33_real <= _zz_132;
      end
      if(_zz_32)begin
        img_reg_array_30_33_real <= _zz_132;
      end
      if(_zz_33)begin
        img_reg_array_31_33_real <= _zz_132;
      end
      if(_zz_34)begin
        img_reg_array_32_33_real <= _zz_132;
      end
      if(_zz_35)begin
        img_reg_array_33_33_real <= _zz_132;
      end
      if(_zz_36)begin
        img_reg_array_34_33_real <= _zz_132;
      end
      if(_zz_37)begin
        img_reg_array_35_33_real <= _zz_132;
      end
      if(_zz_38)begin
        img_reg_array_36_33_real <= _zz_132;
      end
      if(_zz_39)begin
        img_reg_array_37_33_real <= _zz_132;
      end
      if(_zz_40)begin
        img_reg_array_38_33_real <= _zz_132;
      end
      if(_zz_41)begin
        img_reg_array_39_33_real <= _zz_132;
      end
      if(_zz_42)begin
        img_reg_array_40_33_real <= _zz_132;
      end
      if(_zz_43)begin
        img_reg_array_41_33_real <= _zz_132;
      end
      if(_zz_44)begin
        img_reg_array_42_33_real <= _zz_132;
      end
      if(_zz_45)begin
        img_reg_array_43_33_real <= _zz_132;
      end
      if(_zz_46)begin
        img_reg_array_44_33_real <= _zz_132;
      end
      if(_zz_47)begin
        img_reg_array_45_33_real <= _zz_132;
      end
      if(_zz_48)begin
        img_reg_array_46_33_real <= _zz_132;
      end
      if(_zz_49)begin
        img_reg_array_47_33_real <= _zz_132;
      end
      if(_zz_50)begin
        img_reg_array_48_33_real <= _zz_132;
      end
      if(_zz_51)begin
        img_reg_array_49_33_real <= _zz_132;
      end
      if(_zz_52)begin
        img_reg_array_50_33_real <= _zz_132;
      end
      if(_zz_53)begin
        img_reg_array_51_33_real <= _zz_132;
      end
      if(_zz_54)begin
        img_reg_array_52_33_real <= _zz_132;
      end
      if(_zz_55)begin
        img_reg_array_53_33_real <= _zz_132;
      end
      if(_zz_56)begin
        img_reg_array_54_33_real <= _zz_132;
      end
      if(_zz_57)begin
        img_reg_array_55_33_real <= _zz_132;
      end
      if(_zz_58)begin
        img_reg_array_56_33_real <= _zz_132;
      end
      if(_zz_59)begin
        img_reg_array_57_33_real <= _zz_132;
      end
      if(_zz_60)begin
        img_reg_array_58_33_real <= _zz_132;
      end
      if(_zz_61)begin
        img_reg_array_59_33_real <= _zz_132;
      end
      if(_zz_62)begin
        img_reg_array_60_33_real <= _zz_132;
      end
      if(_zz_63)begin
        img_reg_array_61_33_real <= _zz_132;
      end
      if(_zz_64)begin
        img_reg_array_62_33_real <= _zz_132;
      end
      if(_zz_65)begin
        img_reg_array_63_33_real <= _zz_132;
      end
      if(_zz_2)begin
        img_reg_array_0_33_imag <= _zz_133;
      end
      if(_zz_3)begin
        img_reg_array_1_33_imag <= _zz_133;
      end
      if(_zz_4)begin
        img_reg_array_2_33_imag <= _zz_133;
      end
      if(_zz_5)begin
        img_reg_array_3_33_imag <= _zz_133;
      end
      if(_zz_6)begin
        img_reg_array_4_33_imag <= _zz_133;
      end
      if(_zz_7)begin
        img_reg_array_5_33_imag <= _zz_133;
      end
      if(_zz_8)begin
        img_reg_array_6_33_imag <= _zz_133;
      end
      if(_zz_9)begin
        img_reg_array_7_33_imag <= _zz_133;
      end
      if(_zz_10)begin
        img_reg_array_8_33_imag <= _zz_133;
      end
      if(_zz_11)begin
        img_reg_array_9_33_imag <= _zz_133;
      end
      if(_zz_12)begin
        img_reg_array_10_33_imag <= _zz_133;
      end
      if(_zz_13)begin
        img_reg_array_11_33_imag <= _zz_133;
      end
      if(_zz_14)begin
        img_reg_array_12_33_imag <= _zz_133;
      end
      if(_zz_15)begin
        img_reg_array_13_33_imag <= _zz_133;
      end
      if(_zz_16)begin
        img_reg_array_14_33_imag <= _zz_133;
      end
      if(_zz_17)begin
        img_reg_array_15_33_imag <= _zz_133;
      end
      if(_zz_18)begin
        img_reg_array_16_33_imag <= _zz_133;
      end
      if(_zz_19)begin
        img_reg_array_17_33_imag <= _zz_133;
      end
      if(_zz_20)begin
        img_reg_array_18_33_imag <= _zz_133;
      end
      if(_zz_21)begin
        img_reg_array_19_33_imag <= _zz_133;
      end
      if(_zz_22)begin
        img_reg_array_20_33_imag <= _zz_133;
      end
      if(_zz_23)begin
        img_reg_array_21_33_imag <= _zz_133;
      end
      if(_zz_24)begin
        img_reg_array_22_33_imag <= _zz_133;
      end
      if(_zz_25)begin
        img_reg_array_23_33_imag <= _zz_133;
      end
      if(_zz_26)begin
        img_reg_array_24_33_imag <= _zz_133;
      end
      if(_zz_27)begin
        img_reg_array_25_33_imag <= _zz_133;
      end
      if(_zz_28)begin
        img_reg_array_26_33_imag <= _zz_133;
      end
      if(_zz_29)begin
        img_reg_array_27_33_imag <= _zz_133;
      end
      if(_zz_30)begin
        img_reg_array_28_33_imag <= _zz_133;
      end
      if(_zz_31)begin
        img_reg_array_29_33_imag <= _zz_133;
      end
      if(_zz_32)begin
        img_reg_array_30_33_imag <= _zz_133;
      end
      if(_zz_33)begin
        img_reg_array_31_33_imag <= _zz_133;
      end
      if(_zz_34)begin
        img_reg_array_32_33_imag <= _zz_133;
      end
      if(_zz_35)begin
        img_reg_array_33_33_imag <= _zz_133;
      end
      if(_zz_36)begin
        img_reg_array_34_33_imag <= _zz_133;
      end
      if(_zz_37)begin
        img_reg_array_35_33_imag <= _zz_133;
      end
      if(_zz_38)begin
        img_reg_array_36_33_imag <= _zz_133;
      end
      if(_zz_39)begin
        img_reg_array_37_33_imag <= _zz_133;
      end
      if(_zz_40)begin
        img_reg_array_38_33_imag <= _zz_133;
      end
      if(_zz_41)begin
        img_reg_array_39_33_imag <= _zz_133;
      end
      if(_zz_42)begin
        img_reg_array_40_33_imag <= _zz_133;
      end
      if(_zz_43)begin
        img_reg_array_41_33_imag <= _zz_133;
      end
      if(_zz_44)begin
        img_reg_array_42_33_imag <= _zz_133;
      end
      if(_zz_45)begin
        img_reg_array_43_33_imag <= _zz_133;
      end
      if(_zz_46)begin
        img_reg_array_44_33_imag <= _zz_133;
      end
      if(_zz_47)begin
        img_reg_array_45_33_imag <= _zz_133;
      end
      if(_zz_48)begin
        img_reg_array_46_33_imag <= _zz_133;
      end
      if(_zz_49)begin
        img_reg_array_47_33_imag <= _zz_133;
      end
      if(_zz_50)begin
        img_reg_array_48_33_imag <= _zz_133;
      end
      if(_zz_51)begin
        img_reg_array_49_33_imag <= _zz_133;
      end
      if(_zz_52)begin
        img_reg_array_50_33_imag <= _zz_133;
      end
      if(_zz_53)begin
        img_reg_array_51_33_imag <= _zz_133;
      end
      if(_zz_54)begin
        img_reg_array_52_33_imag <= _zz_133;
      end
      if(_zz_55)begin
        img_reg_array_53_33_imag <= _zz_133;
      end
      if(_zz_56)begin
        img_reg_array_54_33_imag <= _zz_133;
      end
      if(_zz_57)begin
        img_reg_array_55_33_imag <= _zz_133;
      end
      if(_zz_58)begin
        img_reg_array_56_33_imag <= _zz_133;
      end
      if(_zz_59)begin
        img_reg_array_57_33_imag <= _zz_133;
      end
      if(_zz_60)begin
        img_reg_array_58_33_imag <= _zz_133;
      end
      if(_zz_61)begin
        img_reg_array_59_33_imag <= _zz_133;
      end
      if(_zz_62)begin
        img_reg_array_60_33_imag <= _zz_133;
      end
      if(_zz_63)begin
        img_reg_array_61_33_imag <= _zz_133;
      end
      if(_zz_64)begin
        img_reg_array_62_33_imag <= _zz_133;
      end
      if(_zz_65)begin
        img_reg_array_63_33_imag <= _zz_133;
      end
      if(_zz_2)begin
        img_reg_array_0_34_real <= _zz_134;
      end
      if(_zz_3)begin
        img_reg_array_1_34_real <= _zz_134;
      end
      if(_zz_4)begin
        img_reg_array_2_34_real <= _zz_134;
      end
      if(_zz_5)begin
        img_reg_array_3_34_real <= _zz_134;
      end
      if(_zz_6)begin
        img_reg_array_4_34_real <= _zz_134;
      end
      if(_zz_7)begin
        img_reg_array_5_34_real <= _zz_134;
      end
      if(_zz_8)begin
        img_reg_array_6_34_real <= _zz_134;
      end
      if(_zz_9)begin
        img_reg_array_7_34_real <= _zz_134;
      end
      if(_zz_10)begin
        img_reg_array_8_34_real <= _zz_134;
      end
      if(_zz_11)begin
        img_reg_array_9_34_real <= _zz_134;
      end
      if(_zz_12)begin
        img_reg_array_10_34_real <= _zz_134;
      end
      if(_zz_13)begin
        img_reg_array_11_34_real <= _zz_134;
      end
      if(_zz_14)begin
        img_reg_array_12_34_real <= _zz_134;
      end
      if(_zz_15)begin
        img_reg_array_13_34_real <= _zz_134;
      end
      if(_zz_16)begin
        img_reg_array_14_34_real <= _zz_134;
      end
      if(_zz_17)begin
        img_reg_array_15_34_real <= _zz_134;
      end
      if(_zz_18)begin
        img_reg_array_16_34_real <= _zz_134;
      end
      if(_zz_19)begin
        img_reg_array_17_34_real <= _zz_134;
      end
      if(_zz_20)begin
        img_reg_array_18_34_real <= _zz_134;
      end
      if(_zz_21)begin
        img_reg_array_19_34_real <= _zz_134;
      end
      if(_zz_22)begin
        img_reg_array_20_34_real <= _zz_134;
      end
      if(_zz_23)begin
        img_reg_array_21_34_real <= _zz_134;
      end
      if(_zz_24)begin
        img_reg_array_22_34_real <= _zz_134;
      end
      if(_zz_25)begin
        img_reg_array_23_34_real <= _zz_134;
      end
      if(_zz_26)begin
        img_reg_array_24_34_real <= _zz_134;
      end
      if(_zz_27)begin
        img_reg_array_25_34_real <= _zz_134;
      end
      if(_zz_28)begin
        img_reg_array_26_34_real <= _zz_134;
      end
      if(_zz_29)begin
        img_reg_array_27_34_real <= _zz_134;
      end
      if(_zz_30)begin
        img_reg_array_28_34_real <= _zz_134;
      end
      if(_zz_31)begin
        img_reg_array_29_34_real <= _zz_134;
      end
      if(_zz_32)begin
        img_reg_array_30_34_real <= _zz_134;
      end
      if(_zz_33)begin
        img_reg_array_31_34_real <= _zz_134;
      end
      if(_zz_34)begin
        img_reg_array_32_34_real <= _zz_134;
      end
      if(_zz_35)begin
        img_reg_array_33_34_real <= _zz_134;
      end
      if(_zz_36)begin
        img_reg_array_34_34_real <= _zz_134;
      end
      if(_zz_37)begin
        img_reg_array_35_34_real <= _zz_134;
      end
      if(_zz_38)begin
        img_reg_array_36_34_real <= _zz_134;
      end
      if(_zz_39)begin
        img_reg_array_37_34_real <= _zz_134;
      end
      if(_zz_40)begin
        img_reg_array_38_34_real <= _zz_134;
      end
      if(_zz_41)begin
        img_reg_array_39_34_real <= _zz_134;
      end
      if(_zz_42)begin
        img_reg_array_40_34_real <= _zz_134;
      end
      if(_zz_43)begin
        img_reg_array_41_34_real <= _zz_134;
      end
      if(_zz_44)begin
        img_reg_array_42_34_real <= _zz_134;
      end
      if(_zz_45)begin
        img_reg_array_43_34_real <= _zz_134;
      end
      if(_zz_46)begin
        img_reg_array_44_34_real <= _zz_134;
      end
      if(_zz_47)begin
        img_reg_array_45_34_real <= _zz_134;
      end
      if(_zz_48)begin
        img_reg_array_46_34_real <= _zz_134;
      end
      if(_zz_49)begin
        img_reg_array_47_34_real <= _zz_134;
      end
      if(_zz_50)begin
        img_reg_array_48_34_real <= _zz_134;
      end
      if(_zz_51)begin
        img_reg_array_49_34_real <= _zz_134;
      end
      if(_zz_52)begin
        img_reg_array_50_34_real <= _zz_134;
      end
      if(_zz_53)begin
        img_reg_array_51_34_real <= _zz_134;
      end
      if(_zz_54)begin
        img_reg_array_52_34_real <= _zz_134;
      end
      if(_zz_55)begin
        img_reg_array_53_34_real <= _zz_134;
      end
      if(_zz_56)begin
        img_reg_array_54_34_real <= _zz_134;
      end
      if(_zz_57)begin
        img_reg_array_55_34_real <= _zz_134;
      end
      if(_zz_58)begin
        img_reg_array_56_34_real <= _zz_134;
      end
      if(_zz_59)begin
        img_reg_array_57_34_real <= _zz_134;
      end
      if(_zz_60)begin
        img_reg_array_58_34_real <= _zz_134;
      end
      if(_zz_61)begin
        img_reg_array_59_34_real <= _zz_134;
      end
      if(_zz_62)begin
        img_reg_array_60_34_real <= _zz_134;
      end
      if(_zz_63)begin
        img_reg_array_61_34_real <= _zz_134;
      end
      if(_zz_64)begin
        img_reg_array_62_34_real <= _zz_134;
      end
      if(_zz_65)begin
        img_reg_array_63_34_real <= _zz_134;
      end
      if(_zz_2)begin
        img_reg_array_0_34_imag <= _zz_135;
      end
      if(_zz_3)begin
        img_reg_array_1_34_imag <= _zz_135;
      end
      if(_zz_4)begin
        img_reg_array_2_34_imag <= _zz_135;
      end
      if(_zz_5)begin
        img_reg_array_3_34_imag <= _zz_135;
      end
      if(_zz_6)begin
        img_reg_array_4_34_imag <= _zz_135;
      end
      if(_zz_7)begin
        img_reg_array_5_34_imag <= _zz_135;
      end
      if(_zz_8)begin
        img_reg_array_6_34_imag <= _zz_135;
      end
      if(_zz_9)begin
        img_reg_array_7_34_imag <= _zz_135;
      end
      if(_zz_10)begin
        img_reg_array_8_34_imag <= _zz_135;
      end
      if(_zz_11)begin
        img_reg_array_9_34_imag <= _zz_135;
      end
      if(_zz_12)begin
        img_reg_array_10_34_imag <= _zz_135;
      end
      if(_zz_13)begin
        img_reg_array_11_34_imag <= _zz_135;
      end
      if(_zz_14)begin
        img_reg_array_12_34_imag <= _zz_135;
      end
      if(_zz_15)begin
        img_reg_array_13_34_imag <= _zz_135;
      end
      if(_zz_16)begin
        img_reg_array_14_34_imag <= _zz_135;
      end
      if(_zz_17)begin
        img_reg_array_15_34_imag <= _zz_135;
      end
      if(_zz_18)begin
        img_reg_array_16_34_imag <= _zz_135;
      end
      if(_zz_19)begin
        img_reg_array_17_34_imag <= _zz_135;
      end
      if(_zz_20)begin
        img_reg_array_18_34_imag <= _zz_135;
      end
      if(_zz_21)begin
        img_reg_array_19_34_imag <= _zz_135;
      end
      if(_zz_22)begin
        img_reg_array_20_34_imag <= _zz_135;
      end
      if(_zz_23)begin
        img_reg_array_21_34_imag <= _zz_135;
      end
      if(_zz_24)begin
        img_reg_array_22_34_imag <= _zz_135;
      end
      if(_zz_25)begin
        img_reg_array_23_34_imag <= _zz_135;
      end
      if(_zz_26)begin
        img_reg_array_24_34_imag <= _zz_135;
      end
      if(_zz_27)begin
        img_reg_array_25_34_imag <= _zz_135;
      end
      if(_zz_28)begin
        img_reg_array_26_34_imag <= _zz_135;
      end
      if(_zz_29)begin
        img_reg_array_27_34_imag <= _zz_135;
      end
      if(_zz_30)begin
        img_reg_array_28_34_imag <= _zz_135;
      end
      if(_zz_31)begin
        img_reg_array_29_34_imag <= _zz_135;
      end
      if(_zz_32)begin
        img_reg_array_30_34_imag <= _zz_135;
      end
      if(_zz_33)begin
        img_reg_array_31_34_imag <= _zz_135;
      end
      if(_zz_34)begin
        img_reg_array_32_34_imag <= _zz_135;
      end
      if(_zz_35)begin
        img_reg_array_33_34_imag <= _zz_135;
      end
      if(_zz_36)begin
        img_reg_array_34_34_imag <= _zz_135;
      end
      if(_zz_37)begin
        img_reg_array_35_34_imag <= _zz_135;
      end
      if(_zz_38)begin
        img_reg_array_36_34_imag <= _zz_135;
      end
      if(_zz_39)begin
        img_reg_array_37_34_imag <= _zz_135;
      end
      if(_zz_40)begin
        img_reg_array_38_34_imag <= _zz_135;
      end
      if(_zz_41)begin
        img_reg_array_39_34_imag <= _zz_135;
      end
      if(_zz_42)begin
        img_reg_array_40_34_imag <= _zz_135;
      end
      if(_zz_43)begin
        img_reg_array_41_34_imag <= _zz_135;
      end
      if(_zz_44)begin
        img_reg_array_42_34_imag <= _zz_135;
      end
      if(_zz_45)begin
        img_reg_array_43_34_imag <= _zz_135;
      end
      if(_zz_46)begin
        img_reg_array_44_34_imag <= _zz_135;
      end
      if(_zz_47)begin
        img_reg_array_45_34_imag <= _zz_135;
      end
      if(_zz_48)begin
        img_reg_array_46_34_imag <= _zz_135;
      end
      if(_zz_49)begin
        img_reg_array_47_34_imag <= _zz_135;
      end
      if(_zz_50)begin
        img_reg_array_48_34_imag <= _zz_135;
      end
      if(_zz_51)begin
        img_reg_array_49_34_imag <= _zz_135;
      end
      if(_zz_52)begin
        img_reg_array_50_34_imag <= _zz_135;
      end
      if(_zz_53)begin
        img_reg_array_51_34_imag <= _zz_135;
      end
      if(_zz_54)begin
        img_reg_array_52_34_imag <= _zz_135;
      end
      if(_zz_55)begin
        img_reg_array_53_34_imag <= _zz_135;
      end
      if(_zz_56)begin
        img_reg_array_54_34_imag <= _zz_135;
      end
      if(_zz_57)begin
        img_reg_array_55_34_imag <= _zz_135;
      end
      if(_zz_58)begin
        img_reg_array_56_34_imag <= _zz_135;
      end
      if(_zz_59)begin
        img_reg_array_57_34_imag <= _zz_135;
      end
      if(_zz_60)begin
        img_reg_array_58_34_imag <= _zz_135;
      end
      if(_zz_61)begin
        img_reg_array_59_34_imag <= _zz_135;
      end
      if(_zz_62)begin
        img_reg_array_60_34_imag <= _zz_135;
      end
      if(_zz_63)begin
        img_reg_array_61_34_imag <= _zz_135;
      end
      if(_zz_64)begin
        img_reg_array_62_34_imag <= _zz_135;
      end
      if(_zz_65)begin
        img_reg_array_63_34_imag <= _zz_135;
      end
      if(_zz_2)begin
        img_reg_array_0_35_real <= _zz_136;
      end
      if(_zz_3)begin
        img_reg_array_1_35_real <= _zz_136;
      end
      if(_zz_4)begin
        img_reg_array_2_35_real <= _zz_136;
      end
      if(_zz_5)begin
        img_reg_array_3_35_real <= _zz_136;
      end
      if(_zz_6)begin
        img_reg_array_4_35_real <= _zz_136;
      end
      if(_zz_7)begin
        img_reg_array_5_35_real <= _zz_136;
      end
      if(_zz_8)begin
        img_reg_array_6_35_real <= _zz_136;
      end
      if(_zz_9)begin
        img_reg_array_7_35_real <= _zz_136;
      end
      if(_zz_10)begin
        img_reg_array_8_35_real <= _zz_136;
      end
      if(_zz_11)begin
        img_reg_array_9_35_real <= _zz_136;
      end
      if(_zz_12)begin
        img_reg_array_10_35_real <= _zz_136;
      end
      if(_zz_13)begin
        img_reg_array_11_35_real <= _zz_136;
      end
      if(_zz_14)begin
        img_reg_array_12_35_real <= _zz_136;
      end
      if(_zz_15)begin
        img_reg_array_13_35_real <= _zz_136;
      end
      if(_zz_16)begin
        img_reg_array_14_35_real <= _zz_136;
      end
      if(_zz_17)begin
        img_reg_array_15_35_real <= _zz_136;
      end
      if(_zz_18)begin
        img_reg_array_16_35_real <= _zz_136;
      end
      if(_zz_19)begin
        img_reg_array_17_35_real <= _zz_136;
      end
      if(_zz_20)begin
        img_reg_array_18_35_real <= _zz_136;
      end
      if(_zz_21)begin
        img_reg_array_19_35_real <= _zz_136;
      end
      if(_zz_22)begin
        img_reg_array_20_35_real <= _zz_136;
      end
      if(_zz_23)begin
        img_reg_array_21_35_real <= _zz_136;
      end
      if(_zz_24)begin
        img_reg_array_22_35_real <= _zz_136;
      end
      if(_zz_25)begin
        img_reg_array_23_35_real <= _zz_136;
      end
      if(_zz_26)begin
        img_reg_array_24_35_real <= _zz_136;
      end
      if(_zz_27)begin
        img_reg_array_25_35_real <= _zz_136;
      end
      if(_zz_28)begin
        img_reg_array_26_35_real <= _zz_136;
      end
      if(_zz_29)begin
        img_reg_array_27_35_real <= _zz_136;
      end
      if(_zz_30)begin
        img_reg_array_28_35_real <= _zz_136;
      end
      if(_zz_31)begin
        img_reg_array_29_35_real <= _zz_136;
      end
      if(_zz_32)begin
        img_reg_array_30_35_real <= _zz_136;
      end
      if(_zz_33)begin
        img_reg_array_31_35_real <= _zz_136;
      end
      if(_zz_34)begin
        img_reg_array_32_35_real <= _zz_136;
      end
      if(_zz_35)begin
        img_reg_array_33_35_real <= _zz_136;
      end
      if(_zz_36)begin
        img_reg_array_34_35_real <= _zz_136;
      end
      if(_zz_37)begin
        img_reg_array_35_35_real <= _zz_136;
      end
      if(_zz_38)begin
        img_reg_array_36_35_real <= _zz_136;
      end
      if(_zz_39)begin
        img_reg_array_37_35_real <= _zz_136;
      end
      if(_zz_40)begin
        img_reg_array_38_35_real <= _zz_136;
      end
      if(_zz_41)begin
        img_reg_array_39_35_real <= _zz_136;
      end
      if(_zz_42)begin
        img_reg_array_40_35_real <= _zz_136;
      end
      if(_zz_43)begin
        img_reg_array_41_35_real <= _zz_136;
      end
      if(_zz_44)begin
        img_reg_array_42_35_real <= _zz_136;
      end
      if(_zz_45)begin
        img_reg_array_43_35_real <= _zz_136;
      end
      if(_zz_46)begin
        img_reg_array_44_35_real <= _zz_136;
      end
      if(_zz_47)begin
        img_reg_array_45_35_real <= _zz_136;
      end
      if(_zz_48)begin
        img_reg_array_46_35_real <= _zz_136;
      end
      if(_zz_49)begin
        img_reg_array_47_35_real <= _zz_136;
      end
      if(_zz_50)begin
        img_reg_array_48_35_real <= _zz_136;
      end
      if(_zz_51)begin
        img_reg_array_49_35_real <= _zz_136;
      end
      if(_zz_52)begin
        img_reg_array_50_35_real <= _zz_136;
      end
      if(_zz_53)begin
        img_reg_array_51_35_real <= _zz_136;
      end
      if(_zz_54)begin
        img_reg_array_52_35_real <= _zz_136;
      end
      if(_zz_55)begin
        img_reg_array_53_35_real <= _zz_136;
      end
      if(_zz_56)begin
        img_reg_array_54_35_real <= _zz_136;
      end
      if(_zz_57)begin
        img_reg_array_55_35_real <= _zz_136;
      end
      if(_zz_58)begin
        img_reg_array_56_35_real <= _zz_136;
      end
      if(_zz_59)begin
        img_reg_array_57_35_real <= _zz_136;
      end
      if(_zz_60)begin
        img_reg_array_58_35_real <= _zz_136;
      end
      if(_zz_61)begin
        img_reg_array_59_35_real <= _zz_136;
      end
      if(_zz_62)begin
        img_reg_array_60_35_real <= _zz_136;
      end
      if(_zz_63)begin
        img_reg_array_61_35_real <= _zz_136;
      end
      if(_zz_64)begin
        img_reg_array_62_35_real <= _zz_136;
      end
      if(_zz_65)begin
        img_reg_array_63_35_real <= _zz_136;
      end
      if(_zz_2)begin
        img_reg_array_0_35_imag <= _zz_137;
      end
      if(_zz_3)begin
        img_reg_array_1_35_imag <= _zz_137;
      end
      if(_zz_4)begin
        img_reg_array_2_35_imag <= _zz_137;
      end
      if(_zz_5)begin
        img_reg_array_3_35_imag <= _zz_137;
      end
      if(_zz_6)begin
        img_reg_array_4_35_imag <= _zz_137;
      end
      if(_zz_7)begin
        img_reg_array_5_35_imag <= _zz_137;
      end
      if(_zz_8)begin
        img_reg_array_6_35_imag <= _zz_137;
      end
      if(_zz_9)begin
        img_reg_array_7_35_imag <= _zz_137;
      end
      if(_zz_10)begin
        img_reg_array_8_35_imag <= _zz_137;
      end
      if(_zz_11)begin
        img_reg_array_9_35_imag <= _zz_137;
      end
      if(_zz_12)begin
        img_reg_array_10_35_imag <= _zz_137;
      end
      if(_zz_13)begin
        img_reg_array_11_35_imag <= _zz_137;
      end
      if(_zz_14)begin
        img_reg_array_12_35_imag <= _zz_137;
      end
      if(_zz_15)begin
        img_reg_array_13_35_imag <= _zz_137;
      end
      if(_zz_16)begin
        img_reg_array_14_35_imag <= _zz_137;
      end
      if(_zz_17)begin
        img_reg_array_15_35_imag <= _zz_137;
      end
      if(_zz_18)begin
        img_reg_array_16_35_imag <= _zz_137;
      end
      if(_zz_19)begin
        img_reg_array_17_35_imag <= _zz_137;
      end
      if(_zz_20)begin
        img_reg_array_18_35_imag <= _zz_137;
      end
      if(_zz_21)begin
        img_reg_array_19_35_imag <= _zz_137;
      end
      if(_zz_22)begin
        img_reg_array_20_35_imag <= _zz_137;
      end
      if(_zz_23)begin
        img_reg_array_21_35_imag <= _zz_137;
      end
      if(_zz_24)begin
        img_reg_array_22_35_imag <= _zz_137;
      end
      if(_zz_25)begin
        img_reg_array_23_35_imag <= _zz_137;
      end
      if(_zz_26)begin
        img_reg_array_24_35_imag <= _zz_137;
      end
      if(_zz_27)begin
        img_reg_array_25_35_imag <= _zz_137;
      end
      if(_zz_28)begin
        img_reg_array_26_35_imag <= _zz_137;
      end
      if(_zz_29)begin
        img_reg_array_27_35_imag <= _zz_137;
      end
      if(_zz_30)begin
        img_reg_array_28_35_imag <= _zz_137;
      end
      if(_zz_31)begin
        img_reg_array_29_35_imag <= _zz_137;
      end
      if(_zz_32)begin
        img_reg_array_30_35_imag <= _zz_137;
      end
      if(_zz_33)begin
        img_reg_array_31_35_imag <= _zz_137;
      end
      if(_zz_34)begin
        img_reg_array_32_35_imag <= _zz_137;
      end
      if(_zz_35)begin
        img_reg_array_33_35_imag <= _zz_137;
      end
      if(_zz_36)begin
        img_reg_array_34_35_imag <= _zz_137;
      end
      if(_zz_37)begin
        img_reg_array_35_35_imag <= _zz_137;
      end
      if(_zz_38)begin
        img_reg_array_36_35_imag <= _zz_137;
      end
      if(_zz_39)begin
        img_reg_array_37_35_imag <= _zz_137;
      end
      if(_zz_40)begin
        img_reg_array_38_35_imag <= _zz_137;
      end
      if(_zz_41)begin
        img_reg_array_39_35_imag <= _zz_137;
      end
      if(_zz_42)begin
        img_reg_array_40_35_imag <= _zz_137;
      end
      if(_zz_43)begin
        img_reg_array_41_35_imag <= _zz_137;
      end
      if(_zz_44)begin
        img_reg_array_42_35_imag <= _zz_137;
      end
      if(_zz_45)begin
        img_reg_array_43_35_imag <= _zz_137;
      end
      if(_zz_46)begin
        img_reg_array_44_35_imag <= _zz_137;
      end
      if(_zz_47)begin
        img_reg_array_45_35_imag <= _zz_137;
      end
      if(_zz_48)begin
        img_reg_array_46_35_imag <= _zz_137;
      end
      if(_zz_49)begin
        img_reg_array_47_35_imag <= _zz_137;
      end
      if(_zz_50)begin
        img_reg_array_48_35_imag <= _zz_137;
      end
      if(_zz_51)begin
        img_reg_array_49_35_imag <= _zz_137;
      end
      if(_zz_52)begin
        img_reg_array_50_35_imag <= _zz_137;
      end
      if(_zz_53)begin
        img_reg_array_51_35_imag <= _zz_137;
      end
      if(_zz_54)begin
        img_reg_array_52_35_imag <= _zz_137;
      end
      if(_zz_55)begin
        img_reg_array_53_35_imag <= _zz_137;
      end
      if(_zz_56)begin
        img_reg_array_54_35_imag <= _zz_137;
      end
      if(_zz_57)begin
        img_reg_array_55_35_imag <= _zz_137;
      end
      if(_zz_58)begin
        img_reg_array_56_35_imag <= _zz_137;
      end
      if(_zz_59)begin
        img_reg_array_57_35_imag <= _zz_137;
      end
      if(_zz_60)begin
        img_reg_array_58_35_imag <= _zz_137;
      end
      if(_zz_61)begin
        img_reg_array_59_35_imag <= _zz_137;
      end
      if(_zz_62)begin
        img_reg_array_60_35_imag <= _zz_137;
      end
      if(_zz_63)begin
        img_reg_array_61_35_imag <= _zz_137;
      end
      if(_zz_64)begin
        img_reg_array_62_35_imag <= _zz_137;
      end
      if(_zz_65)begin
        img_reg_array_63_35_imag <= _zz_137;
      end
      if(_zz_2)begin
        img_reg_array_0_36_real <= _zz_138;
      end
      if(_zz_3)begin
        img_reg_array_1_36_real <= _zz_138;
      end
      if(_zz_4)begin
        img_reg_array_2_36_real <= _zz_138;
      end
      if(_zz_5)begin
        img_reg_array_3_36_real <= _zz_138;
      end
      if(_zz_6)begin
        img_reg_array_4_36_real <= _zz_138;
      end
      if(_zz_7)begin
        img_reg_array_5_36_real <= _zz_138;
      end
      if(_zz_8)begin
        img_reg_array_6_36_real <= _zz_138;
      end
      if(_zz_9)begin
        img_reg_array_7_36_real <= _zz_138;
      end
      if(_zz_10)begin
        img_reg_array_8_36_real <= _zz_138;
      end
      if(_zz_11)begin
        img_reg_array_9_36_real <= _zz_138;
      end
      if(_zz_12)begin
        img_reg_array_10_36_real <= _zz_138;
      end
      if(_zz_13)begin
        img_reg_array_11_36_real <= _zz_138;
      end
      if(_zz_14)begin
        img_reg_array_12_36_real <= _zz_138;
      end
      if(_zz_15)begin
        img_reg_array_13_36_real <= _zz_138;
      end
      if(_zz_16)begin
        img_reg_array_14_36_real <= _zz_138;
      end
      if(_zz_17)begin
        img_reg_array_15_36_real <= _zz_138;
      end
      if(_zz_18)begin
        img_reg_array_16_36_real <= _zz_138;
      end
      if(_zz_19)begin
        img_reg_array_17_36_real <= _zz_138;
      end
      if(_zz_20)begin
        img_reg_array_18_36_real <= _zz_138;
      end
      if(_zz_21)begin
        img_reg_array_19_36_real <= _zz_138;
      end
      if(_zz_22)begin
        img_reg_array_20_36_real <= _zz_138;
      end
      if(_zz_23)begin
        img_reg_array_21_36_real <= _zz_138;
      end
      if(_zz_24)begin
        img_reg_array_22_36_real <= _zz_138;
      end
      if(_zz_25)begin
        img_reg_array_23_36_real <= _zz_138;
      end
      if(_zz_26)begin
        img_reg_array_24_36_real <= _zz_138;
      end
      if(_zz_27)begin
        img_reg_array_25_36_real <= _zz_138;
      end
      if(_zz_28)begin
        img_reg_array_26_36_real <= _zz_138;
      end
      if(_zz_29)begin
        img_reg_array_27_36_real <= _zz_138;
      end
      if(_zz_30)begin
        img_reg_array_28_36_real <= _zz_138;
      end
      if(_zz_31)begin
        img_reg_array_29_36_real <= _zz_138;
      end
      if(_zz_32)begin
        img_reg_array_30_36_real <= _zz_138;
      end
      if(_zz_33)begin
        img_reg_array_31_36_real <= _zz_138;
      end
      if(_zz_34)begin
        img_reg_array_32_36_real <= _zz_138;
      end
      if(_zz_35)begin
        img_reg_array_33_36_real <= _zz_138;
      end
      if(_zz_36)begin
        img_reg_array_34_36_real <= _zz_138;
      end
      if(_zz_37)begin
        img_reg_array_35_36_real <= _zz_138;
      end
      if(_zz_38)begin
        img_reg_array_36_36_real <= _zz_138;
      end
      if(_zz_39)begin
        img_reg_array_37_36_real <= _zz_138;
      end
      if(_zz_40)begin
        img_reg_array_38_36_real <= _zz_138;
      end
      if(_zz_41)begin
        img_reg_array_39_36_real <= _zz_138;
      end
      if(_zz_42)begin
        img_reg_array_40_36_real <= _zz_138;
      end
      if(_zz_43)begin
        img_reg_array_41_36_real <= _zz_138;
      end
      if(_zz_44)begin
        img_reg_array_42_36_real <= _zz_138;
      end
      if(_zz_45)begin
        img_reg_array_43_36_real <= _zz_138;
      end
      if(_zz_46)begin
        img_reg_array_44_36_real <= _zz_138;
      end
      if(_zz_47)begin
        img_reg_array_45_36_real <= _zz_138;
      end
      if(_zz_48)begin
        img_reg_array_46_36_real <= _zz_138;
      end
      if(_zz_49)begin
        img_reg_array_47_36_real <= _zz_138;
      end
      if(_zz_50)begin
        img_reg_array_48_36_real <= _zz_138;
      end
      if(_zz_51)begin
        img_reg_array_49_36_real <= _zz_138;
      end
      if(_zz_52)begin
        img_reg_array_50_36_real <= _zz_138;
      end
      if(_zz_53)begin
        img_reg_array_51_36_real <= _zz_138;
      end
      if(_zz_54)begin
        img_reg_array_52_36_real <= _zz_138;
      end
      if(_zz_55)begin
        img_reg_array_53_36_real <= _zz_138;
      end
      if(_zz_56)begin
        img_reg_array_54_36_real <= _zz_138;
      end
      if(_zz_57)begin
        img_reg_array_55_36_real <= _zz_138;
      end
      if(_zz_58)begin
        img_reg_array_56_36_real <= _zz_138;
      end
      if(_zz_59)begin
        img_reg_array_57_36_real <= _zz_138;
      end
      if(_zz_60)begin
        img_reg_array_58_36_real <= _zz_138;
      end
      if(_zz_61)begin
        img_reg_array_59_36_real <= _zz_138;
      end
      if(_zz_62)begin
        img_reg_array_60_36_real <= _zz_138;
      end
      if(_zz_63)begin
        img_reg_array_61_36_real <= _zz_138;
      end
      if(_zz_64)begin
        img_reg_array_62_36_real <= _zz_138;
      end
      if(_zz_65)begin
        img_reg_array_63_36_real <= _zz_138;
      end
      if(_zz_2)begin
        img_reg_array_0_36_imag <= _zz_139;
      end
      if(_zz_3)begin
        img_reg_array_1_36_imag <= _zz_139;
      end
      if(_zz_4)begin
        img_reg_array_2_36_imag <= _zz_139;
      end
      if(_zz_5)begin
        img_reg_array_3_36_imag <= _zz_139;
      end
      if(_zz_6)begin
        img_reg_array_4_36_imag <= _zz_139;
      end
      if(_zz_7)begin
        img_reg_array_5_36_imag <= _zz_139;
      end
      if(_zz_8)begin
        img_reg_array_6_36_imag <= _zz_139;
      end
      if(_zz_9)begin
        img_reg_array_7_36_imag <= _zz_139;
      end
      if(_zz_10)begin
        img_reg_array_8_36_imag <= _zz_139;
      end
      if(_zz_11)begin
        img_reg_array_9_36_imag <= _zz_139;
      end
      if(_zz_12)begin
        img_reg_array_10_36_imag <= _zz_139;
      end
      if(_zz_13)begin
        img_reg_array_11_36_imag <= _zz_139;
      end
      if(_zz_14)begin
        img_reg_array_12_36_imag <= _zz_139;
      end
      if(_zz_15)begin
        img_reg_array_13_36_imag <= _zz_139;
      end
      if(_zz_16)begin
        img_reg_array_14_36_imag <= _zz_139;
      end
      if(_zz_17)begin
        img_reg_array_15_36_imag <= _zz_139;
      end
      if(_zz_18)begin
        img_reg_array_16_36_imag <= _zz_139;
      end
      if(_zz_19)begin
        img_reg_array_17_36_imag <= _zz_139;
      end
      if(_zz_20)begin
        img_reg_array_18_36_imag <= _zz_139;
      end
      if(_zz_21)begin
        img_reg_array_19_36_imag <= _zz_139;
      end
      if(_zz_22)begin
        img_reg_array_20_36_imag <= _zz_139;
      end
      if(_zz_23)begin
        img_reg_array_21_36_imag <= _zz_139;
      end
      if(_zz_24)begin
        img_reg_array_22_36_imag <= _zz_139;
      end
      if(_zz_25)begin
        img_reg_array_23_36_imag <= _zz_139;
      end
      if(_zz_26)begin
        img_reg_array_24_36_imag <= _zz_139;
      end
      if(_zz_27)begin
        img_reg_array_25_36_imag <= _zz_139;
      end
      if(_zz_28)begin
        img_reg_array_26_36_imag <= _zz_139;
      end
      if(_zz_29)begin
        img_reg_array_27_36_imag <= _zz_139;
      end
      if(_zz_30)begin
        img_reg_array_28_36_imag <= _zz_139;
      end
      if(_zz_31)begin
        img_reg_array_29_36_imag <= _zz_139;
      end
      if(_zz_32)begin
        img_reg_array_30_36_imag <= _zz_139;
      end
      if(_zz_33)begin
        img_reg_array_31_36_imag <= _zz_139;
      end
      if(_zz_34)begin
        img_reg_array_32_36_imag <= _zz_139;
      end
      if(_zz_35)begin
        img_reg_array_33_36_imag <= _zz_139;
      end
      if(_zz_36)begin
        img_reg_array_34_36_imag <= _zz_139;
      end
      if(_zz_37)begin
        img_reg_array_35_36_imag <= _zz_139;
      end
      if(_zz_38)begin
        img_reg_array_36_36_imag <= _zz_139;
      end
      if(_zz_39)begin
        img_reg_array_37_36_imag <= _zz_139;
      end
      if(_zz_40)begin
        img_reg_array_38_36_imag <= _zz_139;
      end
      if(_zz_41)begin
        img_reg_array_39_36_imag <= _zz_139;
      end
      if(_zz_42)begin
        img_reg_array_40_36_imag <= _zz_139;
      end
      if(_zz_43)begin
        img_reg_array_41_36_imag <= _zz_139;
      end
      if(_zz_44)begin
        img_reg_array_42_36_imag <= _zz_139;
      end
      if(_zz_45)begin
        img_reg_array_43_36_imag <= _zz_139;
      end
      if(_zz_46)begin
        img_reg_array_44_36_imag <= _zz_139;
      end
      if(_zz_47)begin
        img_reg_array_45_36_imag <= _zz_139;
      end
      if(_zz_48)begin
        img_reg_array_46_36_imag <= _zz_139;
      end
      if(_zz_49)begin
        img_reg_array_47_36_imag <= _zz_139;
      end
      if(_zz_50)begin
        img_reg_array_48_36_imag <= _zz_139;
      end
      if(_zz_51)begin
        img_reg_array_49_36_imag <= _zz_139;
      end
      if(_zz_52)begin
        img_reg_array_50_36_imag <= _zz_139;
      end
      if(_zz_53)begin
        img_reg_array_51_36_imag <= _zz_139;
      end
      if(_zz_54)begin
        img_reg_array_52_36_imag <= _zz_139;
      end
      if(_zz_55)begin
        img_reg_array_53_36_imag <= _zz_139;
      end
      if(_zz_56)begin
        img_reg_array_54_36_imag <= _zz_139;
      end
      if(_zz_57)begin
        img_reg_array_55_36_imag <= _zz_139;
      end
      if(_zz_58)begin
        img_reg_array_56_36_imag <= _zz_139;
      end
      if(_zz_59)begin
        img_reg_array_57_36_imag <= _zz_139;
      end
      if(_zz_60)begin
        img_reg_array_58_36_imag <= _zz_139;
      end
      if(_zz_61)begin
        img_reg_array_59_36_imag <= _zz_139;
      end
      if(_zz_62)begin
        img_reg_array_60_36_imag <= _zz_139;
      end
      if(_zz_63)begin
        img_reg_array_61_36_imag <= _zz_139;
      end
      if(_zz_64)begin
        img_reg_array_62_36_imag <= _zz_139;
      end
      if(_zz_65)begin
        img_reg_array_63_36_imag <= _zz_139;
      end
      if(_zz_2)begin
        img_reg_array_0_37_real <= _zz_140;
      end
      if(_zz_3)begin
        img_reg_array_1_37_real <= _zz_140;
      end
      if(_zz_4)begin
        img_reg_array_2_37_real <= _zz_140;
      end
      if(_zz_5)begin
        img_reg_array_3_37_real <= _zz_140;
      end
      if(_zz_6)begin
        img_reg_array_4_37_real <= _zz_140;
      end
      if(_zz_7)begin
        img_reg_array_5_37_real <= _zz_140;
      end
      if(_zz_8)begin
        img_reg_array_6_37_real <= _zz_140;
      end
      if(_zz_9)begin
        img_reg_array_7_37_real <= _zz_140;
      end
      if(_zz_10)begin
        img_reg_array_8_37_real <= _zz_140;
      end
      if(_zz_11)begin
        img_reg_array_9_37_real <= _zz_140;
      end
      if(_zz_12)begin
        img_reg_array_10_37_real <= _zz_140;
      end
      if(_zz_13)begin
        img_reg_array_11_37_real <= _zz_140;
      end
      if(_zz_14)begin
        img_reg_array_12_37_real <= _zz_140;
      end
      if(_zz_15)begin
        img_reg_array_13_37_real <= _zz_140;
      end
      if(_zz_16)begin
        img_reg_array_14_37_real <= _zz_140;
      end
      if(_zz_17)begin
        img_reg_array_15_37_real <= _zz_140;
      end
      if(_zz_18)begin
        img_reg_array_16_37_real <= _zz_140;
      end
      if(_zz_19)begin
        img_reg_array_17_37_real <= _zz_140;
      end
      if(_zz_20)begin
        img_reg_array_18_37_real <= _zz_140;
      end
      if(_zz_21)begin
        img_reg_array_19_37_real <= _zz_140;
      end
      if(_zz_22)begin
        img_reg_array_20_37_real <= _zz_140;
      end
      if(_zz_23)begin
        img_reg_array_21_37_real <= _zz_140;
      end
      if(_zz_24)begin
        img_reg_array_22_37_real <= _zz_140;
      end
      if(_zz_25)begin
        img_reg_array_23_37_real <= _zz_140;
      end
      if(_zz_26)begin
        img_reg_array_24_37_real <= _zz_140;
      end
      if(_zz_27)begin
        img_reg_array_25_37_real <= _zz_140;
      end
      if(_zz_28)begin
        img_reg_array_26_37_real <= _zz_140;
      end
      if(_zz_29)begin
        img_reg_array_27_37_real <= _zz_140;
      end
      if(_zz_30)begin
        img_reg_array_28_37_real <= _zz_140;
      end
      if(_zz_31)begin
        img_reg_array_29_37_real <= _zz_140;
      end
      if(_zz_32)begin
        img_reg_array_30_37_real <= _zz_140;
      end
      if(_zz_33)begin
        img_reg_array_31_37_real <= _zz_140;
      end
      if(_zz_34)begin
        img_reg_array_32_37_real <= _zz_140;
      end
      if(_zz_35)begin
        img_reg_array_33_37_real <= _zz_140;
      end
      if(_zz_36)begin
        img_reg_array_34_37_real <= _zz_140;
      end
      if(_zz_37)begin
        img_reg_array_35_37_real <= _zz_140;
      end
      if(_zz_38)begin
        img_reg_array_36_37_real <= _zz_140;
      end
      if(_zz_39)begin
        img_reg_array_37_37_real <= _zz_140;
      end
      if(_zz_40)begin
        img_reg_array_38_37_real <= _zz_140;
      end
      if(_zz_41)begin
        img_reg_array_39_37_real <= _zz_140;
      end
      if(_zz_42)begin
        img_reg_array_40_37_real <= _zz_140;
      end
      if(_zz_43)begin
        img_reg_array_41_37_real <= _zz_140;
      end
      if(_zz_44)begin
        img_reg_array_42_37_real <= _zz_140;
      end
      if(_zz_45)begin
        img_reg_array_43_37_real <= _zz_140;
      end
      if(_zz_46)begin
        img_reg_array_44_37_real <= _zz_140;
      end
      if(_zz_47)begin
        img_reg_array_45_37_real <= _zz_140;
      end
      if(_zz_48)begin
        img_reg_array_46_37_real <= _zz_140;
      end
      if(_zz_49)begin
        img_reg_array_47_37_real <= _zz_140;
      end
      if(_zz_50)begin
        img_reg_array_48_37_real <= _zz_140;
      end
      if(_zz_51)begin
        img_reg_array_49_37_real <= _zz_140;
      end
      if(_zz_52)begin
        img_reg_array_50_37_real <= _zz_140;
      end
      if(_zz_53)begin
        img_reg_array_51_37_real <= _zz_140;
      end
      if(_zz_54)begin
        img_reg_array_52_37_real <= _zz_140;
      end
      if(_zz_55)begin
        img_reg_array_53_37_real <= _zz_140;
      end
      if(_zz_56)begin
        img_reg_array_54_37_real <= _zz_140;
      end
      if(_zz_57)begin
        img_reg_array_55_37_real <= _zz_140;
      end
      if(_zz_58)begin
        img_reg_array_56_37_real <= _zz_140;
      end
      if(_zz_59)begin
        img_reg_array_57_37_real <= _zz_140;
      end
      if(_zz_60)begin
        img_reg_array_58_37_real <= _zz_140;
      end
      if(_zz_61)begin
        img_reg_array_59_37_real <= _zz_140;
      end
      if(_zz_62)begin
        img_reg_array_60_37_real <= _zz_140;
      end
      if(_zz_63)begin
        img_reg_array_61_37_real <= _zz_140;
      end
      if(_zz_64)begin
        img_reg_array_62_37_real <= _zz_140;
      end
      if(_zz_65)begin
        img_reg_array_63_37_real <= _zz_140;
      end
      if(_zz_2)begin
        img_reg_array_0_37_imag <= _zz_141;
      end
      if(_zz_3)begin
        img_reg_array_1_37_imag <= _zz_141;
      end
      if(_zz_4)begin
        img_reg_array_2_37_imag <= _zz_141;
      end
      if(_zz_5)begin
        img_reg_array_3_37_imag <= _zz_141;
      end
      if(_zz_6)begin
        img_reg_array_4_37_imag <= _zz_141;
      end
      if(_zz_7)begin
        img_reg_array_5_37_imag <= _zz_141;
      end
      if(_zz_8)begin
        img_reg_array_6_37_imag <= _zz_141;
      end
      if(_zz_9)begin
        img_reg_array_7_37_imag <= _zz_141;
      end
      if(_zz_10)begin
        img_reg_array_8_37_imag <= _zz_141;
      end
      if(_zz_11)begin
        img_reg_array_9_37_imag <= _zz_141;
      end
      if(_zz_12)begin
        img_reg_array_10_37_imag <= _zz_141;
      end
      if(_zz_13)begin
        img_reg_array_11_37_imag <= _zz_141;
      end
      if(_zz_14)begin
        img_reg_array_12_37_imag <= _zz_141;
      end
      if(_zz_15)begin
        img_reg_array_13_37_imag <= _zz_141;
      end
      if(_zz_16)begin
        img_reg_array_14_37_imag <= _zz_141;
      end
      if(_zz_17)begin
        img_reg_array_15_37_imag <= _zz_141;
      end
      if(_zz_18)begin
        img_reg_array_16_37_imag <= _zz_141;
      end
      if(_zz_19)begin
        img_reg_array_17_37_imag <= _zz_141;
      end
      if(_zz_20)begin
        img_reg_array_18_37_imag <= _zz_141;
      end
      if(_zz_21)begin
        img_reg_array_19_37_imag <= _zz_141;
      end
      if(_zz_22)begin
        img_reg_array_20_37_imag <= _zz_141;
      end
      if(_zz_23)begin
        img_reg_array_21_37_imag <= _zz_141;
      end
      if(_zz_24)begin
        img_reg_array_22_37_imag <= _zz_141;
      end
      if(_zz_25)begin
        img_reg_array_23_37_imag <= _zz_141;
      end
      if(_zz_26)begin
        img_reg_array_24_37_imag <= _zz_141;
      end
      if(_zz_27)begin
        img_reg_array_25_37_imag <= _zz_141;
      end
      if(_zz_28)begin
        img_reg_array_26_37_imag <= _zz_141;
      end
      if(_zz_29)begin
        img_reg_array_27_37_imag <= _zz_141;
      end
      if(_zz_30)begin
        img_reg_array_28_37_imag <= _zz_141;
      end
      if(_zz_31)begin
        img_reg_array_29_37_imag <= _zz_141;
      end
      if(_zz_32)begin
        img_reg_array_30_37_imag <= _zz_141;
      end
      if(_zz_33)begin
        img_reg_array_31_37_imag <= _zz_141;
      end
      if(_zz_34)begin
        img_reg_array_32_37_imag <= _zz_141;
      end
      if(_zz_35)begin
        img_reg_array_33_37_imag <= _zz_141;
      end
      if(_zz_36)begin
        img_reg_array_34_37_imag <= _zz_141;
      end
      if(_zz_37)begin
        img_reg_array_35_37_imag <= _zz_141;
      end
      if(_zz_38)begin
        img_reg_array_36_37_imag <= _zz_141;
      end
      if(_zz_39)begin
        img_reg_array_37_37_imag <= _zz_141;
      end
      if(_zz_40)begin
        img_reg_array_38_37_imag <= _zz_141;
      end
      if(_zz_41)begin
        img_reg_array_39_37_imag <= _zz_141;
      end
      if(_zz_42)begin
        img_reg_array_40_37_imag <= _zz_141;
      end
      if(_zz_43)begin
        img_reg_array_41_37_imag <= _zz_141;
      end
      if(_zz_44)begin
        img_reg_array_42_37_imag <= _zz_141;
      end
      if(_zz_45)begin
        img_reg_array_43_37_imag <= _zz_141;
      end
      if(_zz_46)begin
        img_reg_array_44_37_imag <= _zz_141;
      end
      if(_zz_47)begin
        img_reg_array_45_37_imag <= _zz_141;
      end
      if(_zz_48)begin
        img_reg_array_46_37_imag <= _zz_141;
      end
      if(_zz_49)begin
        img_reg_array_47_37_imag <= _zz_141;
      end
      if(_zz_50)begin
        img_reg_array_48_37_imag <= _zz_141;
      end
      if(_zz_51)begin
        img_reg_array_49_37_imag <= _zz_141;
      end
      if(_zz_52)begin
        img_reg_array_50_37_imag <= _zz_141;
      end
      if(_zz_53)begin
        img_reg_array_51_37_imag <= _zz_141;
      end
      if(_zz_54)begin
        img_reg_array_52_37_imag <= _zz_141;
      end
      if(_zz_55)begin
        img_reg_array_53_37_imag <= _zz_141;
      end
      if(_zz_56)begin
        img_reg_array_54_37_imag <= _zz_141;
      end
      if(_zz_57)begin
        img_reg_array_55_37_imag <= _zz_141;
      end
      if(_zz_58)begin
        img_reg_array_56_37_imag <= _zz_141;
      end
      if(_zz_59)begin
        img_reg_array_57_37_imag <= _zz_141;
      end
      if(_zz_60)begin
        img_reg_array_58_37_imag <= _zz_141;
      end
      if(_zz_61)begin
        img_reg_array_59_37_imag <= _zz_141;
      end
      if(_zz_62)begin
        img_reg_array_60_37_imag <= _zz_141;
      end
      if(_zz_63)begin
        img_reg_array_61_37_imag <= _zz_141;
      end
      if(_zz_64)begin
        img_reg_array_62_37_imag <= _zz_141;
      end
      if(_zz_65)begin
        img_reg_array_63_37_imag <= _zz_141;
      end
      if(_zz_2)begin
        img_reg_array_0_38_real <= _zz_142;
      end
      if(_zz_3)begin
        img_reg_array_1_38_real <= _zz_142;
      end
      if(_zz_4)begin
        img_reg_array_2_38_real <= _zz_142;
      end
      if(_zz_5)begin
        img_reg_array_3_38_real <= _zz_142;
      end
      if(_zz_6)begin
        img_reg_array_4_38_real <= _zz_142;
      end
      if(_zz_7)begin
        img_reg_array_5_38_real <= _zz_142;
      end
      if(_zz_8)begin
        img_reg_array_6_38_real <= _zz_142;
      end
      if(_zz_9)begin
        img_reg_array_7_38_real <= _zz_142;
      end
      if(_zz_10)begin
        img_reg_array_8_38_real <= _zz_142;
      end
      if(_zz_11)begin
        img_reg_array_9_38_real <= _zz_142;
      end
      if(_zz_12)begin
        img_reg_array_10_38_real <= _zz_142;
      end
      if(_zz_13)begin
        img_reg_array_11_38_real <= _zz_142;
      end
      if(_zz_14)begin
        img_reg_array_12_38_real <= _zz_142;
      end
      if(_zz_15)begin
        img_reg_array_13_38_real <= _zz_142;
      end
      if(_zz_16)begin
        img_reg_array_14_38_real <= _zz_142;
      end
      if(_zz_17)begin
        img_reg_array_15_38_real <= _zz_142;
      end
      if(_zz_18)begin
        img_reg_array_16_38_real <= _zz_142;
      end
      if(_zz_19)begin
        img_reg_array_17_38_real <= _zz_142;
      end
      if(_zz_20)begin
        img_reg_array_18_38_real <= _zz_142;
      end
      if(_zz_21)begin
        img_reg_array_19_38_real <= _zz_142;
      end
      if(_zz_22)begin
        img_reg_array_20_38_real <= _zz_142;
      end
      if(_zz_23)begin
        img_reg_array_21_38_real <= _zz_142;
      end
      if(_zz_24)begin
        img_reg_array_22_38_real <= _zz_142;
      end
      if(_zz_25)begin
        img_reg_array_23_38_real <= _zz_142;
      end
      if(_zz_26)begin
        img_reg_array_24_38_real <= _zz_142;
      end
      if(_zz_27)begin
        img_reg_array_25_38_real <= _zz_142;
      end
      if(_zz_28)begin
        img_reg_array_26_38_real <= _zz_142;
      end
      if(_zz_29)begin
        img_reg_array_27_38_real <= _zz_142;
      end
      if(_zz_30)begin
        img_reg_array_28_38_real <= _zz_142;
      end
      if(_zz_31)begin
        img_reg_array_29_38_real <= _zz_142;
      end
      if(_zz_32)begin
        img_reg_array_30_38_real <= _zz_142;
      end
      if(_zz_33)begin
        img_reg_array_31_38_real <= _zz_142;
      end
      if(_zz_34)begin
        img_reg_array_32_38_real <= _zz_142;
      end
      if(_zz_35)begin
        img_reg_array_33_38_real <= _zz_142;
      end
      if(_zz_36)begin
        img_reg_array_34_38_real <= _zz_142;
      end
      if(_zz_37)begin
        img_reg_array_35_38_real <= _zz_142;
      end
      if(_zz_38)begin
        img_reg_array_36_38_real <= _zz_142;
      end
      if(_zz_39)begin
        img_reg_array_37_38_real <= _zz_142;
      end
      if(_zz_40)begin
        img_reg_array_38_38_real <= _zz_142;
      end
      if(_zz_41)begin
        img_reg_array_39_38_real <= _zz_142;
      end
      if(_zz_42)begin
        img_reg_array_40_38_real <= _zz_142;
      end
      if(_zz_43)begin
        img_reg_array_41_38_real <= _zz_142;
      end
      if(_zz_44)begin
        img_reg_array_42_38_real <= _zz_142;
      end
      if(_zz_45)begin
        img_reg_array_43_38_real <= _zz_142;
      end
      if(_zz_46)begin
        img_reg_array_44_38_real <= _zz_142;
      end
      if(_zz_47)begin
        img_reg_array_45_38_real <= _zz_142;
      end
      if(_zz_48)begin
        img_reg_array_46_38_real <= _zz_142;
      end
      if(_zz_49)begin
        img_reg_array_47_38_real <= _zz_142;
      end
      if(_zz_50)begin
        img_reg_array_48_38_real <= _zz_142;
      end
      if(_zz_51)begin
        img_reg_array_49_38_real <= _zz_142;
      end
      if(_zz_52)begin
        img_reg_array_50_38_real <= _zz_142;
      end
      if(_zz_53)begin
        img_reg_array_51_38_real <= _zz_142;
      end
      if(_zz_54)begin
        img_reg_array_52_38_real <= _zz_142;
      end
      if(_zz_55)begin
        img_reg_array_53_38_real <= _zz_142;
      end
      if(_zz_56)begin
        img_reg_array_54_38_real <= _zz_142;
      end
      if(_zz_57)begin
        img_reg_array_55_38_real <= _zz_142;
      end
      if(_zz_58)begin
        img_reg_array_56_38_real <= _zz_142;
      end
      if(_zz_59)begin
        img_reg_array_57_38_real <= _zz_142;
      end
      if(_zz_60)begin
        img_reg_array_58_38_real <= _zz_142;
      end
      if(_zz_61)begin
        img_reg_array_59_38_real <= _zz_142;
      end
      if(_zz_62)begin
        img_reg_array_60_38_real <= _zz_142;
      end
      if(_zz_63)begin
        img_reg_array_61_38_real <= _zz_142;
      end
      if(_zz_64)begin
        img_reg_array_62_38_real <= _zz_142;
      end
      if(_zz_65)begin
        img_reg_array_63_38_real <= _zz_142;
      end
      if(_zz_2)begin
        img_reg_array_0_38_imag <= _zz_143;
      end
      if(_zz_3)begin
        img_reg_array_1_38_imag <= _zz_143;
      end
      if(_zz_4)begin
        img_reg_array_2_38_imag <= _zz_143;
      end
      if(_zz_5)begin
        img_reg_array_3_38_imag <= _zz_143;
      end
      if(_zz_6)begin
        img_reg_array_4_38_imag <= _zz_143;
      end
      if(_zz_7)begin
        img_reg_array_5_38_imag <= _zz_143;
      end
      if(_zz_8)begin
        img_reg_array_6_38_imag <= _zz_143;
      end
      if(_zz_9)begin
        img_reg_array_7_38_imag <= _zz_143;
      end
      if(_zz_10)begin
        img_reg_array_8_38_imag <= _zz_143;
      end
      if(_zz_11)begin
        img_reg_array_9_38_imag <= _zz_143;
      end
      if(_zz_12)begin
        img_reg_array_10_38_imag <= _zz_143;
      end
      if(_zz_13)begin
        img_reg_array_11_38_imag <= _zz_143;
      end
      if(_zz_14)begin
        img_reg_array_12_38_imag <= _zz_143;
      end
      if(_zz_15)begin
        img_reg_array_13_38_imag <= _zz_143;
      end
      if(_zz_16)begin
        img_reg_array_14_38_imag <= _zz_143;
      end
      if(_zz_17)begin
        img_reg_array_15_38_imag <= _zz_143;
      end
      if(_zz_18)begin
        img_reg_array_16_38_imag <= _zz_143;
      end
      if(_zz_19)begin
        img_reg_array_17_38_imag <= _zz_143;
      end
      if(_zz_20)begin
        img_reg_array_18_38_imag <= _zz_143;
      end
      if(_zz_21)begin
        img_reg_array_19_38_imag <= _zz_143;
      end
      if(_zz_22)begin
        img_reg_array_20_38_imag <= _zz_143;
      end
      if(_zz_23)begin
        img_reg_array_21_38_imag <= _zz_143;
      end
      if(_zz_24)begin
        img_reg_array_22_38_imag <= _zz_143;
      end
      if(_zz_25)begin
        img_reg_array_23_38_imag <= _zz_143;
      end
      if(_zz_26)begin
        img_reg_array_24_38_imag <= _zz_143;
      end
      if(_zz_27)begin
        img_reg_array_25_38_imag <= _zz_143;
      end
      if(_zz_28)begin
        img_reg_array_26_38_imag <= _zz_143;
      end
      if(_zz_29)begin
        img_reg_array_27_38_imag <= _zz_143;
      end
      if(_zz_30)begin
        img_reg_array_28_38_imag <= _zz_143;
      end
      if(_zz_31)begin
        img_reg_array_29_38_imag <= _zz_143;
      end
      if(_zz_32)begin
        img_reg_array_30_38_imag <= _zz_143;
      end
      if(_zz_33)begin
        img_reg_array_31_38_imag <= _zz_143;
      end
      if(_zz_34)begin
        img_reg_array_32_38_imag <= _zz_143;
      end
      if(_zz_35)begin
        img_reg_array_33_38_imag <= _zz_143;
      end
      if(_zz_36)begin
        img_reg_array_34_38_imag <= _zz_143;
      end
      if(_zz_37)begin
        img_reg_array_35_38_imag <= _zz_143;
      end
      if(_zz_38)begin
        img_reg_array_36_38_imag <= _zz_143;
      end
      if(_zz_39)begin
        img_reg_array_37_38_imag <= _zz_143;
      end
      if(_zz_40)begin
        img_reg_array_38_38_imag <= _zz_143;
      end
      if(_zz_41)begin
        img_reg_array_39_38_imag <= _zz_143;
      end
      if(_zz_42)begin
        img_reg_array_40_38_imag <= _zz_143;
      end
      if(_zz_43)begin
        img_reg_array_41_38_imag <= _zz_143;
      end
      if(_zz_44)begin
        img_reg_array_42_38_imag <= _zz_143;
      end
      if(_zz_45)begin
        img_reg_array_43_38_imag <= _zz_143;
      end
      if(_zz_46)begin
        img_reg_array_44_38_imag <= _zz_143;
      end
      if(_zz_47)begin
        img_reg_array_45_38_imag <= _zz_143;
      end
      if(_zz_48)begin
        img_reg_array_46_38_imag <= _zz_143;
      end
      if(_zz_49)begin
        img_reg_array_47_38_imag <= _zz_143;
      end
      if(_zz_50)begin
        img_reg_array_48_38_imag <= _zz_143;
      end
      if(_zz_51)begin
        img_reg_array_49_38_imag <= _zz_143;
      end
      if(_zz_52)begin
        img_reg_array_50_38_imag <= _zz_143;
      end
      if(_zz_53)begin
        img_reg_array_51_38_imag <= _zz_143;
      end
      if(_zz_54)begin
        img_reg_array_52_38_imag <= _zz_143;
      end
      if(_zz_55)begin
        img_reg_array_53_38_imag <= _zz_143;
      end
      if(_zz_56)begin
        img_reg_array_54_38_imag <= _zz_143;
      end
      if(_zz_57)begin
        img_reg_array_55_38_imag <= _zz_143;
      end
      if(_zz_58)begin
        img_reg_array_56_38_imag <= _zz_143;
      end
      if(_zz_59)begin
        img_reg_array_57_38_imag <= _zz_143;
      end
      if(_zz_60)begin
        img_reg_array_58_38_imag <= _zz_143;
      end
      if(_zz_61)begin
        img_reg_array_59_38_imag <= _zz_143;
      end
      if(_zz_62)begin
        img_reg_array_60_38_imag <= _zz_143;
      end
      if(_zz_63)begin
        img_reg_array_61_38_imag <= _zz_143;
      end
      if(_zz_64)begin
        img_reg_array_62_38_imag <= _zz_143;
      end
      if(_zz_65)begin
        img_reg_array_63_38_imag <= _zz_143;
      end
      if(_zz_2)begin
        img_reg_array_0_39_real <= _zz_144;
      end
      if(_zz_3)begin
        img_reg_array_1_39_real <= _zz_144;
      end
      if(_zz_4)begin
        img_reg_array_2_39_real <= _zz_144;
      end
      if(_zz_5)begin
        img_reg_array_3_39_real <= _zz_144;
      end
      if(_zz_6)begin
        img_reg_array_4_39_real <= _zz_144;
      end
      if(_zz_7)begin
        img_reg_array_5_39_real <= _zz_144;
      end
      if(_zz_8)begin
        img_reg_array_6_39_real <= _zz_144;
      end
      if(_zz_9)begin
        img_reg_array_7_39_real <= _zz_144;
      end
      if(_zz_10)begin
        img_reg_array_8_39_real <= _zz_144;
      end
      if(_zz_11)begin
        img_reg_array_9_39_real <= _zz_144;
      end
      if(_zz_12)begin
        img_reg_array_10_39_real <= _zz_144;
      end
      if(_zz_13)begin
        img_reg_array_11_39_real <= _zz_144;
      end
      if(_zz_14)begin
        img_reg_array_12_39_real <= _zz_144;
      end
      if(_zz_15)begin
        img_reg_array_13_39_real <= _zz_144;
      end
      if(_zz_16)begin
        img_reg_array_14_39_real <= _zz_144;
      end
      if(_zz_17)begin
        img_reg_array_15_39_real <= _zz_144;
      end
      if(_zz_18)begin
        img_reg_array_16_39_real <= _zz_144;
      end
      if(_zz_19)begin
        img_reg_array_17_39_real <= _zz_144;
      end
      if(_zz_20)begin
        img_reg_array_18_39_real <= _zz_144;
      end
      if(_zz_21)begin
        img_reg_array_19_39_real <= _zz_144;
      end
      if(_zz_22)begin
        img_reg_array_20_39_real <= _zz_144;
      end
      if(_zz_23)begin
        img_reg_array_21_39_real <= _zz_144;
      end
      if(_zz_24)begin
        img_reg_array_22_39_real <= _zz_144;
      end
      if(_zz_25)begin
        img_reg_array_23_39_real <= _zz_144;
      end
      if(_zz_26)begin
        img_reg_array_24_39_real <= _zz_144;
      end
      if(_zz_27)begin
        img_reg_array_25_39_real <= _zz_144;
      end
      if(_zz_28)begin
        img_reg_array_26_39_real <= _zz_144;
      end
      if(_zz_29)begin
        img_reg_array_27_39_real <= _zz_144;
      end
      if(_zz_30)begin
        img_reg_array_28_39_real <= _zz_144;
      end
      if(_zz_31)begin
        img_reg_array_29_39_real <= _zz_144;
      end
      if(_zz_32)begin
        img_reg_array_30_39_real <= _zz_144;
      end
      if(_zz_33)begin
        img_reg_array_31_39_real <= _zz_144;
      end
      if(_zz_34)begin
        img_reg_array_32_39_real <= _zz_144;
      end
      if(_zz_35)begin
        img_reg_array_33_39_real <= _zz_144;
      end
      if(_zz_36)begin
        img_reg_array_34_39_real <= _zz_144;
      end
      if(_zz_37)begin
        img_reg_array_35_39_real <= _zz_144;
      end
      if(_zz_38)begin
        img_reg_array_36_39_real <= _zz_144;
      end
      if(_zz_39)begin
        img_reg_array_37_39_real <= _zz_144;
      end
      if(_zz_40)begin
        img_reg_array_38_39_real <= _zz_144;
      end
      if(_zz_41)begin
        img_reg_array_39_39_real <= _zz_144;
      end
      if(_zz_42)begin
        img_reg_array_40_39_real <= _zz_144;
      end
      if(_zz_43)begin
        img_reg_array_41_39_real <= _zz_144;
      end
      if(_zz_44)begin
        img_reg_array_42_39_real <= _zz_144;
      end
      if(_zz_45)begin
        img_reg_array_43_39_real <= _zz_144;
      end
      if(_zz_46)begin
        img_reg_array_44_39_real <= _zz_144;
      end
      if(_zz_47)begin
        img_reg_array_45_39_real <= _zz_144;
      end
      if(_zz_48)begin
        img_reg_array_46_39_real <= _zz_144;
      end
      if(_zz_49)begin
        img_reg_array_47_39_real <= _zz_144;
      end
      if(_zz_50)begin
        img_reg_array_48_39_real <= _zz_144;
      end
      if(_zz_51)begin
        img_reg_array_49_39_real <= _zz_144;
      end
      if(_zz_52)begin
        img_reg_array_50_39_real <= _zz_144;
      end
      if(_zz_53)begin
        img_reg_array_51_39_real <= _zz_144;
      end
      if(_zz_54)begin
        img_reg_array_52_39_real <= _zz_144;
      end
      if(_zz_55)begin
        img_reg_array_53_39_real <= _zz_144;
      end
      if(_zz_56)begin
        img_reg_array_54_39_real <= _zz_144;
      end
      if(_zz_57)begin
        img_reg_array_55_39_real <= _zz_144;
      end
      if(_zz_58)begin
        img_reg_array_56_39_real <= _zz_144;
      end
      if(_zz_59)begin
        img_reg_array_57_39_real <= _zz_144;
      end
      if(_zz_60)begin
        img_reg_array_58_39_real <= _zz_144;
      end
      if(_zz_61)begin
        img_reg_array_59_39_real <= _zz_144;
      end
      if(_zz_62)begin
        img_reg_array_60_39_real <= _zz_144;
      end
      if(_zz_63)begin
        img_reg_array_61_39_real <= _zz_144;
      end
      if(_zz_64)begin
        img_reg_array_62_39_real <= _zz_144;
      end
      if(_zz_65)begin
        img_reg_array_63_39_real <= _zz_144;
      end
      if(_zz_2)begin
        img_reg_array_0_39_imag <= _zz_145;
      end
      if(_zz_3)begin
        img_reg_array_1_39_imag <= _zz_145;
      end
      if(_zz_4)begin
        img_reg_array_2_39_imag <= _zz_145;
      end
      if(_zz_5)begin
        img_reg_array_3_39_imag <= _zz_145;
      end
      if(_zz_6)begin
        img_reg_array_4_39_imag <= _zz_145;
      end
      if(_zz_7)begin
        img_reg_array_5_39_imag <= _zz_145;
      end
      if(_zz_8)begin
        img_reg_array_6_39_imag <= _zz_145;
      end
      if(_zz_9)begin
        img_reg_array_7_39_imag <= _zz_145;
      end
      if(_zz_10)begin
        img_reg_array_8_39_imag <= _zz_145;
      end
      if(_zz_11)begin
        img_reg_array_9_39_imag <= _zz_145;
      end
      if(_zz_12)begin
        img_reg_array_10_39_imag <= _zz_145;
      end
      if(_zz_13)begin
        img_reg_array_11_39_imag <= _zz_145;
      end
      if(_zz_14)begin
        img_reg_array_12_39_imag <= _zz_145;
      end
      if(_zz_15)begin
        img_reg_array_13_39_imag <= _zz_145;
      end
      if(_zz_16)begin
        img_reg_array_14_39_imag <= _zz_145;
      end
      if(_zz_17)begin
        img_reg_array_15_39_imag <= _zz_145;
      end
      if(_zz_18)begin
        img_reg_array_16_39_imag <= _zz_145;
      end
      if(_zz_19)begin
        img_reg_array_17_39_imag <= _zz_145;
      end
      if(_zz_20)begin
        img_reg_array_18_39_imag <= _zz_145;
      end
      if(_zz_21)begin
        img_reg_array_19_39_imag <= _zz_145;
      end
      if(_zz_22)begin
        img_reg_array_20_39_imag <= _zz_145;
      end
      if(_zz_23)begin
        img_reg_array_21_39_imag <= _zz_145;
      end
      if(_zz_24)begin
        img_reg_array_22_39_imag <= _zz_145;
      end
      if(_zz_25)begin
        img_reg_array_23_39_imag <= _zz_145;
      end
      if(_zz_26)begin
        img_reg_array_24_39_imag <= _zz_145;
      end
      if(_zz_27)begin
        img_reg_array_25_39_imag <= _zz_145;
      end
      if(_zz_28)begin
        img_reg_array_26_39_imag <= _zz_145;
      end
      if(_zz_29)begin
        img_reg_array_27_39_imag <= _zz_145;
      end
      if(_zz_30)begin
        img_reg_array_28_39_imag <= _zz_145;
      end
      if(_zz_31)begin
        img_reg_array_29_39_imag <= _zz_145;
      end
      if(_zz_32)begin
        img_reg_array_30_39_imag <= _zz_145;
      end
      if(_zz_33)begin
        img_reg_array_31_39_imag <= _zz_145;
      end
      if(_zz_34)begin
        img_reg_array_32_39_imag <= _zz_145;
      end
      if(_zz_35)begin
        img_reg_array_33_39_imag <= _zz_145;
      end
      if(_zz_36)begin
        img_reg_array_34_39_imag <= _zz_145;
      end
      if(_zz_37)begin
        img_reg_array_35_39_imag <= _zz_145;
      end
      if(_zz_38)begin
        img_reg_array_36_39_imag <= _zz_145;
      end
      if(_zz_39)begin
        img_reg_array_37_39_imag <= _zz_145;
      end
      if(_zz_40)begin
        img_reg_array_38_39_imag <= _zz_145;
      end
      if(_zz_41)begin
        img_reg_array_39_39_imag <= _zz_145;
      end
      if(_zz_42)begin
        img_reg_array_40_39_imag <= _zz_145;
      end
      if(_zz_43)begin
        img_reg_array_41_39_imag <= _zz_145;
      end
      if(_zz_44)begin
        img_reg_array_42_39_imag <= _zz_145;
      end
      if(_zz_45)begin
        img_reg_array_43_39_imag <= _zz_145;
      end
      if(_zz_46)begin
        img_reg_array_44_39_imag <= _zz_145;
      end
      if(_zz_47)begin
        img_reg_array_45_39_imag <= _zz_145;
      end
      if(_zz_48)begin
        img_reg_array_46_39_imag <= _zz_145;
      end
      if(_zz_49)begin
        img_reg_array_47_39_imag <= _zz_145;
      end
      if(_zz_50)begin
        img_reg_array_48_39_imag <= _zz_145;
      end
      if(_zz_51)begin
        img_reg_array_49_39_imag <= _zz_145;
      end
      if(_zz_52)begin
        img_reg_array_50_39_imag <= _zz_145;
      end
      if(_zz_53)begin
        img_reg_array_51_39_imag <= _zz_145;
      end
      if(_zz_54)begin
        img_reg_array_52_39_imag <= _zz_145;
      end
      if(_zz_55)begin
        img_reg_array_53_39_imag <= _zz_145;
      end
      if(_zz_56)begin
        img_reg_array_54_39_imag <= _zz_145;
      end
      if(_zz_57)begin
        img_reg_array_55_39_imag <= _zz_145;
      end
      if(_zz_58)begin
        img_reg_array_56_39_imag <= _zz_145;
      end
      if(_zz_59)begin
        img_reg_array_57_39_imag <= _zz_145;
      end
      if(_zz_60)begin
        img_reg_array_58_39_imag <= _zz_145;
      end
      if(_zz_61)begin
        img_reg_array_59_39_imag <= _zz_145;
      end
      if(_zz_62)begin
        img_reg_array_60_39_imag <= _zz_145;
      end
      if(_zz_63)begin
        img_reg_array_61_39_imag <= _zz_145;
      end
      if(_zz_64)begin
        img_reg_array_62_39_imag <= _zz_145;
      end
      if(_zz_65)begin
        img_reg_array_63_39_imag <= _zz_145;
      end
      if(_zz_2)begin
        img_reg_array_0_40_real <= _zz_146;
      end
      if(_zz_3)begin
        img_reg_array_1_40_real <= _zz_146;
      end
      if(_zz_4)begin
        img_reg_array_2_40_real <= _zz_146;
      end
      if(_zz_5)begin
        img_reg_array_3_40_real <= _zz_146;
      end
      if(_zz_6)begin
        img_reg_array_4_40_real <= _zz_146;
      end
      if(_zz_7)begin
        img_reg_array_5_40_real <= _zz_146;
      end
      if(_zz_8)begin
        img_reg_array_6_40_real <= _zz_146;
      end
      if(_zz_9)begin
        img_reg_array_7_40_real <= _zz_146;
      end
      if(_zz_10)begin
        img_reg_array_8_40_real <= _zz_146;
      end
      if(_zz_11)begin
        img_reg_array_9_40_real <= _zz_146;
      end
      if(_zz_12)begin
        img_reg_array_10_40_real <= _zz_146;
      end
      if(_zz_13)begin
        img_reg_array_11_40_real <= _zz_146;
      end
      if(_zz_14)begin
        img_reg_array_12_40_real <= _zz_146;
      end
      if(_zz_15)begin
        img_reg_array_13_40_real <= _zz_146;
      end
      if(_zz_16)begin
        img_reg_array_14_40_real <= _zz_146;
      end
      if(_zz_17)begin
        img_reg_array_15_40_real <= _zz_146;
      end
      if(_zz_18)begin
        img_reg_array_16_40_real <= _zz_146;
      end
      if(_zz_19)begin
        img_reg_array_17_40_real <= _zz_146;
      end
      if(_zz_20)begin
        img_reg_array_18_40_real <= _zz_146;
      end
      if(_zz_21)begin
        img_reg_array_19_40_real <= _zz_146;
      end
      if(_zz_22)begin
        img_reg_array_20_40_real <= _zz_146;
      end
      if(_zz_23)begin
        img_reg_array_21_40_real <= _zz_146;
      end
      if(_zz_24)begin
        img_reg_array_22_40_real <= _zz_146;
      end
      if(_zz_25)begin
        img_reg_array_23_40_real <= _zz_146;
      end
      if(_zz_26)begin
        img_reg_array_24_40_real <= _zz_146;
      end
      if(_zz_27)begin
        img_reg_array_25_40_real <= _zz_146;
      end
      if(_zz_28)begin
        img_reg_array_26_40_real <= _zz_146;
      end
      if(_zz_29)begin
        img_reg_array_27_40_real <= _zz_146;
      end
      if(_zz_30)begin
        img_reg_array_28_40_real <= _zz_146;
      end
      if(_zz_31)begin
        img_reg_array_29_40_real <= _zz_146;
      end
      if(_zz_32)begin
        img_reg_array_30_40_real <= _zz_146;
      end
      if(_zz_33)begin
        img_reg_array_31_40_real <= _zz_146;
      end
      if(_zz_34)begin
        img_reg_array_32_40_real <= _zz_146;
      end
      if(_zz_35)begin
        img_reg_array_33_40_real <= _zz_146;
      end
      if(_zz_36)begin
        img_reg_array_34_40_real <= _zz_146;
      end
      if(_zz_37)begin
        img_reg_array_35_40_real <= _zz_146;
      end
      if(_zz_38)begin
        img_reg_array_36_40_real <= _zz_146;
      end
      if(_zz_39)begin
        img_reg_array_37_40_real <= _zz_146;
      end
      if(_zz_40)begin
        img_reg_array_38_40_real <= _zz_146;
      end
      if(_zz_41)begin
        img_reg_array_39_40_real <= _zz_146;
      end
      if(_zz_42)begin
        img_reg_array_40_40_real <= _zz_146;
      end
      if(_zz_43)begin
        img_reg_array_41_40_real <= _zz_146;
      end
      if(_zz_44)begin
        img_reg_array_42_40_real <= _zz_146;
      end
      if(_zz_45)begin
        img_reg_array_43_40_real <= _zz_146;
      end
      if(_zz_46)begin
        img_reg_array_44_40_real <= _zz_146;
      end
      if(_zz_47)begin
        img_reg_array_45_40_real <= _zz_146;
      end
      if(_zz_48)begin
        img_reg_array_46_40_real <= _zz_146;
      end
      if(_zz_49)begin
        img_reg_array_47_40_real <= _zz_146;
      end
      if(_zz_50)begin
        img_reg_array_48_40_real <= _zz_146;
      end
      if(_zz_51)begin
        img_reg_array_49_40_real <= _zz_146;
      end
      if(_zz_52)begin
        img_reg_array_50_40_real <= _zz_146;
      end
      if(_zz_53)begin
        img_reg_array_51_40_real <= _zz_146;
      end
      if(_zz_54)begin
        img_reg_array_52_40_real <= _zz_146;
      end
      if(_zz_55)begin
        img_reg_array_53_40_real <= _zz_146;
      end
      if(_zz_56)begin
        img_reg_array_54_40_real <= _zz_146;
      end
      if(_zz_57)begin
        img_reg_array_55_40_real <= _zz_146;
      end
      if(_zz_58)begin
        img_reg_array_56_40_real <= _zz_146;
      end
      if(_zz_59)begin
        img_reg_array_57_40_real <= _zz_146;
      end
      if(_zz_60)begin
        img_reg_array_58_40_real <= _zz_146;
      end
      if(_zz_61)begin
        img_reg_array_59_40_real <= _zz_146;
      end
      if(_zz_62)begin
        img_reg_array_60_40_real <= _zz_146;
      end
      if(_zz_63)begin
        img_reg_array_61_40_real <= _zz_146;
      end
      if(_zz_64)begin
        img_reg_array_62_40_real <= _zz_146;
      end
      if(_zz_65)begin
        img_reg_array_63_40_real <= _zz_146;
      end
      if(_zz_2)begin
        img_reg_array_0_40_imag <= _zz_147;
      end
      if(_zz_3)begin
        img_reg_array_1_40_imag <= _zz_147;
      end
      if(_zz_4)begin
        img_reg_array_2_40_imag <= _zz_147;
      end
      if(_zz_5)begin
        img_reg_array_3_40_imag <= _zz_147;
      end
      if(_zz_6)begin
        img_reg_array_4_40_imag <= _zz_147;
      end
      if(_zz_7)begin
        img_reg_array_5_40_imag <= _zz_147;
      end
      if(_zz_8)begin
        img_reg_array_6_40_imag <= _zz_147;
      end
      if(_zz_9)begin
        img_reg_array_7_40_imag <= _zz_147;
      end
      if(_zz_10)begin
        img_reg_array_8_40_imag <= _zz_147;
      end
      if(_zz_11)begin
        img_reg_array_9_40_imag <= _zz_147;
      end
      if(_zz_12)begin
        img_reg_array_10_40_imag <= _zz_147;
      end
      if(_zz_13)begin
        img_reg_array_11_40_imag <= _zz_147;
      end
      if(_zz_14)begin
        img_reg_array_12_40_imag <= _zz_147;
      end
      if(_zz_15)begin
        img_reg_array_13_40_imag <= _zz_147;
      end
      if(_zz_16)begin
        img_reg_array_14_40_imag <= _zz_147;
      end
      if(_zz_17)begin
        img_reg_array_15_40_imag <= _zz_147;
      end
      if(_zz_18)begin
        img_reg_array_16_40_imag <= _zz_147;
      end
      if(_zz_19)begin
        img_reg_array_17_40_imag <= _zz_147;
      end
      if(_zz_20)begin
        img_reg_array_18_40_imag <= _zz_147;
      end
      if(_zz_21)begin
        img_reg_array_19_40_imag <= _zz_147;
      end
      if(_zz_22)begin
        img_reg_array_20_40_imag <= _zz_147;
      end
      if(_zz_23)begin
        img_reg_array_21_40_imag <= _zz_147;
      end
      if(_zz_24)begin
        img_reg_array_22_40_imag <= _zz_147;
      end
      if(_zz_25)begin
        img_reg_array_23_40_imag <= _zz_147;
      end
      if(_zz_26)begin
        img_reg_array_24_40_imag <= _zz_147;
      end
      if(_zz_27)begin
        img_reg_array_25_40_imag <= _zz_147;
      end
      if(_zz_28)begin
        img_reg_array_26_40_imag <= _zz_147;
      end
      if(_zz_29)begin
        img_reg_array_27_40_imag <= _zz_147;
      end
      if(_zz_30)begin
        img_reg_array_28_40_imag <= _zz_147;
      end
      if(_zz_31)begin
        img_reg_array_29_40_imag <= _zz_147;
      end
      if(_zz_32)begin
        img_reg_array_30_40_imag <= _zz_147;
      end
      if(_zz_33)begin
        img_reg_array_31_40_imag <= _zz_147;
      end
      if(_zz_34)begin
        img_reg_array_32_40_imag <= _zz_147;
      end
      if(_zz_35)begin
        img_reg_array_33_40_imag <= _zz_147;
      end
      if(_zz_36)begin
        img_reg_array_34_40_imag <= _zz_147;
      end
      if(_zz_37)begin
        img_reg_array_35_40_imag <= _zz_147;
      end
      if(_zz_38)begin
        img_reg_array_36_40_imag <= _zz_147;
      end
      if(_zz_39)begin
        img_reg_array_37_40_imag <= _zz_147;
      end
      if(_zz_40)begin
        img_reg_array_38_40_imag <= _zz_147;
      end
      if(_zz_41)begin
        img_reg_array_39_40_imag <= _zz_147;
      end
      if(_zz_42)begin
        img_reg_array_40_40_imag <= _zz_147;
      end
      if(_zz_43)begin
        img_reg_array_41_40_imag <= _zz_147;
      end
      if(_zz_44)begin
        img_reg_array_42_40_imag <= _zz_147;
      end
      if(_zz_45)begin
        img_reg_array_43_40_imag <= _zz_147;
      end
      if(_zz_46)begin
        img_reg_array_44_40_imag <= _zz_147;
      end
      if(_zz_47)begin
        img_reg_array_45_40_imag <= _zz_147;
      end
      if(_zz_48)begin
        img_reg_array_46_40_imag <= _zz_147;
      end
      if(_zz_49)begin
        img_reg_array_47_40_imag <= _zz_147;
      end
      if(_zz_50)begin
        img_reg_array_48_40_imag <= _zz_147;
      end
      if(_zz_51)begin
        img_reg_array_49_40_imag <= _zz_147;
      end
      if(_zz_52)begin
        img_reg_array_50_40_imag <= _zz_147;
      end
      if(_zz_53)begin
        img_reg_array_51_40_imag <= _zz_147;
      end
      if(_zz_54)begin
        img_reg_array_52_40_imag <= _zz_147;
      end
      if(_zz_55)begin
        img_reg_array_53_40_imag <= _zz_147;
      end
      if(_zz_56)begin
        img_reg_array_54_40_imag <= _zz_147;
      end
      if(_zz_57)begin
        img_reg_array_55_40_imag <= _zz_147;
      end
      if(_zz_58)begin
        img_reg_array_56_40_imag <= _zz_147;
      end
      if(_zz_59)begin
        img_reg_array_57_40_imag <= _zz_147;
      end
      if(_zz_60)begin
        img_reg_array_58_40_imag <= _zz_147;
      end
      if(_zz_61)begin
        img_reg_array_59_40_imag <= _zz_147;
      end
      if(_zz_62)begin
        img_reg_array_60_40_imag <= _zz_147;
      end
      if(_zz_63)begin
        img_reg_array_61_40_imag <= _zz_147;
      end
      if(_zz_64)begin
        img_reg_array_62_40_imag <= _zz_147;
      end
      if(_zz_65)begin
        img_reg_array_63_40_imag <= _zz_147;
      end
      if(_zz_2)begin
        img_reg_array_0_41_real <= _zz_148;
      end
      if(_zz_3)begin
        img_reg_array_1_41_real <= _zz_148;
      end
      if(_zz_4)begin
        img_reg_array_2_41_real <= _zz_148;
      end
      if(_zz_5)begin
        img_reg_array_3_41_real <= _zz_148;
      end
      if(_zz_6)begin
        img_reg_array_4_41_real <= _zz_148;
      end
      if(_zz_7)begin
        img_reg_array_5_41_real <= _zz_148;
      end
      if(_zz_8)begin
        img_reg_array_6_41_real <= _zz_148;
      end
      if(_zz_9)begin
        img_reg_array_7_41_real <= _zz_148;
      end
      if(_zz_10)begin
        img_reg_array_8_41_real <= _zz_148;
      end
      if(_zz_11)begin
        img_reg_array_9_41_real <= _zz_148;
      end
      if(_zz_12)begin
        img_reg_array_10_41_real <= _zz_148;
      end
      if(_zz_13)begin
        img_reg_array_11_41_real <= _zz_148;
      end
      if(_zz_14)begin
        img_reg_array_12_41_real <= _zz_148;
      end
      if(_zz_15)begin
        img_reg_array_13_41_real <= _zz_148;
      end
      if(_zz_16)begin
        img_reg_array_14_41_real <= _zz_148;
      end
      if(_zz_17)begin
        img_reg_array_15_41_real <= _zz_148;
      end
      if(_zz_18)begin
        img_reg_array_16_41_real <= _zz_148;
      end
      if(_zz_19)begin
        img_reg_array_17_41_real <= _zz_148;
      end
      if(_zz_20)begin
        img_reg_array_18_41_real <= _zz_148;
      end
      if(_zz_21)begin
        img_reg_array_19_41_real <= _zz_148;
      end
      if(_zz_22)begin
        img_reg_array_20_41_real <= _zz_148;
      end
      if(_zz_23)begin
        img_reg_array_21_41_real <= _zz_148;
      end
      if(_zz_24)begin
        img_reg_array_22_41_real <= _zz_148;
      end
      if(_zz_25)begin
        img_reg_array_23_41_real <= _zz_148;
      end
      if(_zz_26)begin
        img_reg_array_24_41_real <= _zz_148;
      end
      if(_zz_27)begin
        img_reg_array_25_41_real <= _zz_148;
      end
      if(_zz_28)begin
        img_reg_array_26_41_real <= _zz_148;
      end
      if(_zz_29)begin
        img_reg_array_27_41_real <= _zz_148;
      end
      if(_zz_30)begin
        img_reg_array_28_41_real <= _zz_148;
      end
      if(_zz_31)begin
        img_reg_array_29_41_real <= _zz_148;
      end
      if(_zz_32)begin
        img_reg_array_30_41_real <= _zz_148;
      end
      if(_zz_33)begin
        img_reg_array_31_41_real <= _zz_148;
      end
      if(_zz_34)begin
        img_reg_array_32_41_real <= _zz_148;
      end
      if(_zz_35)begin
        img_reg_array_33_41_real <= _zz_148;
      end
      if(_zz_36)begin
        img_reg_array_34_41_real <= _zz_148;
      end
      if(_zz_37)begin
        img_reg_array_35_41_real <= _zz_148;
      end
      if(_zz_38)begin
        img_reg_array_36_41_real <= _zz_148;
      end
      if(_zz_39)begin
        img_reg_array_37_41_real <= _zz_148;
      end
      if(_zz_40)begin
        img_reg_array_38_41_real <= _zz_148;
      end
      if(_zz_41)begin
        img_reg_array_39_41_real <= _zz_148;
      end
      if(_zz_42)begin
        img_reg_array_40_41_real <= _zz_148;
      end
      if(_zz_43)begin
        img_reg_array_41_41_real <= _zz_148;
      end
      if(_zz_44)begin
        img_reg_array_42_41_real <= _zz_148;
      end
      if(_zz_45)begin
        img_reg_array_43_41_real <= _zz_148;
      end
      if(_zz_46)begin
        img_reg_array_44_41_real <= _zz_148;
      end
      if(_zz_47)begin
        img_reg_array_45_41_real <= _zz_148;
      end
      if(_zz_48)begin
        img_reg_array_46_41_real <= _zz_148;
      end
      if(_zz_49)begin
        img_reg_array_47_41_real <= _zz_148;
      end
      if(_zz_50)begin
        img_reg_array_48_41_real <= _zz_148;
      end
      if(_zz_51)begin
        img_reg_array_49_41_real <= _zz_148;
      end
      if(_zz_52)begin
        img_reg_array_50_41_real <= _zz_148;
      end
      if(_zz_53)begin
        img_reg_array_51_41_real <= _zz_148;
      end
      if(_zz_54)begin
        img_reg_array_52_41_real <= _zz_148;
      end
      if(_zz_55)begin
        img_reg_array_53_41_real <= _zz_148;
      end
      if(_zz_56)begin
        img_reg_array_54_41_real <= _zz_148;
      end
      if(_zz_57)begin
        img_reg_array_55_41_real <= _zz_148;
      end
      if(_zz_58)begin
        img_reg_array_56_41_real <= _zz_148;
      end
      if(_zz_59)begin
        img_reg_array_57_41_real <= _zz_148;
      end
      if(_zz_60)begin
        img_reg_array_58_41_real <= _zz_148;
      end
      if(_zz_61)begin
        img_reg_array_59_41_real <= _zz_148;
      end
      if(_zz_62)begin
        img_reg_array_60_41_real <= _zz_148;
      end
      if(_zz_63)begin
        img_reg_array_61_41_real <= _zz_148;
      end
      if(_zz_64)begin
        img_reg_array_62_41_real <= _zz_148;
      end
      if(_zz_65)begin
        img_reg_array_63_41_real <= _zz_148;
      end
      if(_zz_2)begin
        img_reg_array_0_41_imag <= _zz_149;
      end
      if(_zz_3)begin
        img_reg_array_1_41_imag <= _zz_149;
      end
      if(_zz_4)begin
        img_reg_array_2_41_imag <= _zz_149;
      end
      if(_zz_5)begin
        img_reg_array_3_41_imag <= _zz_149;
      end
      if(_zz_6)begin
        img_reg_array_4_41_imag <= _zz_149;
      end
      if(_zz_7)begin
        img_reg_array_5_41_imag <= _zz_149;
      end
      if(_zz_8)begin
        img_reg_array_6_41_imag <= _zz_149;
      end
      if(_zz_9)begin
        img_reg_array_7_41_imag <= _zz_149;
      end
      if(_zz_10)begin
        img_reg_array_8_41_imag <= _zz_149;
      end
      if(_zz_11)begin
        img_reg_array_9_41_imag <= _zz_149;
      end
      if(_zz_12)begin
        img_reg_array_10_41_imag <= _zz_149;
      end
      if(_zz_13)begin
        img_reg_array_11_41_imag <= _zz_149;
      end
      if(_zz_14)begin
        img_reg_array_12_41_imag <= _zz_149;
      end
      if(_zz_15)begin
        img_reg_array_13_41_imag <= _zz_149;
      end
      if(_zz_16)begin
        img_reg_array_14_41_imag <= _zz_149;
      end
      if(_zz_17)begin
        img_reg_array_15_41_imag <= _zz_149;
      end
      if(_zz_18)begin
        img_reg_array_16_41_imag <= _zz_149;
      end
      if(_zz_19)begin
        img_reg_array_17_41_imag <= _zz_149;
      end
      if(_zz_20)begin
        img_reg_array_18_41_imag <= _zz_149;
      end
      if(_zz_21)begin
        img_reg_array_19_41_imag <= _zz_149;
      end
      if(_zz_22)begin
        img_reg_array_20_41_imag <= _zz_149;
      end
      if(_zz_23)begin
        img_reg_array_21_41_imag <= _zz_149;
      end
      if(_zz_24)begin
        img_reg_array_22_41_imag <= _zz_149;
      end
      if(_zz_25)begin
        img_reg_array_23_41_imag <= _zz_149;
      end
      if(_zz_26)begin
        img_reg_array_24_41_imag <= _zz_149;
      end
      if(_zz_27)begin
        img_reg_array_25_41_imag <= _zz_149;
      end
      if(_zz_28)begin
        img_reg_array_26_41_imag <= _zz_149;
      end
      if(_zz_29)begin
        img_reg_array_27_41_imag <= _zz_149;
      end
      if(_zz_30)begin
        img_reg_array_28_41_imag <= _zz_149;
      end
      if(_zz_31)begin
        img_reg_array_29_41_imag <= _zz_149;
      end
      if(_zz_32)begin
        img_reg_array_30_41_imag <= _zz_149;
      end
      if(_zz_33)begin
        img_reg_array_31_41_imag <= _zz_149;
      end
      if(_zz_34)begin
        img_reg_array_32_41_imag <= _zz_149;
      end
      if(_zz_35)begin
        img_reg_array_33_41_imag <= _zz_149;
      end
      if(_zz_36)begin
        img_reg_array_34_41_imag <= _zz_149;
      end
      if(_zz_37)begin
        img_reg_array_35_41_imag <= _zz_149;
      end
      if(_zz_38)begin
        img_reg_array_36_41_imag <= _zz_149;
      end
      if(_zz_39)begin
        img_reg_array_37_41_imag <= _zz_149;
      end
      if(_zz_40)begin
        img_reg_array_38_41_imag <= _zz_149;
      end
      if(_zz_41)begin
        img_reg_array_39_41_imag <= _zz_149;
      end
      if(_zz_42)begin
        img_reg_array_40_41_imag <= _zz_149;
      end
      if(_zz_43)begin
        img_reg_array_41_41_imag <= _zz_149;
      end
      if(_zz_44)begin
        img_reg_array_42_41_imag <= _zz_149;
      end
      if(_zz_45)begin
        img_reg_array_43_41_imag <= _zz_149;
      end
      if(_zz_46)begin
        img_reg_array_44_41_imag <= _zz_149;
      end
      if(_zz_47)begin
        img_reg_array_45_41_imag <= _zz_149;
      end
      if(_zz_48)begin
        img_reg_array_46_41_imag <= _zz_149;
      end
      if(_zz_49)begin
        img_reg_array_47_41_imag <= _zz_149;
      end
      if(_zz_50)begin
        img_reg_array_48_41_imag <= _zz_149;
      end
      if(_zz_51)begin
        img_reg_array_49_41_imag <= _zz_149;
      end
      if(_zz_52)begin
        img_reg_array_50_41_imag <= _zz_149;
      end
      if(_zz_53)begin
        img_reg_array_51_41_imag <= _zz_149;
      end
      if(_zz_54)begin
        img_reg_array_52_41_imag <= _zz_149;
      end
      if(_zz_55)begin
        img_reg_array_53_41_imag <= _zz_149;
      end
      if(_zz_56)begin
        img_reg_array_54_41_imag <= _zz_149;
      end
      if(_zz_57)begin
        img_reg_array_55_41_imag <= _zz_149;
      end
      if(_zz_58)begin
        img_reg_array_56_41_imag <= _zz_149;
      end
      if(_zz_59)begin
        img_reg_array_57_41_imag <= _zz_149;
      end
      if(_zz_60)begin
        img_reg_array_58_41_imag <= _zz_149;
      end
      if(_zz_61)begin
        img_reg_array_59_41_imag <= _zz_149;
      end
      if(_zz_62)begin
        img_reg_array_60_41_imag <= _zz_149;
      end
      if(_zz_63)begin
        img_reg_array_61_41_imag <= _zz_149;
      end
      if(_zz_64)begin
        img_reg_array_62_41_imag <= _zz_149;
      end
      if(_zz_65)begin
        img_reg_array_63_41_imag <= _zz_149;
      end
      if(_zz_2)begin
        img_reg_array_0_42_real <= _zz_150;
      end
      if(_zz_3)begin
        img_reg_array_1_42_real <= _zz_150;
      end
      if(_zz_4)begin
        img_reg_array_2_42_real <= _zz_150;
      end
      if(_zz_5)begin
        img_reg_array_3_42_real <= _zz_150;
      end
      if(_zz_6)begin
        img_reg_array_4_42_real <= _zz_150;
      end
      if(_zz_7)begin
        img_reg_array_5_42_real <= _zz_150;
      end
      if(_zz_8)begin
        img_reg_array_6_42_real <= _zz_150;
      end
      if(_zz_9)begin
        img_reg_array_7_42_real <= _zz_150;
      end
      if(_zz_10)begin
        img_reg_array_8_42_real <= _zz_150;
      end
      if(_zz_11)begin
        img_reg_array_9_42_real <= _zz_150;
      end
      if(_zz_12)begin
        img_reg_array_10_42_real <= _zz_150;
      end
      if(_zz_13)begin
        img_reg_array_11_42_real <= _zz_150;
      end
      if(_zz_14)begin
        img_reg_array_12_42_real <= _zz_150;
      end
      if(_zz_15)begin
        img_reg_array_13_42_real <= _zz_150;
      end
      if(_zz_16)begin
        img_reg_array_14_42_real <= _zz_150;
      end
      if(_zz_17)begin
        img_reg_array_15_42_real <= _zz_150;
      end
      if(_zz_18)begin
        img_reg_array_16_42_real <= _zz_150;
      end
      if(_zz_19)begin
        img_reg_array_17_42_real <= _zz_150;
      end
      if(_zz_20)begin
        img_reg_array_18_42_real <= _zz_150;
      end
      if(_zz_21)begin
        img_reg_array_19_42_real <= _zz_150;
      end
      if(_zz_22)begin
        img_reg_array_20_42_real <= _zz_150;
      end
      if(_zz_23)begin
        img_reg_array_21_42_real <= _zz_150;
      end
      if(_zz_24)begin
        img_reg_array_22_42_real <= _zz_150;
      end
      if(_zz_25)begin
        img_reg_array_23_42_real <= _zz_150;
      end
      if(_zz_26)begin
        img_reg_array_24_42_real <= _zz_150;
      end
      if(_zz_27)begin
        img_reg_array_25_42_real <= _zz_150;
      end
      if(_zz_28)begin
        img_reg_array_26_42_real <= _zz_150;
      end
      if(_zz_29)begin
        img_reg_array_27_42_real <= _zz_150;
      end
      if(_zz_30)begin
        img_reg_array_28_42_real <= _zz_150;
      end
      if(_zz_31)begin
        img_reg_array_29_42_real <= _zz_150;
      end
      if(_zz_32)begin
        img_reg_array_30_42_real <= _zz_150;
      end
      if(_zz_33)begin
        img_reg_array_31_42_real <= _zz_150;
      end
      if(_zz_34)begin
        img_reg_array_32_42_real <= _zz_150;
      end
      if(_zz_35)begin
        img_reg_array_33_42_real <= _zz_150;
      end
      if(_zz_36)begin
        img_reg_array_34_42_real <= _zz_150;
      end
      if(_zz_37)begin
        img_reg_array_35_42_real <= _zz_150;
      end
      if(_zz_38)begin
        img_reg_array_36_42_real <= _zz_150;
      end
      if(_zz_39)begin
        img_reg_array_37_42_real <= _zz_150;
      end
      if(_zz_40)begin
        img_reg_array_38_42_real <= _zz_150;
      end
      if(_zz_41)begin
        img_reg_array_39_42_real <= _zz_150;
      end
      if(_zz_42)begin
        img_reg_array_40_42_real <= _zz_150;
      end
      if(_zz_43)begin
        img_reg_array_41_42_real <= _zz_150;
      end
      if(_zz_44)begin
        img_reg_array_42_42_real <= _zz_150;
      end
      if(_zz_45)begin
        img_reg_array_43_42_real <= _zz_150;
      end
      if(_zz_46)begin
        img_reg_array_44_42_real <= _zz_150;
      end
      if(_zz_47)begin
        img_reg_array_45_42_real <= _zz_150;
      end
      if(_zz_48)begin
        img_reg_array_46_42_real <= _zz_150;
      end
      if(_zz_49)begin
        img_reg_array_47_42_real <= _zz_150;
      end
      if(_zz_50)begin
        img_reg_array_48_42_real <= _zz_150;
      end
      if(_zz_51)begin
        img_reg_array_49_42_real <= _zz_150;
      end
      if(_zz_52)begin
        img_reg_array_50_42_real <= _zz_150;
      end
      if(_zz_53)begin
        img_reg_array_51_42_real <= _zz_150;
      end
      if(_zz_54)begin
        img_reg_array_52_42_real <= _zz_150;
      end
      if(_zz_55)begin
        img_reg_array_53_42_real <= _zz_150;
      end
      if(_zz_56)begin
        img_reg_array_54_42_real <= _zz_150;
      end
      if(_zz_57)begin
        img_reg_array_55_42_real <= _zz_150;
      end
      if(_zz_58)begin
        img_reg_array_56_42_real <= _zz_150;
      end
      if(_zz_59)begin
        img_reg_array_57_42_real <= _zz_150;
      end
      if(_zz_60)begin
        img_reg_array_58_42_real <= _zz_150;
      end
      if(_zz_61)begin
        img_reg_array_59_42_real <= _zz_150;
      end
      if(_zz_62)begin
        img_reg_array_60_42_real <= _zz_150;
      end
      if(_zz_63)begin
        img_reg_array_61_42_real <= _zz_150;
      end
      if(_zz_64)begin
        img_reg_array_62_42_real <= _zz_150;
      end
      if(_zz_65)begin
        img_reg_array_63_42_real <= _zz_150;
      end
      if(_zz_2)begin
        img_reg_array_0_42_imag <= _zz_151;
      end
      if(_zz_3)begin
        img_reg_array_1_42_imag <= _zz_151;
      end
      if(_zz_4)begin
        img_reg_array_2_42_imag <= _zz_151;
      end
      if(_zz_5)begin
        img_reg_array_3_42_imag <= _zz_151;
      end
      if(_zz_6)begin
        img_reg_array_4_42_imag <= _zz_151;
      end
      if(_zz_7)begin
        img_reg_array_5_42_imag <= _zz_151;
      end
      if(_zz_8)begin
        img_reg_array_6_42_imag <= _zz_151;
      end
      if(_zz_9)begin
        img_reg_array_7_42_imag <= _zz_151;
      end
      if(_zz_10)begin
        img_reg_array_8_42_imag <= _zz_151;
      end
      if(_zz_11)begin
        img_reg_array_9_42_imag <= _zz_151;
      end
      if(_zz_12)begin
        img_reg_array_10_42_imag <= _zz_151;
      end
      if(_zz_13)begin
        img_reg_array_11_42_imag <= _zz_151;
      end
      if(_zz_14)begin
        img_reg_array_12_42_imag <= _zz_151;
      end
      if(_zz_15)begin
        img_reg_array_13_42_imag <= _zz_151;
      end
      if(_zz_16)begin
        img_reg_array_14_42_imag <= _zz_151;
      end
      if(_zz_17)begin
        img_reg_array_15_42_imag <= _zz_151;
      end
      if(_zz_18)begin
        img_reg_array_16_42_imag <= _zz_151;
      end
      if(_zz_19)begin
        img_reg_array_17_42_imag <= _zz_151;
      end
      if(_zz_20)begin
        img_reg_array_18_42_imag <= _zz_151;
      end
      if(_zz_21)begin
        img_reg_array_19_42_imag <= _zz_151;
      end
      if(_zz_22)begin
        img_reg_array_20_42_imag <= _zz_151;
      end
      if(_zz_23)begin
        img_reg_array_21_42_imag <= _zz_151;
      end
      if(_zz_24)begin
        img_reg_array_22_42_imag <= _zz_151;
      end
      if(_zz_25)begin
        img_reg_array_23_42_imag <= _zz_151;
      end
      if(_zz_26)begin
        img_reg_array_24_42_imag <= _zz_151;
      end
      if(_zz_27)begin
        img_reg_array_25_42_imag <= _zz_151;
      end
      if(_zz_28)begin
        img_reg_array_26_42_imag <= _zz_151;
      end
      if(_zz_29)begin
        img_reg_array_27_42_imag <= _zz_151;
      end
      if(_zz_30)begin
        img_reg_array_28_42_imag <= _zz_151;
      end
      if(_zz_31)begin
        img_reg_array_29_42_imag <= _zz_151;
      end
      if(_zz_32)begin
        img_reg_array_30_42_imag <= _zz_151;
      end
      if(_zz_33)begin
        img_reg_array_31_42_imag <= _zz_151;
      end
      if(_zz_34)begin
        img_reg_array_32_42_imag <= _zz_151;
      end
      if(_zz_35)begin
        img_reg_array_33_42_imag <= _zz_151;
      end
      if(_zz_36)begin
        img_reg_array_34_42_imag <= _zz_151;
      end
      if(_zz_37)begin
        img_reg_array_35_42_imag <= _zz_151;
      end
      if(_zz_38)begin
        img_reg_array_36_42_imag <= _zz_151;
      end
      if(_zz_39)begin
        img_reg_array_37_42_imag <= _zz_151;
      end
      if(_zz_40)begin
        img_reg_array_38_42_imag <= _zz_151;
      end
      if(_zz_41)begin
        img_reg_array_39_42_imag <= _zz_151;
      end
      if(_zz_42)begin
        img_reg_array_40_42_imag <= _zz_151;
      end
      if(_zz_43)begin
        img_reg_array_41_42_imag <= _zz_151;
      end
      if(_zz_44)begin
        img_reg_array_42_42_imag <= _zz_151;
      end
      if(_zz_45)begin
        img_reg_array_43_42_imag <= _zz_151;
      end
      if(_zz_46)begin
        img_reg_array_44_42_imag <= _zz_151;
      end
      if(_zz_47)begin
        img_reg_array_45_42_imag <= _zz_151;
      end
      if(_zz_48)begin
        img_reg_array_46_42_imag <= _zz_151;
      end
      if(_zz_49)begin
        img_reg_array_47_42_imag <= _zz_151;
      end
      if(_zz_50)begin
        img_reg_array_48_42_imag <= _zz_151;
      end
      if(_zz_51)begin
        img_reg_array_49_42_imag <= _zz_151;
      end
      if(_zz_52)begin
        img_reg_array_50_42_imag <= _zz_151;
      end
      if(_zz_53)begin
        img_reg_array_51_42_imag <= _zz_151;
      end
      if(_zz_54)begin
        img_reg_array_52_42_imag <= _zz_151;
      end
      if(_zz_55)begin
        img_reg_array_53_42_imag <= _zz_151;
      end
      if(_zz_56)begin
        img_reg_array_54_42_imag <= _zz_151;
      end
      if(_zz_57)begin
        img_reg_array_55_42_imag <= _zz_151;
      end
      if(_zz_58)begin
        img_reg_array_56_42_imag <= _zz_151;
      end
      if(_zz_59)begin
        img_reg_array_57_42_imag <= _zz_151;
      end
      if(_zz_60)begin
        img_reg_array_58_42_imag <= _zz_151;
      end
      if(_zz_61)begin
        img_reg_array_59_42_imag <= _zz_151;
      end
      if(_zz_62)begin
        img_reg_array_60_42_imag <= _zz_151;
      end
      if(_zz_63)begin
        img_reg_array_61_42_imag <= _zz_151;
      end
      if(_zz_64)begin
        img_reg_array_62_42_imag <= _zz_151;
      end
      if(_zz_65)begin
        img_reg_array_63_42_imag <= _zz_151;
      end
      if(_zz_2)begin
        img_reg_array_0_43_real <= _zz_152;
      end
      if(_zz_3)begin
        img_reg_array_1_43_real <= _zz_152;
      end
      if(_zz_4)begin
        img_reg_array_2_43_real <= _zz_152;
      end
      if(_zz_5)begin
        img_reg_array_3_43_real <= _zz_152;
      end
      if(_zz_6)begin
        img_reg_array_4_43_real <= _zz_152;
      end
      if(_zz_7)begin
        img_reg_array_5_43_real <= _zz_152;
      end
      if(_zz_8)begin
        img_reg_array_6_43_real <= _zz_152;
      end
      if(_zz_9)begin
        img_reg_array_7_43_real <= _zz_152;
      end
      if(_zz_10)begin
        img_reg_array_8_43_real <= _zz_152;
      end
      if(_zz_11)begin
        img_reg_array_9_43_real <= _zz_152;
      end
      if(_zz_12)begin
        img_reg_array_10_43_real <= _zz_152;
      end
      if(_zz_13)begin
        img_reg_array_11_43_real <= _zz_152;
      end
      if(_zz_14)begin
        img_reg_array_12_43_real <= _zz_152;
      end
      if(_zz_15)begin
        img_reg_array_13_43_real <= _zz_152;
      end
      if(_zz_16)begin
        img_reg_array_14_43_real <= _zz_152;
      end
      if(_zz_17)begin
        img_reg_array_15_43_real <= _zz_152;
      end
      if(_zz_18)begin
        img_reg_array_16_43_real <= _zz_152;
      end
      if(_zz_19)begin
        img_reg_array_17_43_real <= _zz_152;
      end
      if(_zz_20)begin
        img_reg_array_18_43_real <= _zz_152;
      end
      if(_zz_21)begin
        img_reg_array_19_43_real <= _zz_152;
      end
      if(_zz_22)begin
        img_reg_array_20_43_real <= _zz_152;
      end
      if(_zz_23)begin
        img_reg_array_21_43_real <= _zz_152;
      end
      if(_zz_24)begin
        img_reg_array_22_43_real <= _zz_152;
      end
      if(_zz_25)begin
        img_reg_array_23_43_real <= _zz_152;
      end
      if(_zz_26)begin
        img_reg_array_24_43_real <= _zz_152;
      end
      if(_zz_27)begin
        img_reg_array_25_43_real <= _zz_152;
      end
      if(_zz_28)begin
        img_reg_array_26_43_real <= _zz_152;
      end
      if(_zz_29)begin
        img_reg_array_27_43_real <= _zz_152;
      end
      if(_zz_30)begin
        img_reg_array_28_43_real <= _zz_152;
      end
      if(_zz_31)begin
        img_reg_array_29_43_real <= _zz_152;
      end
      if(_zz_32)begin
        img_reg_array_30_43_real <= _zz_152;
      end
      if(_zz_33)begin
        img_reg_array_31_43_real <= _zz_152;
      end
      if(_zz_34)begin
        img_reg_array_32_43_real <= _zz_152;
      end
      if(_zz_35)begin
        img_reg_array_33_43_real <= _zz_152;
      end
      if(_zz_36)begin
        img_reg_array_34_43_real <= _zz_152;
      end
      if(_zz_37)begin
        img_reg_array_35_43_real <= _zz_152;
      end
      if(_zz_38)begin
        img_reg_array_36_43_real <= _zz_152;
      end
      if(_zz_39)begin
        img_reg_array_37_43_real <= _zz_152;
      end
      if(_zz_40)begin
        img_reg_array_38_43_real <= _zz_152;
      end
      if(_zz_41)begin
        img_reg_array_39_43_real <= _zz_152;
      end
      if(_zz_42)begin
        img_reg_array_40_43_real <= _zz_152;
      end
      if(_zz_43)begin
        img_reg_array_41_43_real <= _zz_152;
      end
      if(_zz_44)begin
        img_reg_array_42_43_real <= _zz_152;
      end
      if(_zz_45)begin
        img_reg_array_43_43_real <= _zz_152;
      end
      if(_zz_46)begin
        img_reg_array_44_43_real <= _zz_152;
      end
      if(_zz_47)begin
        img_reg_array_45_43_real <= _zz_152;
      end
      if(_zz_48)begin
        img_reg_array_46_43_real <= _zz_152;
      end
      if(_zz_49)begin
        img_reg_array_47_43_real <= _zz_152;
      end
      if(_zz_50)begin
        img_reg_array_48_43_real <= _zz_152;
      end
      if(_zz_51)begin
        img_reg_array_49_43_real <= _zz_152;
      end
      if(_zz_52)begin
        img_reg_array_50_43_real <= _zz_152;
      end
      if(_zz_53)begin
        img_reg_array_51_43_real <= _zz_152;
      end
      if(_zz_54)begin
        img_reg_array_52_43_real <= _zz_152;
      end
      if(_zz_55)begin
        img_reg_array_53_43_real <= _zz_152;
      end
      if(_zz_56)begin
        img_reg_array_54_43_real <= _zz_152;
      end
      if(_zz_57)begin
        img_reg_array_55_43_real <= _zz_152;
      end
      if(_zz_58)begin
        img_reg_array_56_43_real <= _zz_152;
      end
      if(_zz_59)begin
        img_reg_array_57_43_real <= _zz_152;
      end
      if(_zz_60)begin
        img_reg_array_58_43_real <= _zz_152;
      end
      if(_zz_61)begin
        img_reg_array_59_43_real <= _zz_152;
      end
      if(_zz_62)begin
        img_reg_array_60_43_real <= _zz_152;
      end
      if(_zz_63)begin
        img_reg_array_61_43_real <= _zz_152;
      end
      if(_zz_64)begin
        img_reg_array_62_43_real <= _zz_152;
      end
      if(_zz_65)begin
        img_reg_array_63_43_real <= _zz_152;
      end
      if(_zz_2)begin
        img_reg_array_0_43_imag <= _zz_153;
      end
      if(_zz_3)begin
        img_reg_array_1_43_imag <= _zz_153;
      end
      if(_zz_4)begin
        img_reg_array_2_43_imag <= _zz_153;
      end
      if(_zz_5)begin
        img_reg_array_3_43_imag <= _zz_153;
      end
      if(_zz_6)begin
        img_reg_array_4_43_imag <= _zz_153;
      end
      if(_zz_7)begin
        img_reg_array_5_43_imag <= _zz_153;
      end
      if(_zz_8)begin
        img_reg_array_6_43_imag <= _zz_153;
      end
      if(_zz_9)begin
        img_reg_array_7_43_imag <= _zz_153;
      end
      if(_zz_10)begin
        img_reg_array_8_43_imag <= _zz_153;
      end
      if(_zz_11)begin
        img_reg_array_9_43_imag <= _zz_153;
      end
      if(_zz_12)begin
        img_reg_array_10_43_imag <= _zz_153;
      end
      if(_zz_13)begin
        img_reg_array_11_43_imag <= _zz_153;
      end
      if(_zz_14)begin
        img_reg_array_12_43_imag <= _zz_153;
      end
      if(_zz_15)begin
        img_reg_array_13_43_imag <= _zz_153;
      end
      if(_zz_16)begin
        img_reg_array_14_43_imag <= _zz_153;
      end
      if(_zz_17)begin
        img_reg_array_15_43_imag <= _zz_153;
      end
      if(_zz_18)begin
        img_reg_array_16_43_imag <= _zz_153;
      end
      if(_zz_19)begin
        img_reg_array_17_43_imag <= _zz_153;
      end
      if(_zz_20)begin
        img_reg_array_18_43_imag <= _zz_153;
      end
      if(_zz_21)begin
        img_reg_array_19_43_imag <= _zz_153;
      end
      if(_zz_22)begin
        img_reg_array_20_43_imag <= _zz_153;
      end
      if(_zz_23)begin
        img_reg_array_21_43_imag <= _zz_153;
      end
      if(_zz_24)begin
        img_reg_array_22_43_imag <= _zz_153;
      end
      if(_zz_25)begin
        img_reg_array_23_43_imag <= _zz_153;
      end
      if(_zz_26)begin
        img_reg_array_24_43_imag <= _zz_153;
      end
      if(_zz_27)begin
        img_reg_array_25_43_imag <= _zz_153;
      end
      if(_zz_28)begin
        img_reg_array_26_43_imag <= _zz_153;
      end
      if(_zz_29)begin
        img_reg_array_27_43_imag <= _zz_153;
      end
      if(_zz_30)begin
        img_reg_array_28_43_imag <= _zz_153;
      end
      if(_zz_31)begin
        img_reg_array_29_43_imag <= _zz_153;
      end
      if(_zz_32)begin
        img_reg_array_30_43_imag <= _zz_153;
      end
      if(_zz_33)begin
        img_reg_array_31_43_imag <= _zz_153;
      end
      if(_zz_34)begin
        img_reg_array_32_43_imag <= _zz_153;
      end
      if(_zz_35)begin
        img_reg_array_33_43_imag <= _zz_153;
      end
      if(_zz_36)begin
        img_reg_array_34_43_imag <= _zz_153;
      end
      if(_zz_37)begin
        img_reg_array_35_43_imag <= _zz_153;
      end
      if(_zz_38)begin
        img_reg_array_36_43_imag <= _zz_153;
      end
      if(_zz_39)begin
        img_reg_array_37_43_imag <= _zz_153;
      end
      if(_zz_40)begin
        img_reg_array_38_43_imag <= _zz_153;
      end
      if(_zz_41)begin
        img_reg_array_39_43_imag <= _zz_153;
      end
      if(_zz_42)begin
        img_reg_array_40_43_imag <= _zz_153;
      end
      if(_zz_43)begin
        img_reg_array_41_43_imag <= _zz_153;
      end
      if(_zz_44)begin
        img_reg_array_42_43_imag <= _zz_153;
      end
      if(_zz_45)begin
        img_reg_array_43_43_imag <= _zz_153;
      end
      if(_zz_46)begin
        img_reg_array_44_43_imag <= _zz_153;
      end
      if(_zz_47)begin
        img_reg_array_45_43_imag <= _zz_153;
      end
      if(_zz_48)begin
        img_reg_array_46_43_imag <= _zz_153;
      end
      if(_zz_49)begin
        img_reg_array_47_43_imag <= _zz_153;
      end
      if(_zz_50)begin
        img_reg_array_48_43_imag <= _zz_153;
      end
      if(_zz_51)begin
        img_reg_array_49_43_imag <= _zz_153;
      end
      if(_zz_52)begin
        img_reg_array_50_43_imag <= _zz_153;
      end
      if(_zz_53)begin
        img_reg_array_51_43_imag <= _zz_153;
      end
      if(_zz_54)begin
        img_reg_array_52_43_imag <= _zz_153;
      end
      if(_zz_55)begin
        img_reg_array_53_43_imag <= _zz_153;
      end
      if(_zz_56)begin
        img_reg_array_54_43_imag <= _zz_153;
      end
      if(_zz_57)begin
        img_reg_array_55_43_imag <= _zz_153;
      end
      if(_zz_58)begin
        img_reg_array_56_43_imag <= _zz_153;
      end
      if(_zz_59)begin
        img_reg_array_57_43_imag <= _zz_153;
      end
      if(_zz_60)begin
        img_reg_array_58_43_imag <= _zz_153;
      end
      if(_zz_61)begin
        img_reg_array_59_43_imag <= _zz_153;
      end
      if(_zz_62)begin
        img_reg_array_60_43_imag <= _zz_153;
      end
      if(_zz_63)begin
        img_reg_array_61_43_imag <= _zz_153;
      end
      if(_zz_64)begin
        img_reg_array_62_43_imag <= _zz_153;
      end
      if(_zz_65)begin
        img_reg_array_63_43_imag <= _zz_153;
      end
      if(_zz_2)begin
        img_reg_array_0_44_real <= _zz_154;
      end
      if(_zz_3)begin
        img_reg_array_1_44_real <= _zz_154;
      end
      if(_zz_4)begin
        img_reg_array_2_44_real <= _zz_154;
      end
      if(_zz_5)begin
        img_reg_array_3_44_real <= _zz_154;
      end
      if(_zz_6)begin
        img_reg_array_4_44_real <= _zz_154;
      end
      if(_zz_7)begin
        img_reg_array_5_44_real <= _zz_154;
      end
      if(_zz_8)begin
        img_reg_array_6_44_real <= _zz_154;
      end
      if(_zz_9)begin
        img_reg_array_7_44_real <= _zz_154;
      end
      if(_zz_10)begin
        img_reg_array_8_44_real <= _zz_154;
      end
      if(_zz_11)begin
        img_reg_array_9_44_real <= _zz_154;
      end
      if(_zz_12)begin
        img_reg_array_10_44_real <= _zz_154;
      end
      if(_zz_13)begin
        img_reg_array_11_44_real <= _zz_154;
      end
      if(_zz_14)begin
        img_reg_array_12_44_real <= _zz_154;
      end
      if(_zz_15)begin
        img_reg_array_13_44_real <= _zz_154;
      end
      if(_zz_16)begin
        img_reg_array_14_44_real <= _zz_154;
      end
      if(_zz_17)begin
        img_reg_array_15_44_real <= _zz_154;
      end
      if(_zz_18)begin
        img_reg_array_16_44_real <= _zz_154;
      end
      if(_zz_19)begin
        img_reg_array_17_44_real <= _zz_154;
      end
      if(_zz_20)begin
        img_reg_array_18_44_real <= _zz_154;
      end
      if(_zz_21)begin
        img_reg_array_19_44_real <= _zz_154;
      end
      if(_zz_22)begin
        img_reg_array_20_44_real <= _zz_154;
      end
      if(_zz_23)begin
        img_reg_array_21_44_real <= _zz_154;
      end
      if(_zz_24)begin
        img_reg_array_22_44_real <= _zz_154;
      end
      if(_zz_25)begin
        img_reg_array_23_44_real <= _zz_154;
      end
      if(_zz_26)begin
        img_reg_array_24_44_real <= _zz_154;
      end
      if(_zz_27)begin
        img_reg_array_25_44_real <= _zz_154;
      end
      if(_zz_28)begin
        img_reg_array_26_44_real <= _zz_154;
      end
      if(_zz_29)begin
        img_reg_array_27_44_real <= _zz_154;
      end
      if(_zz_30)begin
        img_reg_array_28_44_real <= _zz_154;
      end
      if(_zz_31)begin
        img_reg_array_29_44_real <= _zz_154;
      end
      if(_zz_32)begin
        img_reg_array_30_44_real <= _zz_154;
      end
      if(_zz_33)begin
        img_reg_array_31_44_real <= _zz_154;
      end
      if(_zz_34)begin
        img_reg_array_32_44_real <= _zz_154;
      end
      if(_zz_35)begin
        img_reg_array_33_44_real <= _zz_154;
      end
      if(_zz_36)begin
        img_reg_array_34_44_real <= _zz_154;
      end
      if(_zz_37)begin
        img_reg_array_35_44_real <= _zz_154;
      end
      if(_zz_38)begin
        img_reg_array_36_44_real <= _zz_154;
      end
      if(_zz_39)begin
        img_reg_array_37_44_real <= _zz_154;
      end
      if(_zz_40)begin
        img_reg_array_38_44_real <= _zz_154;
      end
      if(_zz_41)begin
        img_reg_array_39_44_real <= _zz_154;
      end
      if(_zz_42)begin
        img_reg_array_40_44_real <= _zz_154;
      end
      if(_zz_43)begin
        img_reg_array_41_44_real <= _zz_154;
      end
      if(_zz_44)begin
        img_reg_array_42_44_real <= _zz_154;
      end
      if(_zz_45)begin
        img_reg_array_43_44_real <= _zz_154;
      end
      if(_zz_46)begin
        img_reg_array_44_44_real <= _zz_154;
      end
      if(_zz_47)begin
        img_reg_array_45_44_real <= _zz_154;
      end
      if(_zz_48)begin
        img_reg_array_46_44_real <= _zz_154;
      end
      if(_zz_49)begin
        img_reg_array_47_44_real <= _zz_154;
      end
      if(_zz_50)begin
        img_reg_array_48_44_real <= _zz_154;
      end
      if(_zz_51)begin
        img_reg_array_49_44_real <= _zz_154;
      end
      if(_zz_52)begin
        img_reg_array_50_44_real <= _zz_154;
      end
      if(_zz_53)begin
        img_reg_array_51_44_real <= _zz_154;
      end
      if(_zz_54)begin
        img_reg_array_52_44_real <= _zz_154;
      end
      if(_zz_55)begin
        img_reg_array_53_44_real <= _zz_154;
      end
      if(_zz_56)begin
        img_reg_array_54_44_real <= _zz_154;
      end
      if(_zz_57)begin
        img_reg_array_55_44_real <= _zz_154;
      end
      if(_zz_58)begin
        img_reg_array_56_44_real <= _zz_154;
      end
      if(_zz_59)begin
        img_reg_array_57_44_real <= _zz_154;
      end
      if(_zz_60)begin
        img_reg_array_58_44_real <= _zz_154;
      end
      if(_zz_61)begin
        img_reg_array_59_44_real <= _zz_154;
      end
      if(_zz_62)begin
        img_reg_array_60_44_real <= _zz_154;
      end
      if(_zz_63)begin
        img_reg_array_61_44_real <= _zz_154;
      end
      if(_zz_64)begin
        img_reg_array_62_44_real <= _zz_154;
      end
      if(_zz_65)begin
        img_reg_array_63_44_real <= _zz_154;
      end
      if(_zz_2)begin
        img_reg_array_0_44_imag <= _zz_155;
      end
      if(_zz_3)begin
        img_reg_array_1_44_imag <= _zz_155;
      end
      if(_zz_4)begin
        img_reg_array_2_44_imag <= _zz_155;
      end
      if(_zz_5)begin
        img_reg_array_3_44_imag <= _zz_155;
      end
      if(_zz_6)begin
        img_reg_array_4_44_imag <= _zz_155;
      end
      if(_zz_7)begin
        img_reg_array_5_44_imag <= _zz_155;
      end
      if(_zz_8)begin
        img_reg_array_6_44_imag <= _zz_155;
      end
      if(_zz_9)begin
        img_reg_array_7_44_imag <= _zz_155;
      end
      if(_zz_10)begin
        img_reg_array_8_44_imag <= _zz_155;
      end
      if(_zz_11)begin
        img_reg_array_9_44_imag <= _zz_155;
      end
      if(_zz_12)begin
        img_reg_array_10_44_imag <= _zz_155;
      end
      if(_zz_13)begin
        img_reg_array_11_44_imag <= _zz_155;
      end
      if(_zz_14)begin
        img_reg_array_12_44_imag <= _zz_155;
      end
      if(_zz_15)begin
        img_reg_array_13_44_imag <= _zz_155;
      end
      if(_zz_16)begin
        img_reg_array_14_44_imag <= _zz_155;
      end
      if(_zz_17)begin
        img_reg_array_15_44_imag <= _zz_155;
      end
      if(_zz_18)begin
        img_reg_array_16_44_imag <= _zz_155;
      end
      if(_zz_19)begin
        img_reg_array_17_44_imag <= _zz_155;
      end
      if(_zz_20)begin
        img_reg_array_18_44_imag <= _zz_155;
      end
      if(_zz_21)begin
        img_reg_array_19_44_imag <= _zz_155;
      end
      if(_zz_22)begin
        img_reg_array_20_44_imag <= _zz_155;
      end
      if(_zz_23)begin
        img_reg_array_21_44_imag <= _zz_155;
      end
      if(_zz_24)begin
        img_reg_array_22_44_imag <= _zz_155;
      end
      if(_zz_25)begin
        img_reg_array_23_44_imag <= _zz_155;
      end
      if(_zz_26)begin
        img_reg_array_24_44_imag <= _zz_155;
      end
      if(_zz_27)begin
        img_reg_array_25_44_imag <= _zz_155;
      end
      if(_zz_28)begin
        img_reg_array_26_44_imag <= _zz_155;
      end
      if(_zz_29)begin
        img_reg_array_27_44_imag <= _zz_155;
      end
      if(_zz_30)begin
        img_reg_array_28_44_imag <= _zz_155;
      end
      if(_zz_31)begin
        img_reg_array_29_44_imag <= _zz_155;
      end
      if(_zz_32)begin
        img_reg_array_30_44_imag <= _zz_155;
      end
      if(_zz_33)begin
        img_reg_array_31_44_imag <= _zz_155;
      end
      if(_zz_34)begin
        img_reg_array_32_44_imag <= _zz_155;
      end
      if(_zz_35)begin
        img_reg_array_33_44_imag <= _zz_155;
      end
      if(_zz_36)begin
        img_reg_array_34_44_imag <= _zz_155;
      end
      if(_zz_37)begin
        img_reg_array_35_44_imag <= _zz_155;
      end
      if(_zz_38)begin
        img_reg_array_36_44_imag <= _zz_155;
      end
      if(_zz_39)begin
        img_reg_array_37_44_imag <= _zz_155;
      end
      if(_zz_40)begin
        img_reg_array_38_44_imag <= _zz_155;
      end
      if(_zz_41)begin
        img_reg_array_39_44_imag <= _zz_155;
      end
      if(_zz_42)begin
        img_reg_array_40_44_imag <= _zz_155;
      end
      if(_zz_43)begin
        img_reg_array_41_44_imag <= _zz_155;
      end
      if(_zz_44)begin
        img_reg_array_42_44_imag <= _zz_155;
      end
      if(_zz_45)begin
        img_reg_array_43_44_imag <= _zz_155;
      end
      if(_zz_46)begin
        img_reg_array_44_44_imag <= _zz_155;
      end
      if(_zz_47)begin
        img_reg_array_45_44_imag <= _zz_155;
      end
      if(_zz_48)begin
        img_reg_array_46_44_imag <= _zz_155;
      end
      if(_zz_49)begin
        img_reg_array_47_44_imag <= _zz_155;
      end
      if(_zz_50)begin
        img_reg_array_48_44_imag <= _zz_155;
      end
      if(_zz_51)begin
        img_reg_array_49_44_imag <= _zz_155;
      end
      if(_zz_52)begin
        img_reg_array_50_44_imag <= _zz_155;
      end
      if(_zz_53)begin
        img_reg_array_51_44_imag <= _zz_155;
      end
      if(_zz_54)begin
        img_reg_array_52_44_imag <= _zz_155;
      end
      if(_zz_55)begin
        img_reg_array_53_44_imag <= _zz_155;
      end
      if(_zz_56)begin
        img_reg_array_54_44_imag <= _zz_155;
      end
      if(_zz_57)begin
        img_reg_array_55_44_imag <= _zz_155;
      end
      if(_zz_58)begin
        img_reg_array_56_44_imag <= _zz_155;
      end
      if(_zz_59)begin
        img_reg_array_57_44_imag <= _zz_155;
      end
      if(_zz_60)begin
        img_reg_array_58_44_imag <= _zz_155;
      end
      if(_zz_61)begin
        img_reg_array_59_44_imag <= _zz_155;
      end
      if(_zz_62)begin
        img_reg_array_60_44_imag <= _zz_155;
      end
      if(_zz_63)begin
        img_reg_array_61_44_imag <= _zz_155;
      end
      if(_zz_64)begin
        img_reg_array_62_44_imag <= _zz_155;
      end
      if(_zz_65)begin
        img_reg_array_63_44_imag <= _zz_155;
      end
      if(_zz_2)begin
        img_reg_array_0_45_real <= _zz_156;
      end
      if(_zz_3)begin
        img_reg_array_1_45_real <= _zz_156;
      end
      if(_zz_4)begin
        img_reg_array_2_45_real <= _zz_156;
      end
      if(_zz_5)begin
        img_reg_array_3_45_real <= _zz_156;
      end
      if(_zz_6)begin
        img_reg_array_4_45_real <= _zz_156;
      end
      if(_zz_7)begin
        img_reg_array_5_45_real <= _zz_156;
      end
      if(_zz_8)begin
        img_reg_array_6_45_real <= _zz_156;
      end
      if(_zz_9)begin
        img_reg_array_7_45_real <= _zz_156;
      end
      if(_zz_10)begin
        img_reg_array_8_45_real <= _zz_156;
      end
      if(_zz_11)begin
        img_reg_array_9_45_real <= _zz_156;
      end
      if(_zz_12)begin
        img_reg_array_10_45_real <= _zz_156;
      end
      if(_zz_13)begin
        img_reg_array_11_45_real <= _zz_156;
      end
      if(_zz_14)begin
        img_reg_array_12_45_real <= _zz_156;
      end
      if(_zz_15)begin
        img_reg_array_13_45_real <= _zz_156;
      end
      if(_zz_16)begin
        img_reg_array_14_45_real <= _zz_156;
      end
      if(_zz_17)begin
        img_reg_array_15_45_real <= _zz_156;
      end
      if(_zz_18)begin
        img_reg_array_16_45_real <= _zz_156;
      end
      if(_zz_19)begin
        img_reg_array_17_45_real <= _zz_156;
      end
      if(_zz_20)begin
        img_reg_array_18_45_real <= _zz_156;
      end
      if(_zz_21)begin
        img_reg_array_19_45_real <= _zz_156;
      end
      if(_zz_22)begin
        img_reg_array_20_45_real <= _zz_156;
      end
      if(_zz_23)begin
        img_reg_array_21_45_real <= _zz_156;
      end
      if(_zz_24)begin
        img_reg_array_22_45_real <= _zz_156;
      end
      if(_zz_25)begin
        img_reg_array_23_45_real <= _zz_156;
      end
      if(_zz_26)begin
        img_reg_array_24_45_real <= _zz_156;
      end
      if(_zz_27)begin
        img_reg_array_25_45_real <= _zz_156;
      end
      if(_zz_28)begin
        img_reg_array_26_45_real <= _zz_156;
      end
      if(_zz_29)begin
        img_reg_array_27_45_real <= _zz_156;
      end
      if(_zz_30)begin
        img_reg_array_28_45_real <= _zz_156;
      end
      if(_zz_31)begin
        img_reg_array_29_45_real <= _zz_156;
      end
      if(_zz_32)begin
        img_reg_array_30_45_real <= _zz_156;
      end
      if(_zz_33)begin
        img_reg_array_31_45_real <= _zz_156;
      end
      if(_zz_34)begin
        img_reg_array_32_45_real <= _zz_156;
      end
      if(_zz_35)begin
        img_reg_array_33_45_real <= _zz_156;
      end
      if(_zz_36)begin
        img_reg_array_34_45_real <= _zz_156;
      end
      if(_zz_37)begin
        img_reg_array_35_45_real <= _zz_156;
      end
      if(_zz_38)begin
        img_reg_array_36_45_real <= _zz_156;
      end
      if(_zz_39)begin
        img_reg_array_37_45_real <= _zz_156;
      end
      if(_zz_40)begin
        img_reg_array_38_45_real <= _zz_156;
      end
      if(_zz_41)begin
        img_reg_array_39_45_real <= _zz_156;
      end
      if(_zz_42)begin
        img_reg_array_40_45_real <= _zz_156;
      end
      if(_zz_43)begin
        img_reg_array_41_45_real <= _zz_156;
      end
      if(_zz_44)begin
        img_reg_array_42_45_real <= _zz_156;
      end
      if(_zz_45)begin
        img_reg_array_43_45_real <= _zz_156;
      end
      if(_zz_46)begin
        img_reg_array_44_45_real <= _zz_156;
      end
      if(_zz_47)begin
        img_reg_array_45_45_real <= _zz_156;
      end
      if(_zz_48)begin
        img_reg_array_46_45_real <= _zz_156;
      end
      if(_zz_49)begin
        img_reg_array_47_45_real <= _zz_156;
      end
      if(_zz_50)begin
        img_reg_array_48_45_real <= _zz_156;
      end
      if(_zz_51)begin
        img_reg_array_49_45_real <= _zz_156;
      end
      if(_zz_52)begin
        img_reg_array_50_45_real <= _zz_156;
      end
      if(_zz_53)begin
        img_reg_array_51_45_real <= _zz_156;
      end
      if(_zz_54)begin
        img_reg_array_52_45_real <= _zz_156;
      end
      if(_zz_55)begin
        img_reg_array_53_45_real <= _zz_156;
      end
      if(_zz_56)begin
        img_reg_array_54_45_real <= _zz_156;
      end
      if(_zz_57)begin
        img_reg_array_55_45_real <= _zz_156;
      end
      if(_zz_58)begin
        img_reg_array_56_45_real <= _zz_156;
      end
      if(_zz_59)begin
        img_reg_array_57_45_real <= _zz_156;
      end
      if(_zz_60)begin
        img_reg_array_58_45_real <= _zz_156;
      end
      if(_zz_61)begin
        img_reg_array_59_45_real <= _zz_156;
      end
      if(_zz_62)begin
        img_reg_array_60_45_real <= _zz_156;
      end
      if(_zz_63)begin
        img_reg_array_61_45_real <= _zz_156;
      end
      if(_zz_64)begin
        img_reg_array_62_45_real <= _zz_156;
      end
      if(_zz_65)begin
        img_reg_array_63_45_real <= _zz_156;
      end
      if(_zz_2)begin
        img_reg_array_0_45_imag <= _zz_157;
      end
      if(_zz_3)begin
        img_reg_array_1_45_imag <= _zz_157;
      end
      if(_zz_4)begin
        img_reg_array_2_45_imag <= _zz_157;
      end
      if(_zz_5)begin
        img_reg_array_3_45_imag <= _zz_157;
      end
      if(_zz_6)begin
        img_reg_array_4_45_imag <= _zz_157;
      end
      if(_zz_7)begin
        img_reg_array_5_45_imag <= _zz_157;
      end
      if(_zz_8)begin
        img_reg_array_6_45_imag <= _zz_157;
      end
      if(_zz_9)begin
        img_reg_array_7_45_imag <= _zz_157;
      end
      if(_zz_10)begin
        img_reg_array_8_45_imag <= _zz_157;
      end
      if(_zz_11)begin
        img_reg_array_9_45_imag <= _zz_157;
      end
      if(_zz_12)begin
        img_reg_array_10_45_imag <= _zz_157;
      end
      if(_zz_13)begin
        img_reg_array_11_45_imag <= _zz_157;
      end
      if(_zz_14)begin
        img_reg_array_12_45_imag <= _zz_157;
      end
      if(_zz_15)begin
        img_reg_array_13_45_imag <= _zz_157;
      end
      if(_zz_16)begin
        img_reg_array_14_45_imag <= _zz_157;
      end
      if(_zz_17)begin
        img_reg_array_15_45_imag <= _zz_157;
      end
      if(_zz_18)begin
        img_reg_array_16_45_imag <= _zz_157;
      end
      if(_zz_19)begin
        img_reg_array_17_45_imag <= _zz_157;
      end
      if(_zz_20)begin
        img_reg_array_18_45_imag <= _zz_157;
      end
      if(_zz_21)begin
        img_reg_array_19_45_imag <= _zz_157;
      end
      if(_zz_22)begin
        img_reg_array_20_45_imag <= _zz_157;
      end
      if(_zz_23)begin
        img_reg_array_21_45_imag <= _zz_157;
      end
      if(_zz_24)begin
        img_reg_array_22_45_imag <= _zz_157;
      end
      if(_zz_25)begin
        img_reg_array_23_45_imag <= _zz_157;
      end
      if(_zz_26)begin
        img_reg_array_24_45_imag <= _zz_157;
      end
      if(_zz_27)begin
        img_reg_array_25_45_imag <= _zz_157;
      end
      if(_zz_28)begin
        img_reg_array_26_45_imag <= _zz_157;
      end
      if(_zz_29)begin
        img_reg_array_27_45_imag <= _zz_157;
      end
      if(_zz_30)begin
        img_reg_array_28_45_imag <= _zz_157;
      end
      if(_zz_31)begin
        img_reg_array_29_45_imag <= _zz_157;
      end
      if(_zz_32)begin
        img_reg_array_30_45_imag <= _zz_157;
      end
      if(_zz_33)begin
        img_reg_array_31_45_imag <= _zz_157;
      end
      if(_zz_34)begin
        img_reg_array_32_45_imag <= _zz_157;
      end
      if(_zz_35)begin
        img_reg_array_33_45_imag <= _zz_157;
      end
      if(_zz_36)begin
        img_reg_array_34_45_imag <= _zz_157;
      end
      if(_zz_37)begin
        img_reg_array_35_45_imag <= _zz_157;
      end
      if(_zz_38)begin
        img_reg_array_36_45_imag <= _zz_157;
      end
      if(_zz_39)begin
        img_reg_array_37_45_imag <= _zz_157;
      end
      if(_zz_40)begin
        img_reg_array_38_45_imag <= _zz_157;
      end
      if(_zz_41)begin
        img_reg_array_39_45_imag <= _zz_157;
      end
      if(_zz_42)begin
        img_reg_array_40_45_imag <= _zz_157;
      end
      if(_zz_43)begin
        img_reg_array_41_45_imag <= _zz_157;
      end
      if(_zz_44)begin
        img_reg_array_42_45_imag <= _zz_157;
      end
      if(_zz_45)begin
        img_reg_array_43_45_imag <= _zz_157;
      end
      if(_zz_46)begin
        img_reg_array_44_45_imag <= _zz_157;
      end
      if(_zz_47)begin
        img_reg_array_45_45_imag <= _zz_157;
      end
      if(_zz_48)begin
        img_reg_array_46_45_imag <= _zz_157;
      end
      if(_zz_49)begin
        img_reg_array_47_45_imag <= _zz_157;
      end
      if(_zz_50)begin
        img_reg_array_48_45_imag <= _zz_157;
      end
      if(_zz_51)begin
        img_reg_array_49_45_imag <= _zz_157;
      end
      if(_zz_52)begin
        img_reg_array_50_45_imag <= _zz_157;
      end
      if(_zz_53)begin
        img_reg_array_51_45_imag <= _zz_157;
      end
      if(_zz_54)begin
        img_reg_array_52_45_imag <= _zz_157;
      end
      if(_zz_55)begin
        img_reg_array_53_45_imag <= _zz_157;
      end
      if(_zz_56)begin
        img_reg_array_54_45_imag <= _zz_157;
      end
      if(_zz_57)begin
        img_reg_array_55_45_imag <= _zz_157;
      end
      if(_zz_58)begin
        img_reg_array_56_45_imag <= _zz_157;
      end
      if(_zz_59)begin
        img_reg_array_57_45_imag <= _zz_157;
      end
      if(_zz_60)begin
        img_reg_array_58_45_imag <= _zz_157;
      end
      if(_zz_61)begin
        img_reg_array_59_45_imag <= _zz_157;
      end
      if(_zz_62)begin
        img_reg_array_60_45_imag <= _zz_157;
      end
      if(_zz_63)begin
        img_reg_array_61_45_imag <= _zz_157;
      end
      if(_zz_64)begin
        img_reg_array_62_45_imag <= _zz_157;
      end
      if(_zz_65)begin
        img_reg_array_63_45_imag <= _zz_157;
      end
      if(_zz_2)begin
        img_reg_array_0_46_real <= _zz_158;
      end
      if(_zz_3)begin
        img_reg_array_1_46_real <= _zz_158;
      end
      if(_zz_4)begin
        img_reg_array_2_46_real <= _zz_158;
      end
      if(_zz_5)begin
        img_reg_array_3_46_real <= _zz_158;
      end
      if(_zz_6)begin
        img_reg_array_4_46_real <= _zz_158;
      end
      if(_zz_7)begin
        img_reg_array_5_46_real <= _zz_158;
      end
      if(_zz_8)begin
        img_reg_array_6_46_real <= _zz_158;
      end
      if(_zz_9)begin
        img_reg_array_7_46_real <= _zz_158;
      end
      if(_zz_10)begin
        img_reg_array_8_46_real <= _zz_158;
      end
      if(_zz_11)begin
        img_reg_array_9_46_real <= _zz_158;
      end
      if(_zz_12)begin
        img_reg_array_10_46_real <= _zz_158;
      end
      if(_zz_13)begin
        img_reg_array_11_46_real <= _zz_158;
      end
      if(_zz_14)begin
        img_reg_array_12_46_real <= _zz_158;
      end
      if(_zz_15)begin
        img_reg_array_13_46_real <= _zz_158;
      end
      if(_zz_16)begin
        img_reg_array_14_46_real <= _zz_158;
      end
      if(_zz_17)begin
        img_reg_array_15_46_real <= _zz_158;
      end
      if(_zz_18)begin
        img_reg_array_16_46_real <= _zz_158;
      end
      if(_zz_19)begin
        img_reg_array_17_46_real <= _zz_158;
      end
      if(_zz_20)begin
        img_reg_array_18_46_real <= _zz_158;
      end
      if(_zz_21)begin
        img_reg_array_19_46_real <= _zz_158;
      end
      if(_zz_22)begin
        img_reg_array_20_46_real <= _zz_158;
      end
      if(_zz_23)begin
        img_reg_array_21_46_real <= _zz_158;
      end
      if(_zz_24)begin
        img_reg_array_22_46_real <= _zz_158;
      end
      if(_zz_25)begin
        img_reg_array_23_46_real <= _zz_158;
      end
      if(_zz_26)begin
        img_reg_array_24_46_real <= _zz_158;
      end
      if(_zz_27)begin
        img_reg_array_25_46_real <= _zz_158;
      end
      if(_zz_28)begin
        img_reg_array_26_46_real <= _zz_158;
      end
      if(_zz_29)begin
        img_reg_array_27_46_real <= _zz_158;
      end
      if(_zz_30)begin
        img_reg_array_28_46_real <= _zz_158;
      end
      if(_zz_31)begin
        img_reg_array_29_46_real <= _zz_158;
      end
      if(_zz_32)begin
        img_reg_array_30_46_real <= _zz_158;
      end
      if(_zz_33)begin
        img_reg_array_31_46_real <= _zz_158;
      end
      if(_zz_34)begin
        img_reg_array_32_46_real <= _zz_158;
      end
      if(_zz_35)begin
        img_reg_array_33_46_real <= _zz_158;
      end
      if(_zz_36)begin
        img_reg_array_34_46_real <= _zz_158;
      end
      if(_zz_37)begin
        img_reg_array_35_46_real <= _zz_158;
      end
      if(_zz_38)begin
        img_reg_array_36_46_real <= _zz_158;
      end
      if(_zz_39)begin
        img_reg_array_37_46_real <= _zz_158;
      end
      if(_zz_40)begin
        img_reg_array_38_46_real <= _zz_158;
      end
      if(_zz_41)begin
        img_reg_array_39_46_real <= _zz_158;
      end
      if(_zz_42)begin
        img_reg_array_40_46_real <= _zz_158;
      end
      if(_zz_43)begin
        img_reg_array_41_46_real <= _zz_158;
      end
      if(_zz_44)begin
        img_reg_array_42_46_real <= _zz_158;
      end
      if(_zz_45)begin
        img_reg_array_43_46_real <= _zz_158;
      end
      if(_zz_46)begin
        img_reg_array_44_46_real <= _zz_158;
      end
      if(_zz_47)begin
        img_reg_array_45_46_real <= _zz_158;
      end
      if(_zz_48)begin
        img_reg_array_46_46_real <= _zz_158;
      end
      if(_zz_49)begin
        img_reg_array_47_46_real <= _zz_158;
      end
      if(_zz_50)begin
        img_reg_array_48_46_real <= _zz_158;
      end
      if(_zz_51)begin
        img_reg_array_49_46_real <= _zz_158;
      end
      if(_zz_52)begin
        img_reg_array_50_46_real <= _zz_158;
      end
      if(_zz_53)begin
        img_reg_array_51_46_real <= _zz_158;
      end
      if(_zz_54)begin
        img_reg_array_52_46_real <= _zz_158;
      end
      if(_zz_55)begin
        img_reg_array_53_46_real <= _zz_158;
      end
      if(_zz_56)begin
        img_reg_array_54_46_real <= _zz_158;
      end
      if(_zz_57)begin
        img_reg_array_55_46_real <= _zz_158;
      end
      if(_zz_58)begin
        img_reg_array_56_46_real <= _zz_158;
      end
      if(_zz_59)begin
        img_reg_array_57_46_real <= _zz_158;
      end
      if(_zz_60)begin
        img_reg_array_58_46_real <= _zz_158;
      end
      if(_zz_61)begin
        img_reg_array_59_46_real <= _zz_158;
      end
      if(_zz_62)begin
        img_reg_array_60_46_real <= _zz_158;
      end
      if(_zz_63)begin
        img_reg_array_61_46_real <= _zz_158;
      end
      if(_zz_64)begin
        img_reg_array_62_46_real <= _zz_158;
      end
      if(_zz_65)begin
        img_reg_array_63_46_real <= _zz_158;
      end
      if(_zz_2)begin
        img_reg_array_0_46_imag <= _zz_159;
      end
      if(_zz_3)begin
        img_reg_array_1_46_imag <= _zz_159;
      end
      if(_zz_4)begin
        img_reg_array_2_46_imag <= _zz_159;
      end
      if(_zz_5)begin
        img_reg_array_3_46_imag <= _zz_159;
      end
      if(_zz_6)begin
        img_reg_array_4_46_imag <= _zz_159;
      end
      if(_zz_7)begin
        img_reg_array_5_46_imag <= _zz_159;
      end
      if(_zz_8)begin
        img_reg_array_6_46_imag <= _zz_159;
      end
      if(_zz_9)begin
        img_reg_array_7_46_imag <= _zz_159;
      end
      if(_zz_10)begin
        img_reg_array_8_46_imag <= _zz_159;
      end
      if(_zz_11)begin
        img_reg_array_9_46_imag <= _zz_159;
      end
      if(_zz_12)begin
        img_reg_array_10_46_imag <= _zz_159;
      end
      if(_zz_13)begin
        img_reg_array_11_46_imag <= _zz_159;
      end
      if(_zz_14)begin
        img_reg_array_12_46_imag <= _zz_159;
      end
      if(_zz_15)begin
        img_reg_array_13_46_imag <= _zz_159;
      end
      if(_zz_16)begin
        img_reg_array_14_46_imag <= _zz_159;
      end
      if(_zz_17)begin
        img_reg_array_15_46_imag <= _zz_159;
      end
      if(_zz_18)begin
        img_reg_array_16_46_imag <= _zz_159;
      end
      if(_zz_19)begin
        img_reg_array_17_46_imag <= _zz_159;
      end
      if(_zz_20)begin
        img_reg_array_18_46_imag <= _zz_159;
      end
      if(_zz_21)begin
        img_reg_array_19_46_imag <= _zz_159;
      end
      if(_zz_22)begin
        img_reg_array_20_46_imag <= _zz_159;
      end
      if(_zz_23)begin
        img_reg_array_21_46_imag <= _zz_159;
      end
      if(_zz_24)begin
        img_reg_array_22_46_imag <= _zz_159;
      end
      if(_zz_25)begin
        img_reg_array_23_46_imag <= _zz_159;
      end
      if(_zz_26)begin
        img_reg_array_24_46_imag <= _zz_159;
      end
      if(_zz_27)begin
        img_reg_array_25_46_imag <= _zz_159;
      end
      if(_zz_28)begin
        img_reg_array_26_46_imag <= _zz_159;
      end
      if(_zz_29)begin
        img_reg_array_27_46_imag <= _zz_159;
      end
      if(_zz_30)begin
        img_reg_array_28_46_imag <= _zz_159;
      end
      if(_zz_31)begin
        img_reg_array_29_46_imag <= _zz_159;
      end
      if(_zz_32)begin
        img_reg_array_30_46_imag <= _zz_159;
      end
      if(_zz_33)begin
        img_reg_array_31_46_imag <= _zz_159;
      end
      if(_zz_34)begin
        img_reg_array_32_46_imag <= _zz_159;
      end
      if(_zz_35)begin
        img_reg_array_33_46_imag <= _zz_159;
      end
      if(_zz_36)begin
        img_reg_array_34_46_imag <= _zz_159;
      end
      if(_zz_37)begin
        img_reg_array_35_46_imag <= _zz_159;
      end
      if(_zz_38)begin
        img_reg_array_36_46_imag <= _zz_159;
      end
      if(_zz_39)begin
        img_reg_array_37_46_imag <= _zz_159;
      end
      if(_zz_40)begin
        img_reg_array_38_46_imag <= _zz_159;
      end
      if(_zz_41)begin
        img_reg_array_39_46_imag <= _zz_159;
      end
      if(_zz_42)begin
        img_reg_array_40_46_imag <= _zz_159;
      end
      if(_zz_43)begin
        img_reg_array_41_46_imag <= _zz_159;
      end
      if(_zz_44)begin
        img_reg_array_42_46_imag <= _zz_159;
      end
      if(_zz_45)begin
        img_reg_array_43_46_imag <= _zz_159;
      end
      if(_zz_46)begin
        img_reg_array_44_46_imag <= _zz_159;
      end
      if(_zz_47)begin
        img_reg_array_45_46_imag <= _zz_159;
      end
      if(_zz_48)begin
        img_reg_array_46_46_imag <= _zz_159;
      end
      if(_zz_49)begin
        img_reg_array_47_46_imag <= _zz_159;
      end
      if(_zz_50)begin
        img_reg_array_48_46_imag <= _zz_159;
      end
      if(_zz_51)begin
        img_reg_array_49_46_imag <= _zz_159;
      end
      if(_zz_52)begin
        img_reg_array_50_46_imag <= _zz_159;
      end
      if(_zz_53)begin
        img_reg_array_51_46_imag <= _zz_159;
      end
      if(_zz_54)begin
        img_reg_array_52_46_imag <= _zz_159;
      end
      if(_zz_55)begin
        img_reg_array_53_46_imag <= _zz_159;
      end
      if(_zz_56)begin
        img_reg_array_54_46_imag <= _zz_159;
      end
      if(_zz_57)begin
        img_reg_array_55_46_imag <= _zz_159;
      end
      if(_zz_58)begin
        img_reg_array_56_46_imag <= _zz_159;
      end
      if(_zz_59)begin
        img_reg_array_57_46_imag <= _zz_159;
      end
      if(_zz_60)begin
        img_reg_array_58_46_imag <= _zz_159;
      end
      if(_zz_61)begin
        img_reg_array_59_46_imag <= _zz_159;
      end
      if(_zz_62)begin
        img_reg_array_60_46_imag <= _zz_159;
      end
      if(_zz_63)begin
        img_reg_array_61_46_imag <= _zz_159;
      end
      if(_zz_64)begin
        img_reg_array_62_46_imag <= _zz_159;
      end
      if(_zz_65)begin
        img_reg_array_63_46_imag <= _zz_159;
      end
      if(_zz_2)begin
        img_reg_array_0_47_real <= _zz_160;
      end
      if(_zz_3)begin
        img_reg_array_1_47_real <= _zz_160;
      end
      if(_zz_4)begin
        img_reg_array_2_47_real <= _zz_160;
      end
      if(_zz_5)begin
        img_reg_array_3_47_real <= _zz_160;
      end
      if(_zz_6)begin
        img_reg_array_4_47_real <= _zz_160;
      end
      if(_zz_7)begin
        img_reg_array_5_47_real <= _zz_160;
      end
      if(_zz_8)begin
        img_reg_array_6_47_real <= _zz_160;
      end
      if(_zz_9)begin
        img_reg_array_7_47_real <= _zz_160;
      end
      if(_zz_10)begin
        img_reg_array_8_47_real <= _zz_160;
      end
      if(_zz_11)begin
        img_reg_array_9_47_real <= _zz_160;
      end
      if(_zz_12)begin
        img_reg_array_10_47_real <= _zz_160;
      end
      if(_zz_13)begin
        img_reg_array_11_47_real <= _zz_160;
      end
      if(_zz_14)begin
        img_reg_array_12_47_real <= _zz_160;
      end
      if(_zz_15)begin
        img_reg_array_13_47_real <= _zz_160;
      end
      if(_zz_16)begin
        img_reg_array_14_47_real <= _zz_160;
      end
      if(_zz_17)begin
        img_reg_array_15_47_real <= _zz_160;
      end
      if(_zz_18)begin
        img_reg_array_16_47_real <= _zz_160;
      end
      if(_zz_19)begin
        img_reg_array_17_47_real <= _zz_160;
      end
      if(_zz_20)begin
        img_reg_array_18_47_real <= _zz_160;
      end
      if(_zz_21)begin
        img_reg_array_19_47_real <= _zz_160;
      end
      if(_zz_22)begin
        img_reg_array_20_47_real <= _zz_160;
      end
      if(_zz_23)begin
        img_reg_array_21_47_real <= _zz_160;
      end
      if(_zz_24)begin
        img_reg_array_22_47_real <= _zz_160;
      end
      if(_zz_25)begin
        img_reg_array_23_47_real <= _zz_160;
      end
      if(_zz_26)begin
        img_reg_array_24_47_real <= _zz_160;
      end
      if(_zz_27)begin
        img_reg_array_25_47_real <= _zz_160;
      end
      if(_zz_28)begin
        img_reg_array_26_47_real <= _zz_160;
      end
      if(_zz_29)begin
        img_reg_array_27_47_real <= _zz_160;
      end
      if(_zz_30)begin
        img_reg_array_28_47_real <= _zz_160;
      end
      if(_zz_31)begin
        img_reg_array_29_47_real <= _zz_160;
      end
      if(_zz_32)begin
        img_reg_array_30_47_real <= _zz_160;
      end
      if(_zz_33)begin
        img_reg_array_31_47_real <= _zz_160;
      end
      if(_zz_34)begin
        img_reg_array_32_47_real <= _zz_160;
      end
      if(_zz_35)begin
        img_reg_array_33_47_real <= _zz_160;
      end
      if(_zz_36)begin
        img_reg_array_34_47_real <= _zz_160;
      end
      if(_zz_37)begin
        img_reg_array_35_47_real <= _zz_160;
      end
      if(_zz_38)begin
        img_reg_array_36_47_real <= _zz_160;
      end
      if(_zz_39)begin
        img_reg_array_37_47_real <= _zz_160;
      end
      if(_zz_40)begin
        img_reg_array_38_47_real <= _zz_160;
      end
      if(_zz_41)begin
        img_reg_array_39_47_real <= _zz_160;
      end
      if(_zz_42)begin
        img_reg_array_40_47_real <= _zz_160;
      end
      if(_zz_43)begin
        img_reg_array_41_47_real <= _zz_160;
      end
      if(_zz_44)begin
        img_reg_array_42_47_real <= _zz_160;
      end
      if(_zz_45)begin
        img_reg_array_43_47_real <= _zz_160;
      end
      if(_zz_46)begin
        img_reg_array_44_47_real <= _zz_160;
      end
      if(_zz_47)begin
        img_reg_array_45_47_real <= _zz_160;
      end
      if(_zz_48)begin
        img_reg_array_46_47_real <= _zz_160;
      end
      if(_zz_49)begin
        img_reg_array_47_47_real <= _zz_160;
      end
      if(_zz_50)begin
        img_reg_array_48_47_real <= _zz_160;
      end
      if(_zz_51)begin
        img_reg_array_49_47_real <= _zz_160;
      end
      if(_zz_52)begin
        img_reg_array_50_47_real <= _zz_160;
      end
      if(_zz_53)begin
        img_reg_array_51_47_real <= _zz_160;
      end
      if(_zz_54)begin
        img_reg_array_52_47_real <= _zz_160;
      end
      if(_zz_55)begin
        img_reg_array_53_47_real <= _zz_160;
      end
      if(_zz_56)begin
        img_reg_array_54_47_real <= _zz_160;
      end
      if(_zz_57)begin
        img_reg_array_55_47_real <= _zz_160;
      end
      if(_zz_58)begin
        img_reg_array_56_47_real <= _zz_160;
      end
      if(_zz_59)begin
        img_reg_array_57_47_real <= _zz_160;
      end
      if(_zz_60)begin
        img_reg_array_58_47_real <= _zz_160;
      end
      if(_zz_61)begin
        img_reg_array_59_47_real <= _zz_160;
      end
      if(_zz_62)begin
        img_reg_array_60_47_real <= _zz_160;
      end
      if(_zz_63)begin
        img_reg_array_61_47_real <= _zz_160;
      end
      if(_zz_64)begin
        img_reg_array_62_47_real <= _zz_160;
      end
      if(_zz_65)begin
        img_reg_array_63_47_real <= _zz_160;
      end
      if(_zz_2)begin
        img_reg_array_0_47_imag <= _zz_161;
      end
      if(_zz_3)begin
        img_reg_array_1_47_imag <= _zz_161;
      end
      if(_zz_4)begin
        img_reg_array_2_47_imag <= _zz_161;
      end
      if(_zz_5)begin
        img_reg_array_3_47_imag <= _zz_161;
      end
      if(_zz_6)begin
        img_reg_array_4_47_imag <= _zz_161;
      end
      if(_zz_7)begin
        img_reg_array_5_47_imag <= _zz_161;
      end
      if(_zz_8)begin
        img_reg_array_6_47_imag <= _zz_161;
      end
      if(_zz_9)begin
        img_reg_array_7_47_imag <= _zz_161;
      end
      if(_zz_10)begin
        img_reg_array_8_47_imag <= _zz_161;
      end
      if(_zz_11)begin
        img_reg_array_9_47_imag <= _zz_161;
      end
      if(_zz_12)begin
        img_reg_array_10_47_imag <= _zz_161;
      end
      if(_zz_13)begin
        img_reg_array_11_47_imag <= _zz_161;
      end
      if(_zz_14)begin
        img_reg_array_12_47_imag <= _zz_161;
      end
      if(_zz_15)begin
        img_reg_array_13_47_imag <= _zz_161;
      end
      if(_zz_16)begin
        img_reg_array_14_47_imag <= _zz_161;
      end
      if(_zz_17)begin
        img_reg_array_15_47_imag <= _zz_161;
      end
      if(_zz_18)begin
        img_reg_array_16_47_imag <= _zz_161;
      end
      if(_zz_19)begin
        img_reg_array_17_47_imag <= _zz_161;
      end
      if(_zz_20)begin
        img_reg_array_18_47_imag <= _zz_161;
      end
      if(_zz_21)begin
        img_reg_array_19_47_imag <= _zz_161;
      end
      if(_zz_22)begin
        img_reg_array_20_47_imag <= _zz_161;
      end
      if(_zz_23)begin
        img_reg_array_21_47_imag <= _zz_161;
      end
      if(_zz_24)begin
        img_reg_array_22_47_imag <= _zz_161;
      end
      if(_zz_25)begin
        img_reg_array_23_47_imag <= _zz_161;
      end
      if(_zz_26)begin
        img_reg_array_24_47_imag <= _zz_161;
      end
      if(_zz_27)begin
        img_reg_array_25_47_imag <= _zz_161;
      end
      if(_zz_28)begin
        img_reg_array_26_47_imag <= _zz_161;
      end
      if(_zz_29)begin
        img_reg_array_27_47_imag <= _zz_161;
      end
      if(_zz_30)begin
        img_reg_array_28_47_imag <= _zz_161;
      end
      if(_zz_31)begin
        img_reg_array_29_47_imag <= _zz_161;
      end
      if(_zz_32)begin
        img_reg_array_30_47_imag <= _zz_161;
      end
      if(_zz_33)begin
        img_reg_array_31_47_imag <= _zz_161;
      end
      if(_zz_34)begin
        img_reg_array_32_47_imag <= _zz_161;
      end
      if(_zz_35)begin
        img_reg_array_33_47_imag <= _zz_161;
      end
      if(_zz_36)begin
        img_reg_array_34_47_imag <= _zz_161;
      end
      if(_zz_37)begin
        img_reg_array_35_47_imag <= _zz_161;
      end
      if(_zz_38)begin
        img_reg_array_36_47_imag <= _zz_161;
      end
      if(_zz_39)begin
        img_reg_array_37_47_imag <= _zz_161;
      end
      if(_zz_40)begin
        img_reg_array_38_47_imag <= _zz_161;
      end
      if(_zz_41)begin
        img_reg_array_39_47_imag <= _zz_161;
      end
      if(_zz_42)begin
        img_reg_array_40_47_imag <= _zz_161;
      end
      if(_zz_43)begin
        img_reg_array_41_47_imag <= _zz_161;
      end
      if(_zz_44)begin
        img_reg_array_42_47_imag <= _zz_161;
      end
      if(_zz_45)begin
        img_reg_array_43_47_imag <= _zz_161;
      end
      if(_zz_46)begin
        img_reg_array_44_47_imag <= _zz_161;
      end
      if(_zz_47)begin
        img_reg_array_45_47_imag <= _zz_161;
      end
      if(_zz_48)begin
        img_reg_array_46_47_imag <= _zz_161;
      end
      if(_zz_49)begin
        img_reg_array_47_47_imag <= _zz_161;
      end
      if(_zz_50)begin
        img_reg_array_48_47_imag <= _zz_161;
      end
      if(_zz_51)begin
        img_reg_array_49_47_imag <= _zz_161;
      end
      if(_zz_52)begin
        img_reg_array_50_47_imag <= _zz_161;
      end
      if(_zz_53)begin
        img_reg_array_51_47_imag <= _zz_161;
      end
      if(_zz_54)begin
        img_reg_array_52_47_imag <= _zz_161;
      end
      if(_zz_55)begin
        img_reg_array_53_47_imag <= _zz_161;
      end
      if(_zz_56)begin
        img_reg_array_54_47_imag <= _zz_161;
      end
      if(_zz_57)begin
        img_reg_array_55_47_imag <= _zz_161;
      end
      if(_zz_58)begin
        img_reg_array_56_47_imag <= _zz_161;
      end
      if(_zz_59)begin
        img_reg_array_57_47_imag <= _zz_161;
      end
      if(_zz_60)begin
        img_reg_array_58_47_imag <= _zz_161;
      end
      if(_zz_61)begin
        img_reg_array_59_47_imag <= _zz_161;
      end
      if(_zz_62)begin
        img_reg_array_60_47_imag <= _zz_161;
      end
      if(_zz_63)begin
        img_reg_array_61_47_imag <= _zz_161;
      end
      if(_zz_64)begin
        img_reg_array_62_47_imag <= _zz_161;
      end
      if(_zz_65)begin
        img_reg_array_63_47_imag <= _zz_161;
      end
      if(_zz_2)begin
        img_reg_array_0_48_real <= _zz_162;
      end
      if(_zz_3)begin
        img_reg_array_1_48_real <= _zz_162;
      end
      if(_zz_4)begin
        img_reg_array_2_48_real <= _zz_162;
      end
      if(_zz_5)begin
        img_reg_array_3_48_real <= _zz_162;
      end
      if(_zz_6)begin
        img_reg_array_4_48_real <= _zz_162;
      end
      if(_zz_7)begin
        img_reg_array_5_48_real <= _zz_162;
      end
      if(_zz_8)begin
        img_reg_array_6_48_real <= _zz_162;
      end
      if(_zz_9)begin
        img_reg_array_7_48_real <= _zz_162;
      end
      if(_zz_10)begin
        img_reg_array_8_48_real <= _zz_162;
      end
      if(_zz_11)begin
        img_reg_array_9_48_real <= _zz_162;
      end
      if(_zz_12)begin
        img_reg_array_10_48_real <= _zz_162;
      end
      if(_zz_13)begin
        img_reg_array_11_48_real <= _zz_162;
      end
      if(_zz_14)begin
        img_reg_array_12_48_real <= _zz_162;
      end
      if(_zz_15)begin
        img_reg_array_13_48_real <= _zz_162;
      end
      if(_zz_16)begin
        img_reg_array_14_48_real <= _zz_162;
      end
      if(_zz_17)begin
        img_reg_array_15_48_real <= _zz_162;
      end
      if(_zz_18)begin
        img_reg_array_16_48_real <= _zz_162;
      end
      if(_zz_19)begin
        img_reg_array_17_48_real <= _zz_162;
      end
      if(_zz_20)begin
        img_reg_array_18_48_real <= _zz_162;
      end
      if(_zz_21)begin
        img_reg_array_19_48_real <= _zz_162;
      end
      if(_zz_22)begin
        img_reg_array_20_48_real <= _zz_162;
      end
      if(_zz_23)begin
        img_reg_array_21_48_real <= _zz_162;
      end
      if(_zz_24)begin
        img_reg_array_22_48_real <= _zz_162;
      end
      if(_zz_25)begin
        img_reg_array_23_48_real <= _zz_162;
      end
      if(_zz_26)begin
        img_reg_array_24_48_real <= _zz_162;
      end
      if(_zz_27)begin
        img_reg_array_25_48_real <= _zz_162;
      end
      if(_zz_28)begin
        img_reg_array_26_48_real <= _zz_162;
      end
      if(_zz_29)begin
        img_reg_array_27_48_real <= _zz_162;
      end
      if(_zz_30)begin
        img_reg_array_28_48_real <= _zz_162;
      end
      if(_zz_31)begin
        img_reg_array_29_48_real <= _zz_162;
      end
      if(_zz_32)begin
        img_reg_array_30_48_real <= _zz_162;
      end
      if(_zz_33)begin
        img_reg_array_31_48_real <= _zz_162;
      end
      if(_zz_34)begin
        img_reg_array_32_48_real <= _zz_162;
      end
      if(_zz_35)begin
        img_reg_array_33_48_real <= _zz_162;
      end
      if(_zz_36)begin
        img_reg_array_34_48_real <= _zz_162;
      end
      if(_zz_37)begin
        img_reg_array_35_48_real <= _zz_162;
      end
      if(_zz_38)begin
        img_reg_array_36_48_real <= _zz_162;
      end
      if(_zz_39)begin
        img_reg_array_37_48_real <= _zz_162;
      end
      if(_zz_40)begin
        img_reg_array_38_48_real <= _zz_162;
      end
      if(_zz_41)begin
        img_reg_array_39_48_real <= _zz_162;
      end
      if(_zz_42)begin
        img_reg_array_40_48_real <= _zz_162;
      end
      if(_zz_43)begin
        img_reg_array_41_48_real <= _zz_162;
      end
      if(_zz_44)begin
        img_reg_array_42_48_real <= _zz_162;
      end
      if(_zz_45)begin
        img_reg_array_43_48_real <= _zz_162;
      end
      if(_zz_46)begin
        img_reg_array_44_48_real <= _zz_162;
      end
      if(_zz_47)begin
        img_reg_array_45_48_real <= _zz_162;
      end
      if(_zz_48)begin
        img_reg_array_46_48_real <= _zz_162;
      end
      if(_zz_49)begin
        img_reg_array_47_48_real <= _zz_162;
      end
      if(_zz_50)begin
        img_reg_array_48_48_real <= _zz_162;
      end
      if(_zz_51)begin
        img_reg_array_49_48_real <= _zz_162;
      end
      if(_zz_52)begin
        img_reg_array_50_48_real <= _zz_162;
      end
      if(_zz_53)begin
        img_reg_array_51_48_real <= _zz_162;
      end
      if(_zz_54)begin
        img_reg_array_52_48_real <= _zz_162;
      end
      if(_zz_55)begin
        img_reg_array_53_48_real <= _zz_162;
      end
      if(_zz_56)begin
        img_reg_array_54_48_real <= _zz_162;
      end
      if(_zz_57)begin
        img_reg_array_55_48_real <= _zz_162;
      end
      if(_zz_58)begin
        img_reg_array_56_48_real <= _zz_162;
      end
      if(_zz_59)begin
        img_reg_array_57_48_real <= _zz_162;
      end
      if(_zz_60)begin
        img_reg_array_58_48_real <= _zz_162;
      end
      if(_zz_61)begin
        img_reg_array_59_48_real <= _zz_162;
      end
      if(_zz_62)begin
        img_reg_array_60_48_real <= _zz_162;
      end
      if(_zz_63)begin
        img_reg_array_61_48_real <= _zz_162;
      end
      if(_zz_64)begin
        img_reg_array_62_48_real <= _zz_162;
      end
      if(_zz_65)begin
        img_reg_array_63_48_real <= _zz_162;
      end
      if(_zz_2)begin
        img_reg_array_0_48_imag <= _zz_163;
      end
      if(_zz_3)begin
        img_reg_array_1_48_imag <= _zz_163;
      end
      if(_zz_4)begin
        img_reg_array_2_48_imag <= _zz_163;
      end
      if(_zz_5)begin
        img_reg_array_3_48_imag <= _zz_163;
      end
      if(_zz_6)begin
        img_reg_array_4_48_imag <= _zz_163;
      end
      if(_zz_7)begin
        img_reg_array_5_48_imag <= _zz_163;
      end
      if(_zz_8)begin
        img_reg_array_6_48_imag <= _zz_163;
      end
      if(_zz_9)begin
        img_reg_array_7_48_imag <= _zz_163;
      end
      if(_zz_10)begin
        img_reg_array_8_48_imag <= _zz_163;
      end
      if(_zz_11)begin
        img_reg_array_9_48_imag <= _zz_163;
      end
      if(_zz_12)begin
        img_reg_array_10_48_imag <= _zz_163;
      end
      if(_zz_13)begin
        img_reg_array_11_48_imag <= _zz_163;
      end
      if(_zz_14)begin
        img_reg_array_12_48_imag <= _zz_163;
      end
      if(_zz_15)begin
        img_reg_array_13_48_imag <= _zz_163;
      end
      if(_zz_16)begin
        img_reg_array_14_48_imag <= _zz_163;
      end
      if(_zz_17)begin
        img_reg_array_15_48_imag <= _zz_163;
      end
      if(_zz_18)begin
        img_reg_array_16_48_imag <= _zz_163;
      end
      if(_zz_19)begin
        img_reg_array_17_48_imag <= _zz_163;
      end
      if(_zz_20)begin
        img_reg_array_18_48_imag <= _zz_163;
      end
      if(_zz_21)begin
        img_reg_array_19_48_imag <= _zz_163;
      end
      if(_zz_22)begin
        img_reg_array_20_48_imag <= _zz_163;
      end
      if(_zz_23)begin
        img_reg_array_21_48_imag <= _zz_163;
      end
      if(_zz_24)begin
        img_reg_array_22_48_imag <= _zz_163;
      end
      if(_zz_25)begin
        img_reg_array_23_48_imag <= _zz_163;
      end
      if(_zz_26)begin
        img_reg_array_24_48_imag <= _zz_163;
      end
      if(_zz_27)begin
        img_reg_array_25_48_imag <= _zz_163;
      end
      if(_zz_28)begin
        img_reg_array_26_48_imag <= _zz_163;
      end
      if(_zz_29)begin
        img_reg_array_27_48_imag <= _zz_163;
      end
      if(_zz_30)begin
        img_reg_array_28_48_imag <= _zz_163;
      end
      if(_zz_31)begin
        img_reg_array_29_48_imag <= _zz_163;
      end
      if(_zz_32)begin
        img_reg_array_30_48_imag <= _zz_163;
      end
      if(_zz_33)begin
        img_reg_array_31_48_imag <= _zz_163;
      end
      if(_zz_34)begin
        img_reg_array_32_48_imag <= _zz_163;
      end
      if(_zz_35)begin
        img_reg_array_33_48_imag <= _zz_163;
      end
      if(_zz_36)begin
        img_reg_array_34_48_imag <= _zz_163;
      end
      if(_zz_37)begin
        img_reg_array_35_48_imag <= _zz_163;
      end
      if(_zz_38)begin
        img_reg_array_36_48_imag <= _zz_163;
      end
      if(_zz_39)begin
        img_reg_array_37_48_imag <= _zz_163;
      end
      if(_zz_40)begin
        img_reg_array_38_48_imag <= _zz_163;
      end
      if(_zz_41)begin
        img_reg_array_39_48_imag <= _zz_163;
      end
      if(_zz_42)begin
        img_reg_array_40_48_imag <= _zz_163;
      end
      if(_zz_43)begin
        img_reg_array_41_48_imag <= _zz_163;
      end
      if(_zz_44)begin
        img_reg_array_42_48_imag <= _zz_163;
      end
      if(_zz_45)begin
        img_reg_array_43_48_imag <= _zz_163;
      end
      if(_zz_46)begin
        img_reg_array_44_48_imag <= _zz_163;
      end
      if(_zz_47)begin
        img_reg_array_45_48_imag <= _zz_163;
      end
      if(_zz_48)begin
        img_reg_array_46_48_imag <= _zz_163;
      end
      if(_zz_49)begin
        img_reg_array_47_48_imag <= _zz_163;
      end
      if(_zz_50)begin
        img_reg_array_48_48_imag <= _zz_163;
      end
      if(_zz_51)begin
        img_reg_array_49_48_imag <= _zz_163;
      end
      if(_zz_52)begin
        img_reg_array_50_48_imag <= _zz_163;
      end
      if(_zz_53)begin
        img_reg_array_51_48_imag <= _zz_163;
      end
      if(_zz_54)begin
        img_reg_array_52_48_imag <= _zz_163;
      end
      if(_zz_55)begin
        img_reg_array_53_48_imag <= _zz_163;
      end
      if(_zz_56)begin
        img_reg_array_54_48_imag <= _zz_163;
      end
      if(_zz_57)begin
        img_reg_array_55_48_imag <= _zz_163;
      end
      if(_zz_58)begin
        img_reg_array_56_48_imag <= _zz_163;
      end
      if(_zz_59)begin
        img_reg_array_57_48_imag <= _zz_163;
      end
      if(_zz_60)begin
        img_reg_array_58_48_imag <= _zz_163;
      end
      if(_zz_61)begin
        img_reg_array_59_48_imag <= _zz_163;
      end
      if(_zz_62)begin
        img_reg_array_60_48_imag <= _zz_163;
      end
      if(_zz_63)begin
        img_reg_array_61_48_imag <= _zz_163;
      end
      if(_zz_64)begin
        img_reg_array_62_48_imag <= _zz_163;
      end
      if(_zz_65)begin
        img_reg_array_63_48_imag <= _zz_163;
      end
      if(_zz_2)begin
        img_reg_array_0_49_real <= _zz_164;
      end
      if(_zz_3)begin
        img_reg_array_1_49_real <= _zz_164;
      end
      if(_zz_4)begin
        img_reg_array_2_49_real <= _zz_164;
      end
      if(_zz_5)begin
        img_reg_array_3_49_real <= _zz_164;
      end
      if(_zz_6)begin
        img_reg_array_4_49_real <= _zz_164;
      end
      if(_zz_7)begin
        img_reg_array_5_49_real <= _zz_164;
      end
      if(_zz_8)begin
        img_reg_array_6_49_real <= _zz_164;
      end
      if(_zz_9)begin
        img_reg_array_7_49_real <= _zz_164;
      end
      if(_zz_10)begin
        img_reg_array_8_49_real <= _zz_164;
      end
      if(_zz_11)begin
        img_reg_array_9_49_real <= _zz_164;
      end
      if(_zz_12)begin
        img_reg_array_10_49_real <= _zz_164;
      end
      if(_zz_13)begin
        img_reg_array_11_49_real <= _zz_164;
      end
      if(_zz_14)begin
        img_reg_array_12_49_real <= _zz_164;
      end
      if(_zz_15)begin
        img_reg_array_13_49_real <= _zz_164;
      end
      if(_zz_16)begin
        img_reg_array_14_49_real <= _zz_164;
      end
      if(_zz_17)begin
        img_reg_array_15_49_real <= _zz_164;
      end
      if(_zz_18)begin
        img_reg_array_16_49_real <= _zz_164;
      end
      if(_zz_19)begin
        img_reg_array_17_49_real <= _zz_164;
      end
      if(_zz_20)begin
        img_reg_array_18_49_real <= _zz_164;
      end
      if(_zz_21)begin
        img_reg_array_19_49_real <= _zz_164;
      end
      if(_zz_22)begin
        img_reg_array_20_49_real <= _zz_164;
      end
      if(_zz_23)begin
        img_reg_array_21_49_real <= _zz_164;
      end
      if(_zz_24)begin
        img_reg_array_22_49_real <= _zz_164;
      end
      if(_zz_25)begin
        img_reg_array_23_49_real <= _zz_164;
      end
      if(_zz_26)begin
        img_reg_array_24_49_real <= _zz_164;
      end
      if(_zz_27)begin
        img_reg_array_25_49_real <= _zz_164;
      end
      if(_zz_28)begin
        img_reg_array_26_49_real <= _zz_164;
      end
      if(_zz_29)begin
        img_reg_array_27_49_real <= _zz_164;
      end
      if(_zz_30)begin
        img_reg_array_28_49_real <= _zz_164;
      end
      if(_zz_31)begin
        img_reg_array_29_49_real <= _zz_164;
      end
      if(_zz_32)begin
        img_reg_array_30_49_real <= _zz_164;
      end
      if(_zz_33)begin
        img_reg_array_31_49_real <= _zz_164;
      end
      if(_zz_34)begin
        img_reg_array_32_49_real <= _zz_164;
      end
      if(_zz_35)begin
        img_reg_array_33_49_real <= _zz_164;
      end
      if(_zz_36)begin
        img_reg_array_34_49_real <= _zz_164;
      end
      if(_zz_37)begin
        img_reg_array_35_49_real <= _zz_164;
      end
      if(_zz_38)begin
        img_reg_array_36_49_real <= _zz_164;
      end
      if(_zz_39)begin
        img_reg_array_37_49_real <= _zz_164;
      end
      if(_zz_40)begin
        img_reg_array_38_49_real <= _zz_164;
      end
      if(_zz_41)begin
        img_reg_array_39_49_real <= _zz_164;
      end
      if(_zz_42)begin
        img_reg_array_40_49_real <= _zz_164;
      end
      if(_zz_43)begin
        img_reg_array_41_49_real <= _zz_164;
      end
      if(_zz_44)begin
        img_reg_array_42_49_real <= _zz_164;
      end
      if(_zz_45)begin
        img_reg_array_43_49_real <= _zz_164;
      end
      if(_zz_46)begin
        img_reg_array_44_49_real <= _zz_164;
      end
      if(_zz_47)begin
        img_reg_array_45_49_real <= _zz_164;
      end
      if(_zz_48)begin
        img_reg_array_46_49_real <= _zz_164;
      end
      if(_zz_49)begin
        img_reg_array_47_49_real <= _zz_164;
      end
      if(_zz_50)begin
        img_reg_array_48_49_real <= _zz_164;
      end
      if(_zz_51)begin
        img_reg_array_49_49_real <= _zz_164;
      end
      if(_zz_52)begin
        img_reg_array_50_49_real <= _zz_164;
      end
      if(_zz_53)begin
        img_reg_array_51_49_real <= _zz_164;
      end
      if(_zz_54)begin
        img_reg_array_52_49_real <= _zz_164;
      end
      if(_zz_55)begin
        img_reg_array_53_49_real <= _zz_164;
      end
      if(_zz_56)begin
        img_reg_array_54_49_real <= _zz_164;
      end
      if(_zz_57)begin
        img_reg_array_55_49_real <= _zz_164;
      end
      if(_zz_58)begin
        img_reg_array_56_49_real <= _zz_164;
      end
      if(_zz_59)begin
        img_reg_array_57_49_real <= _zz_164;
      end
      if(_zz_60)begin
        img_reg_array_58_49_real <= _zz_164;
      end
      if(_zz_61)begin
        img_reg_array_59_49_real <= _zz_164;
      end
      if(_zz_62)begin
        img_reg_array_60_49_real <= _zz_164;
      end
      if(_zz_63)begin
        img_reg_array_61_49_real <= _zz_164;
      end
      if(_zz_64)begin
        img_reg_array_62_49_real <= _zz_164;
      end
      if(_zz_65)begin
        img_reg_array_63_49_real <= _zz_164;
      end
      if(_zz_2)begin
        img_reg_array_0_49_imag <= _zz_165;
      end
      if(_zz_3)begin
        img_reg_array_1_49_imag <= _zz_165;
      end
      if(_zz_4)begin
        img_reg_array_2_49_imag <= _zz_165;
      end
      if(_zz_5)begin
        img_reg_array_3_49_imag <= _zz_165;
      end
      if(_zz_6)begin
        img_reg_array_4_49_imag <= _zz_165;
      end
      if(_zz_7)begin
        img_reg_array_5_49_imag <= _zz_165;
      end
      if(_zz_8)begin
        img_reg_array_6_49_imag <= _zz_165;
      end
      if(_zz_9)begin
        img_reg_array_7_49_imag <= _zz_165;
      end
      if(_zz_10)begin
        img_reg_array_8_49_imag <= _zz_165;
      end
      if(_zz_11)begin
        img_reg_array_9_49_imag <= _zz_165;
      end
      if(_zz_12)begin
        img_reg_array_10_49_imag <= _zz_165;
      end
      if(_zz_13)begin
        img_reg_array_11_49_imag <= _zz_165;
      end
      if(_zz_14)begin
        img_reg_array_12_49_imag <= _zz_165;
      end
      if(_zz_15)begin
        img_reg_array_13_49_imag <= _zz_165;
      end
      if(_zz_16)begin
        img_reg_array_14_49_imag <= _zz_165;
      end
      if(_zz_17)begin
        img_reg_array_15_49_imag <= _zz_165;
      end
      if(_zz_18)begin
        img_reg_array_16_49_imag <= _zz_165;
      end
      if(_zz_19)begin
        img_reg_array_17_49_imag <= _zz_165;
      end
      if(_zz_20)begin
        img_reg_array_18_49_imag <= _zz_165;
      end
      if(_zz_21)begin
        img_reg_array_19_49_imag <= _zz_165;
      end
      if(_zz_22)begin
        img_reg_array_20_49_imag <= _zz_165;
      end
      if(_zz_23)begin
        img_reg_array_21_49_imag <= _zz_165;
      end
      if(_zz_24)begin
        img_reg_array_22_49_imag <= _zz_165;
      end
      if(_zz_25)begin
        img_reg_array_23_49_imag <= _zz_165;
      end
      if(_zz_26)begin
        img_reg_array_24_49_imag <= _zz_165;
      end
      if(_zz_27)begin
        img_reg_array_25_49_imag <= _zz_165;
      end
      if(_zz_28)begin
        img_reg_array_26_49_imag <= _zz_165;
      end
      if(_zz_29)begin
        img_reg_array_27_49_imag <= _zz_165;
      end
      if(_zz_30)begin
        img_reg_array_28_49_imag <= _zz_165;
      end
      if(_zz_31)begin
        img_reg_array_29_49_imag <= _zz_165;
      end
      if(_zz_32)begin
        img_reg_array_30_49_imag <= _zz_165;
      end
      if(_zz_33)begin
        img_reg_array_31_49_imag <= _zz_165;
      end
      if(_zz_34)begin
        img_reg_array_32_49_imag <= _zz_165;
      end
      if(_zz_35)begin
        img_reg_array_33_49_imag <= _zz_165;
      end
      if(_zz_36)begin
        img_reg_array_34_49_imag <= _zz_165;
      end
      if(_zz_37)begin
        img_reg_array_35_49_imag <= _zz_165;
      end
      if(_zz_38)begin
        img_reg_array_36_49_imag <= _zz_165;
      end
      if(_zz_39)begin
        img_reg_array_37_49_imag <= _zz_165;
      end
      if(_zz_40)begin
        img_reg_array_38_49_imag <= _zz_165;
      end
      if(_zz_41)begin
        img_reg_array_39_49_imag <= _zz_165;
      end
      if(_zz_42)begin
        img_reg_array_40_49_imag <= _zz_165;
      end
      if(_zz_43)begin
        img_reg_array_41_49_imag <= _zz_165;
      end
      if(_zz_44)begin
        img_reg_array_42_49_imag <= _zz_165;
      end
      if(_zz_45)begin
        img_reg_array_43_49_imag <= _zz_165;
      end
      if(_zz_46)begin
        img_reg_array_44_49_imag <= _zz_165;
      end
      if(_zz_47)begin
        img_reg_array_45_49_imag <= _zz_165;
      end
      if(_zz_48)begin
        img_reg_array_46_49_imag <= _zz_165;
      end
      if(_zz_49)begin
        img_reg_array_47_49_imag <= _zz_165;
      end
      if(_zz_50)begin
        img_reg_array_48_49_imag <= _zz_165;
      end
      if(_zz_51)begin
        img_reg_array_49_49_imag <= _zz_165;
      end
      if(_zz_52)begin
        img_reg_array_50_49_imag <= _zz_165;
      end
      if(_zz_53)begin
        img_reg_array_51_49_imag <= _zz_165;
      end
      if(_zz_54)begin
        img_reg_array_52_49_imag <= _zz_165;
      end
      if(_zz_55)begin
        img_reg_array_53_49_imag <= _zz_165;
      end
      if(_zz_56)begin
        img_reg_array_54_49_imag <= _zz_165;
      end
      if(_zz_57)begin
        img_reg_array_55_49_imag <= _zz_165;
      end
      if(_zz_58)begin
        img_reg_array_56_49_imag <= _zz_165;
      end
      if(_zz_59)begin
        img_reg_array_57_49_imag <= _zz_165;
      end
      if(_zz_60)begin
        img_reg_array_58_49_imag <= _zz_165;
      end
      if(_zz_61)begin
        img_reg_array_59_49_imag <= _zz_165;
      end
      if(_zz_62)begin
        img_reg_array_60_49_imag <= _zz_165;
      end
      if(_zz_63)begin
        img_reg_array_61_49_imag <= _zz_165;
      end
      if(_zz_64)begin
        img_reg_array_62_49_imag <= _zz_165;
      end
      if(_zz_65)begin
        img_reg_array_63_49_imag <= _zz_165;
      end
      if(_zz_2)begin
        img_reg_array_0_50_real <= _zz_166;
      end
      if(_zz_3)begin
        img_reg_array_1_50_real <= _zz_166;
      end
      if(_zz_4)begin
        img_reg_array_2_50_real <= _zz_166;
      end
      if(_zz_5)begin
        img_reg_array_3_50_real <= _zz_166;
      end
      if(_zz_6)begin
        img_reg_array_4_50_real <= _zz_166;
      end
      if(_zz_7)begin
        img_reg_array_5_50_real <= _zz_166;
      end
      if(_zz_8)begin
        img_reg_array_6_50_real <= _zz_166;
      end
      if(_zz_9)begin
        img_reg_array_7_50_real <= _zz_166;
      end
      if(_zz_10)begin
        img_reg_array_8_50_real <= _zz_166;
      end
      if(_zz_11)begin
        img_reg_array_9_50_real <= _zz_166;
      end
      if(_zz_12)begin
        img_reg_array_10_50_real <= _zz_166;
      end
      if(_zz_13)begin
        img_reg_array_11_50_real <= _zz_166;
      end
      if(_zz_14)begin
        img_reg_array_12_50_real <= _zz_166;
      end
      if(_zz_15)begin
        img_reg_array_13_50_real <= _zz_166;
      end
      if(_zz_16)begin
        img_reg_array_14_50_real <= _zz_166;
      end
      if(_zz_17)begin
        img_reg_array_15_50_real <= _zz_166;
      end
      if(_zz_18)begin
        img_reg_array_16_50_real <= _zz_166;
      end
      if(_zz_19)begin
        img_reg_array_17_50_real <= _zz_166;
      end
      if(_zz_20)begin
        img_reg_array_18_50_real <= _zz_166;
      end
      if(_zz_21)begin
        img_reg_array_19_50_real <= _zz_166;
      end
      if(_zz_22)begin
        img_reg_array_20_50_real <= _zz_166;
      end
      if(_zz_23)begin
        img_reg_array_21_50_real <= _zz_166;
      end
      if(_zz_24)begin
        img_reg_array_22_50_real <= _zz_166;
      end
      if(_zz_25)begin
        img_reg_array_23_50_real <= _zz_166;
      end
      if(_zz_26)begin
        img_reg_array_24_50_real <= _zz_166;
      end
      if(_zz_27)begin
        img_reg_array_25_50_real <= _zz_166;
      end
      if(_zz_28)begin
        img_reg_array_26_50_real <= _zz_166;
      end
      if(_zz_29)begin
        img_reg_array_27_50_real <= _zz_166;
      end
      if(_zz_30)begin
        img_reg_array_28_50_real <= _zz_166;
      end
      if(_zz_31)begin
        img_reg_array_29_50_real <= _zz_166;
      end
      if(_zz_32)begin
        img_reg_array_30_50_real <= _zz_166;
      end
      if(_zz_33)begin
        img_reg_array_31_50_real <= _zz_166;
      end
      if(_zz_34)begin
        img_reg_array_32_50_real <= _zz_166;
      end
      if(_zz_35)begin
        img_reg_array_33_50_real <= _zz_166;
      end
      if(_zz_36)begin
        img_reg_array_34_50_real <= _zz_166;
      end
      if(_zz_37)begin
        img_reg_array_35_50_real <= _zz_166;
      end
      if(_zz_38)begin
        img_reg_array_36_50_real <= _zz_166;
      end
      if(_zz_39)begin
        img_reg_array_37_50_real <= _zz_166;
      end
      if(_zz_40)begin
        img_reg_array_38_50_real <= _zz_166;
      end
      if(_zz_41)begin
        img_reg_array_39_50_real <= _zz_166;
      end
      if(_zz_42)begin
        img_reg_array_40_50_real <= _zz_166;
      end
      if(_zz_43)begin
        img_reg_array_41_50_real <= _zz_166;
      end
      if(_zz_44)begin
        img_reg_array_42_50_real <= _zz_166;
      end
      if(_zz_45)begin
        img_reg_array_43_50_real <= _zz_166;
      end
      if(_zz_46)begin
        img_reg_array_44_50_real <= _zz_166;
      end
      if(_zz_47)begin
        img_reg_array_45_50_real <= _zz_166;
      end
      if(_zz_48)begin
        img_reg_array_46_50_real <= _zz_166;
      end
      if(_zz_49)begin
        img_reg_array_47_50_real <= _zz_166;
      end
      if(_zz_50)begin
        img_reg_array_48_50_real <= _zz_166;
      end
      if(_zz_51)begin
        img_reg_array_49_50_real <= _zz_166;
      end
      if(_zz_52)begin
        img_reg_array_50_50_real <= _zz_166;
      end
      if(_zz_53)begin
        img_reg_array_51_50_real <= _zz_166;
      end
      if(_zz_54)begin
        img_reg_array_52_50_real <= _zz_166;
      end
      if(_zz_55)begin
        img_reg_array_53_50_real <= _zz_166;
      end
      if(_zz_56)begin
        img_reg_array_54_50_real <= _zz_166;
      end
      if(_zz_57)begin
        img_reg_array_55_50_real <= _zz_166;
      end
      if(_zz_58)begin
        img_reg_array_56_50_real <= _zz_166;
      end
      if(_zz_59)begin
        img_reg_array_57_50_real <= _zz_166;
      end
      if(_zz_60)begin
        img_reg_array_58_50_real <= _zz_166;
      end
      if(_zz_61)begin
        img_reg_array_59_50_real <= _zz_166;
      end
      if(_zz_62)begin
        img_reg_array_60_50_real <= _zz_166;
      end
      if(_zz_63)begin
        img_reg_array_61_50_real <= _zz_166;
      end
      if(_zz_64)begin
        img_reg_array_62_50_real <= _zz_166;
      end
      if(_zz_65)begin
        img_reg_array_63_50_real <= _zz_166;
      end
      if(_zz_2)begin
        img_reg_array_0_50_imag <= _zz_167;
      end
      if(_zz_3)begin
        img_reg_array_1_50_imag <= _zz_167;
      end
      if(_zz_4)begin
        img_reg_array_2_50_imag <= _zz_167;
      end
      if(_zz_5)begin
        img_reg_array_3_50_imag <= _zz_167;
      end
      if(_zz_6)begin
        img_reg_array_4_50_imag <= _zz_167;
      end
      if(_zz_7)begin
        img_reg_array_5_50_imag <= _zz_167;
      end
      if(_zz_8)begin
        img_reg_array_6_50_imag <= _zz_167;
      end
      if(_zz_9)begin
        img_reg_array_7_50_imag <= _zz_167;
      end
      if(_zz_10)begin
        img_reg_array_8_50_imag <= _zz_167;
      end
      if(_zz_11)begin
        img_reg_array_9_50_imag <= _zz_167;
      end
      if(_zz_12)begin
        img_reg_array_10_50_imag <= _zz_167;
      end
      if(_zz_13)begin
        img_reg_array_11_50_imag <= _zz_167;
      end
      if(_zz_14)begin
        img_reg_array_12_50_imag <= _zz_167;
      end
      if(_zz_15)begin
        img_reg_array_13_50_imag <= _zz_167;
      end
      if(_zz_16)begin
        img_reg_array_14_50_imag <= _zz_167;
      end
      if(_zz_17)begin
        img_reg_array_15_50_imag <= _zz_167;
      end
      if(_zz_18)begin
        img_reg_array_16_50_imag <= _zz_167;
      end
      if(_zz_19)begin
        img_reg_array_17_50_imag <= _zz_167;
      end
      if(_zz_20)begin
        img_reg_array_18_50_imag <= _zz_167;
      end
      if(_zz_21)begin
        img_reg_array_19_50_imag <= _zz_167;
      end
      if(_zz_22)begin
        img_reg_array_20_50_imag <= _zz_167;
      end
      if(_zz_23)begin
        img_reg_array_21_50_imag <= _zz_167;
      end
      if(_zz_24)begin
        img_reg_array_22_50_imag <= _zz_167;
      end
      if(_zz_25)begin
        img_reg_array_23_50_imag <= _zz_167;
      end
      if(_zz_26)begin
        img_reg_array_24_50_imag <= _zz_167;
      end
      if(_zz_27)begin
        img_reg_array_25_50_imag <= _zz_167;
      end
      if(_zz_28)begin
        img_reg_array_26_50_imag <= _zz_167;
      end
      if(_zz_29)begin
        img_reg_array_27_50_imag <= _zz_167;
      end
      if(_zz_30)begin
        img_reg_array_28_50_imag <= _zz_167;
      end
      if(_zz_31)begin
        img_reg_array_29_50_imag <= _zz_167;
      end
      if(_zz_32)begin
        img_reg_array_30_50_imag <= _zz_167;
      end
      if(_zz_33)begin
        img_reg_array_31_50_imag <= _zz_167;
      end
      if(_zz_34)begin
        img_reg_array_32_50_imag <= _zz_167;
      end
      if(_zz_35)begin
        img_reg_array_33_50_imag <= _zz_167;
      end
      if(_zz_36)begin
        img_reg_array_34_50_imag <= _zz_167;
      end
      if(_zz_37)begin
        img_reg_array_35_50_imag <= _zz_167;
      end
      if(_zz_38)begin
        img_reg_array_36_50_imag <= _zz_167;
      end
      if(_zz_39)begin
        img_reg_array_37_50_imag <= _zz_167;
      end
      if(_zz_40)begin
        img_reg_array_38_50_imag <= _zz_167;
      end
      if(_zz_41)begin
        img_reg_array_39_50_imag <= _zz_167;
      end
      if(_zz_42)begin
        img_reg_array_40_50_imag <= _zz_167;
      end
      if(_zz_43)begin
        img_reg_array_41_50_imag <= _zz_167;
      end
      if(_zz_44)begin
        img_reg_array_42_50_imag <= _zz_167;
      end
      if(_zz_45)begin
        img_reg_array_43_50_imag <= _zz_167;
      end
      if(_zz_46)begin
        img_reg_array_44_50_imag <= _zz_167;
      end
      if(_zz_47)begin
        img_reg_array_45_50_imag <= _zz_167;
      end
      if(_zz_48)begin
        img_reg_array_46_50_imag <= _zz_167;
      end
      if(_zz_49)begin
        img_reg_array_47_50_imag <= _zz_167;
      end
      if(_zz_50)begin
        img_reg_array_48_50_imag <= _zz_167;
      end
      if(_zz_51)begin
        img_reg_array_49_50_imag <= _zz_167;
      end
      if(_zz_52)begin
        img_reg_array_50_50_imag <= _zz_167;
      end
      if(_zz_53)begin
        img_reg_array_51_50_imag <= _zz_167;
      end
      if(_zz_54)begin
        img_reg_array_52_50_imag <= _zz_167;
      end
      if(_zz_55)begin
        img_reg_array_53_50_imag <= _zz_167;
      end
      if(_zz_56)begin
        img_reg_array_54_50_imag <= _zz_167;
      end
      if(_zz_57)begin
        img_reg_array_55_50_imag <= _zz_167;
      end
      if(_zz_58)begin
        img_reg_array_56_50_imag <= _zz_167;
      end
      if(_zz_59)begin
        img_reg_array_57_50_imag <= _zz_167;
      end
      if(_zz_60)begin
        img_reg_array_58_50_imag <= _zz_167;
      end
      if(_zz_61)begin
        img_reg_array_59_50_imag <= _zz_167;
      end
      if(_zz_62)begin
        img_reg_array_60_50_imag <= _zz_167;
      end
      if(_zz_63)begin
        img_reg_array_61_50_imag <= _zz_167;
      end
      if(_zz_64)begin
        img_reg_array_62_50_imag <= _zz_167;
      end
      if(_zz_65)begin
        img_reg_array_63_50_imag <= _zz_167;
      end
      if(_zz_2)begin
        img_reg_array_0_51_real <= _zz_168;
      end
      if(_zz_3)begin
        img_reg_array_1_51_real <= _zz_168;
      end
      if(_zz_4)begin
        img_reg_array_2_51_real <= _zz_168;
      end
      if(_zz_5)begin
        img_reg_array_3_51_real <= _zz_168;
      end
      if(_zz_6)begin
        img_reg_array_4_51_real <= _zz_168;
      end
      if(_zz_7)begin
        img_reg_array_5_51_real <= _zz_168;
      end
      if(_zz_8)begin
        img_reg_array_6_51_real <= _zz_168;
      end
      if(_zz_9)begin
        img_reg_array_7_51_real <= _zz_168;
      end
      if(_zz_10)begin
        img_reg_array_8_51_real <= _zz_168;
      end
      if(_zz_11)begin
        img_reg_array_9_51_real <= _zz_168;
      end
      if(_zz_12)begin
        img_reg_array_10_51_real <= _zz_168;
      end
      if(_zz_13)begin
        img_reg_array_11_51_real <= _zz_168;
      end
      if(_zz_14)begin
        img_reg_array_12_51_real <= _zz_168;
      end
      if(_zz_15)begin
        img_reg_array_13_51_real <= _zz_168;
      end
      if(_zz_16)begin
        img_reg_array_14_51_real <= _zz_168;
      end
      if(_zz_17)begin
        img_reg_array_15_51_real <= _zz_168;
      end
      if(_zz_18)begin
        img_reg_array_16_51_real <= _zz_168;
      end
      if(_zz_19)begin
        img_reg_array_17_51_real <= _zz_168;
      end
      if(_zz_20)begin
        img_reg_array_18_51_real <= _zz_168;
      end
      if(_zz_21)begin
        img_reg_array_19_51_real <= _zz_168;
      end
      if(_zz_22)begin
        img_reg_array_20_51_real <= _zz_168;
      end
      if(_zz_23)begin
        img_reg_array_21_51_real <= _zz_168;
      end
      if(_zz_24)begin
        img_reg_array_22_51_real <= _zz_168;
      end
      if(_zz_25)begin
        img_reg_array_23_51_real <= _zz_168;
      end
      if(_zz_26)begin
        img_reg_array_24_51_real <= _zz_168;
      end
      if(_zz_27)begin
        img_reg_array_25_51_real <= _zz_168;
      end
      if(_zz_28)begin
        img_reg_array_26_51_real <= _zz_168;
      end
      if(_zz_29)begin
        img_reg_array_27_51_real <= _zz_168;
      end
      if(_zz_30)begin
        img_reg_array_28_51_real <= _zz_168;
      end
      if(_zz_31)begin
        img_reg_array_29_51_real <= _zz_168;
      end
      if(_zz_32)begin
        img_reg_array_30_51_real <= _zz_168;
      end
      if(_zz_33)begin
        img_reg_array_31_51_real <= _zz_168;
      end
      if(_zz_34)begin
        img_reg_array_32_51_real <= _zz_168;
      end
      if(_zz_35)begin
        img_reg_array_33_51_real <= _zz_168;
      end
      if(_zz_36)begin
        img_reg_array_34_51_real <= _zz_168;
      end
      if(_zz_37)begin
        img_reg_array_35_51_real <= _zz_168;
      end
      if(_zz_38)begin
        img_reg_array_36_51_real <= _zz_168;
      end
      if(_zz_39)begin
        img_reg_array_37_51_real <= _zz_168;
      end
      if(_zz_40)begin
        img_reg_array_38_51_real <= _zz_168;
      end
      if(_zz_41)begin
        img_reg_array_39_51_real <= _zz_168;
      end
      if(_zz_42)begin
        img_reg_array_40_51_real <= _zz_168;
      end
      if(_zz_43)begin
        img_reg_array_41_51_real <= _zz_168;
      end
      if(_zz_44)begin
        img_reg_array_42_51_real <= _zz_168;
      end
      if(_zz_45)begin
        img_reg_array_43_51_real <= _zz_168;
      end
      if(_zz_46)begin
        img_reg_array_44_51_real <= _zz_168;
      end
      if(_zz_47)begin
        img_reg_array_45_51_real <= _zz_168;
      end
      if(_zz_48)begin
        img_reg_array_46_51_real <= _zz_168;
      end
      if(_zz_49)begin
        img_reg_array_47_51_real <= _zz_168;
      end
      if(_zz_50)begin
        img_reg_array_48_51_real <= _zz_168;
      end
      if(_zz_51)begin
        img_reg_array_49_51_real <= _zz_168;
      end
      if(_zz_52)begin
        img_reg_array_50_51_real <= _zz_168;
      end
      if(_zz_53)begin
        img_reg_array_51_51_real <= _zz_168;
      end
      if(_zz_54)begin
        img_reg_array_52_51_real <= _zz_168;
      end
      if(_zz_55)begin
        img_reg_array_53_51_real <= _zz_168;
      end
      if(_zz_56)begin
        img_reg_array_54_51_real <= _zz_168;
      end
      if(_zz_57)begin
        img_reg_array_55_51_real <= _zz_168;
      end
      if(_zz_58)begin
        img_reg_array_56_51_real <= _zz_168;
      end
      if(_zz_59)begin
        img_reg_array_57_51_real <= _zz_168;
      end
      if(_zz_60)begin
        img_reg_array_58_51_real <= _zz_168;
      end
      if(_zz_61)begin
        img_reg_array_59_51_real <= _zz_168;
      end
      if(_zz_62)begin
        img_reg_array_60_51_real <= _zz_168;
      end
      if(_zz_63)begin
        img_reg_array_61_51_real <= _zz_168;
      end
      if(_zz_64)begin
        img_reg_array_62_51_real <= _zz_168;
      end
      if(_zz_65)begin
        img_reg_array_63_51_real <= _zz_168;
      end
      if(_zz_2)begin
        img_reg_array_0_51_imag <= _zz_169;
      end
      if(_zz_3)begin
        img_reg_array_1_51_imag <= _zz_169;
      end
      if(_zz_4)begin
        img_reg_array_2_51_imag <= _zz_169;
      end
      if(_zz_5)begin
        img_reg_array_3_51_imag <= _zz_169;
      end
      if(_zz_6)begin
        img_reg_array_4_51_imag <= _zz_169;
      end
      if(_zz_7)begin
        img_reg_array_5_51_imag <= _zz_169;
      end
      if(_zz_8)begin
        img_reg_array_6_51_imag <= _zz_169;
      end
      if(_zz_9)begin
        img_reg_array_7_51_imag <= _zz_169;
      end
      if(_zz_10)begin
        img_reg_array_8_51_imag <= _zz_169;
      end
      if(_zz_11)begin
        img_reg_array_9_51_imag <= _zz_169;
      end
      if(_zz_12)begin
        img_reg_array_10_51_imag <= _zz_169;
      end
      if(_zz_13)begin
        img_reg_array_11_51_imag <= _zz_169;
      end
      if(_zz_14)begin
        img_reg_array_12_51_imag <= _zz_169;
      end
      if(_zz_15)begin
        img_reg_array_13_51_imag <= _zz_169;
      end
      if(_zz_16)begin
        img_reg_array_14_51_imag <= _zz_169;
      end
      if(_zz_17)begin
        img_reg_array_15_51_imag <= _zz_169;
      end
      if(_zz_18)begin
        img_reg_array_16_51_imag <= _zz_169;
      end
      if(_zz_19)begin
        img_reg_array_17_51_imag <= _zz_169;
      end
      if(_zz_20)begin
        img_reg_array_18_51_imag <= _zz_169;
      end
      if(_zz_21)begin
        img_reg_array_19_51_imag <= _zz_169;
      end
      if(_zz_22)begin
        img_reg_array_20_51_imag <= _zz_169;
      end
      if(_zz_23)begin
        img_reg_array_21_51_imag <= _zz_169;
      end
      if(_zz_24)begin
        img_reg_array_22_51_imag <= _zz_169;
      end
      if(_zz_25)begin
        img_reg_array_23_51_imag <= _zz_169;
      end
      if(_zz_26)begin
        img_reg_array_24_51_imag <= _zz_169;
      end
      if(_zz_27)begin
        img_reg_array_25_51_imag <= _zz_169;
      end
      if(_zz_28)begin
        img_reg_array_26_51_imag <= _zz_169;
      end
      if(_zz_29)begin
        img_reg_array_27_51_imag <= _zz_169;
      end
      if(_zz_30)begin
        img_reg_array_28_51_imag <= _zz_169;
      end
      if(_zz_31)begin
        img_reg_array_29_51_imag <= _zz_169;
      end
      if(_zz_32)begin
        img_reg_array_30_51_imag <= _zz_169;
      end
      if(_zz_33)begin
        img_reg_array_31_51_imag <= _zz_169;
      end
      if(_zz_34)begin
        img_reg_array_32_51_imag <= _zz_169;
      end
      if(_zz_35)begin
        img_reg_array_33_51_imag <= _zz_169;
      end
      if(_zz_36)begin
        img_reg_array_34_51_imag <= _zz_169;
      end
      if(_zz_37)begin
        img_reg_array_35_51_imag <= _zz_169;
      end
      if(_zz_38)begin
        img_reg_array_36_51_imag <= _zz_169;
      end
      if(_zz_39)begin
        img_reg_array_37_51_imag <= _zz_169;
      end
      if(_zz_40)begin
        img_reg_array_38_51_imag <= _zz_169;
      end
      if(_zz_41)begin
        img_reg_array_39_51_imag <= _zz_169;
      end
      if(_zz_42)begin
        img_reg_array_40_51_imag <= _zz_169;
      end
      if(_zz_43)begin
        img_reg_array_41_51_imag <= _zz_169;
      end
      if(_zz_44)begin
        img_reg_array_42_51_imag <= _zz_169;
      end
      if(_zz_45)begin
        img_reg_array_43_51_imag <= _zz_169;
      end
      if(_zz_46)begin
        img_reg_array_44_51_imag <= _zz_169;
      end
      if(_zz_47)begin
        img_reg_array_45_51_imag <= _zz_169;
      end
      if(_zz_48)begin
        img_reg_array_46_51_imag <= _zz_169;
      end
      if(_zz_49)begin
        img_reg_array_47_51_imag <= _zz_169;
      end
      if(_zz_50)begin
        img_reg_array_48_51_imag <= _zz_169;
      end
      if(_zz_51)begin
        img_reg_array_49_51_imag <= _zz_169;
      end
      if(_zz_52)begin
        img_reg_array_50_51_imag <= _zz_169;
      end
      if(_zz_53)begin
        img_reg_array_51_51_imag <= _zz_169;
      end
      if(_zz_54)begin
        img_reg_array_52_51_imag <= _zz_169;
      end
      if(_zz_55)begin
        img_reg_array_53_51_imag <= _zz_169;
      end
      if(_zz_56)begin
        img_reg_array_54_51_imag <= _zz_169;
      end
      if(_zz_57)begin
        img_reg_array_55_51_imag <= _zz_169;
      end
      if(_zz_58)begin
        img_reg_array_56_51_imag <= _zz_169;
      end
      if(_zz_59)begin
        img_reg_array_57_51_imag <= _zz_169;
      end
      if(_zz_60)begin
        img_reg_array_58_51_imag <= _zz_169;
      end
      if(_zz_61)begin
        img_reg_array_59_51_imag <= _zz_169;
      end
      if(_zz_62)begin
        img_reg_array_60_51_imag <= _zz_169;
      end
      if(_zz_63)begin
        img_reg_array_61_51_imag <= _zz_169;
      end
      if(_zz_64)begin
        img_reg_array_62_51_imag <= _zz_169;
      end
      if(_zz_65)begin
        img_reg_array_63_51_imag <= _zz_169;
      end
      if(_zz_2)begin
        img_reg_array_0_52_real <= _zz_170;
      end
      if(_zz_3)begin
        img_reg_array_1_52_real <= _zz_170;
      end
      if(_zz_4)begin
        img_reg_array_2_52_real <= _zz_170;
      end
      if(_zz_5)begin
        img_reg_array_3_52_real <= _zz_170;
      end
      if(_zz_6)begin
        img_reg_array_4_52_real <= _zz_170;
      end
      if(_zz_7)begin
        img_reg_array_5_52_real <= _zz_170;
      end
      if(_zz_8)begin
        img_reg_array_6_52_real <= _zz_170;
      end
      if(_zz_9)begin
        img_reg_array_7_52_real <= _zz_170;
      end
      if(_zz_10)begin
        img_reg_array_8_52_real <= _zz_170;
      end
      if(_zz_11)begin
        img_reg_array_9_52_real <= _zz_170;
      end
      if(_zz_12)begin
        img_reg_array_10_52_real <= _zz_170;
      end
      if(_zz_13)begin
        img_reg_array_11_52_real <= _zz_170;
      end
      if(_zz_14)begin
        img_reg_array_12_52_real <= _zz_170;
      end
      if(_zz_15)begin
        img_reg_array_13_52_real <= _zz_170;
      end
      if(_zz_16)begin
        img_reg_array_14_52_real <= _zz_170;
      end
      if(_zz_17)begin
        img_reg_array_15_52_real <= _zz_170;
      end
      if(_zz_18)begin
        img_reg_array_16_52_real <= _zz_170;
      end
      if(_zz_19)begin
        img_reg_array_17_52_real <= _zz_170;
      end
      if(_zz_20)begin
        img_reg_array_18_52_real <= _zz_170;
      end
      if(_zz_21)begin
        img_reg_array_19_52_real <= _zz_170;
      end
      if(_zz_22)begin
        img_reg_array_20_52_real <= _zz_170;
      end
      if(_zz_23)begin
        img_reg_array_21_52_real <= _zz_170;
      end
      if(_zz_24)begin
        img_reg_array_22_52_real <= _zz_170;
      end
      if(_zz_25)begin
        img_reg_array_23_52_real <= _zz_170;
      end
      if(_zz_26)begin
        img_reg_array_24_52_real <= _zz_170;
      end
      if(_zz_27)begin
        img_reg_array_25_52_real <= _zz_170;
      end
      if(_zz_28)begin
        img_reg_array_26_52_real <= _zz_170;
      end
      if(_zz_29)begin
        img_reg_array_27_52_real <= _zz_170;
      end
      if(_zz_30)begin
        img_reg_array_28_52_real <= _zz_170;
      end
      if(_zz_31)begin
        img_reg_array_29_52_real <= _zz_170;
      end
      if(_zz_32)begin
        img_reg_array_30_52_real <= _zz_170;
      end
      if(_zz_33)begin
        img_reg_array_31_52_real <= _zz_170;
      end
      if(_zz_34)begin
        img_reg_array_32_52_real <= _zz_170;
      end
      if(_zz_35)begin
        img_reg_array_33_52_real <= _zz_170;
      end
      if(_zz_36)begin
        img_reg_array_34_52_real <= _zz_170;
      end
      if(_zz_37)begin
        img_reg_array_35_52_real <= _zz_170;
      end
      if(_zz_38)begin
        img_reg_array_36_52_real <= _zz_170;
      end
      if(_zz_39)begin
        img_reg_array_37_52_real <= _zz_170;
      end
      if(_zz_40)begin
        img_reg_array_38_52_real <= _zz_170;
      end
      if(_zz_41)begin
        img_reg_array_39_52_real <= _zz_170;
      end
      if(_zz_42)begin
        img_reg_array_40_52_real <= _zz_170;
      end
      if(_zz_43)begin
        img_reg_array_41_52_real <= _zz_170;
      end
      if(_zz_44)begin
        img_reg_array_42_52_real <= _zz_170;
      end
      if(_zz_45)begin
        img_reg_array_43_52_real <= _zz_170;
      end
      if(_zz_46)begin
        img_reg_array_44_52_real <= _zz_170;
      end
      if(_zz_47)begin
        img_reg_array_45_52_real <= _zz_170;
      end
      if(_zz_48)begin
        img_reg_array_46_52_real <= _zz_170;
      end
      if(_zz_49)begin
        img_reg_array_47_52_real <= _zz_170;
      end
      if(_zz_50)begin
        img_reg_array_48_52_real <= _zz_170;
      end
      if(_zz_51)begin
        img_reg_array_49_52_real <= _zz_170;
      end
      if(_zz_52)begin
        img_reg_array_50_52_real <= _zz_170;
      end
      if(_zz_53)begin
        img_reg_array_51_52_real <= _zz_170;
      end
      if(_zz_54)begin
        img_reg_array_52_52_real <= _zz_170;
      end
      if(_zz_55)begin
        img_reg_array_53_52_real <= _zz_170;
      end
      if(_zz_56)begin
        img_reg_array_54_52_real <= _zz_170;
      end
      if(_zz_57)begin
        img_reg_array_55_52_real <= _zz_170;
      end
      if(_zz_58)begin
        img_reg_array_56_52_real <= _zz_170;
      end
      if(_zz_59)begin
        img_reg_array_57_52_real <= _zz_170;
      end
      if(_zz_60)begin
        img_reg_array_58_52_real <= _zz_170;
      end
      if(_zz_61)begin
        img_reg_array_59_52_real <= _zz_170;
      end
      if(_zz_62)begin
        img_reg_array_60_52_real <= _zz_170;
      end
      if(_zz_63)begin
        img_reg_array_61_52_real <= _zz_170;
      end
      if(_zz_64)begin
        img_reg_array_62_52_real <= _zz_170;
      end
      if(_zz_65)begin
        img_reg_array_63_52_real <= _zz_170;
      end
      if(_zz_2)begin
        img_reg_array_0_52_imag <= _zz_171;
      end
      if(_zz_3)begin
        img_reg_array_1_52_imag <= _zz_171;
      end
      if(_zz_4)begin
        img_reg_array_2_52_imag <= _zz_171;
      end
      if(_zz_5)begin
        img_reg_array_3_52_imag <= _zz_171;
      end
      if(_zz_6)begin
        img_reg_array_4_52_imag <= _zz_171;
      end
      if(_zz_7)begin
        img_reg_array_5_52_imag <= _zz_171;
      end
      if(_zz_8)begin
        img_reg_array_6_52_imag <= _zz_171;
      end
      if(_zz_9)begin
        img_reg_array_7_52_imag <= _zz_171;
      end
      if(_zz_10)begin
        img_reg_array_8_52_imag <= _zz_171;
      end
      if(_zz_11)begin
        img_reg_array_9_52_imag <= _zz_171;
      end
      if(_zz_12)begin
        img_reg_array_10_52_imag <= _zz_171;
      end
      if(_zz_13)begin
        img_reg_array_11_52_imag <= _zz_171;
      end
      if(_zz_14)begin
        img_reg_array_12_52_imag <= _zz_171;
      end
      if(_zz_15)begin
        img_reg_array_13_52_imag <= _zz_171;
      end
      if(_zz_16)begin
        img_reg_array_14_52_imag <= _zz_171;
      end
      if(_zz_17)begin
        img_reg_array_15_52_imag <= _zz_171;
      end
      if(_zz_18)begin
        img_reg_array_16_52_imag <= _zz_171;
      end
      if(_zz_19)begin
        img_reg_array_17_52_imag <= _zz_171;
      end
      if(_zz_20)begin
        img_reg_array_18_52_imag <= _zz_171;
      end
      if(_zz_21)begin
        img_reg_array_19_52_imag <= _zz_171;
      end
      if(_zz_22)begin
        img_reg_array_20_52_imag <= _zz_171;
      end
      if(_zz_23)begin
        img_reg_array_21_52_imag <= _zz_171;
      end
      if(_zz_24)begin
        img_reg_array_22_52_imag <= _zz_171;
      end
      if(_zz_25)begin
        img_reg_array_23_52_imag <= _zz_171;
      end
      if(_zz_26)begin
        img_reg_array_24_52_imag <= _zz_171;
      end
      if(_zz_27)begin
        img_reg_array_25_52_imag <= _zz_171;
      end
      if(_zz_28)begin
        img_reg_array_26_52_imag <= _zz_171;
      end
      if(_zz_29)begin
        img_reg_array_27_52_imag <= _zz_171;
      end
      if(_zz_30)begin
        img_reg_array_28_52_imag <= _zz_171;
      end
      if(_zz_31)begin
        img_reg_array_29_52_imag <= _zz_171;
      end
      if(_zz_32)begin
        img_reg_array_30_52_imag <= _zz_171;
      end
      if(_zz_33)begin
        img_reg_array_31_52_imag <= _zz_171;
      end
      if(_zz_34)begin
        img_reg_array_32_52_imag <= _zz_171;
      end
      if(_zz_35)begin
        img_reg_array_33_52_imag <= _zz_171;
      end
      if(_zz_36)begin
        img_reg_array_34_52_imag <= _zz_171;
      end
      if(_zz_37)begin
        img_reg_array_35_52_imag <= _zz_171;
      end
      if(_zz_38)begin
        img_reg_array_36_52_imag <= _zz_171;
      end
      if(_zz_39)begin
        img_reg_array_37_52_imag <= _zz_171;
      end
      if(_zz_40)begin
        img_reg_array_38_52_imag <= _zz_171;
      end
      if(_zz_41)begin
        img_reg_array_39_52_imag <= _zz_171;
      end
      if(_zz_42)begin
        img_reg_array_40_52_imag <= _zz_171;
      end
      if(_zz_43)begin
        img_reg_array_41_52_imag <= _zz_171;
      end
      if(_zz_44)begin
        img_reg_array_42_52_imag <= _zz_171;
      end
      if(_zz_45)begin
        img_reg_array_43_52_imag <= _zz_171;
      end
      if(_zz_46)begin
        img_reg_array_44_52_imag <= _zz_171;
      end
      if(_zz_47)begin
        img_reg_array_45_52_imag <= _zz_171;
      end
      if(_zz_48)begin
        img_reg_array_46_52_imag <= _zz_171;
      end
      if(_zz_49)begin
        img_reg_array_47_52_imag <= _zz_171;
      end
      if(_zz_50)begin
        img_reg_array_48_52_imag <= _zz_171;
      end
      if(_zz_51)begin
        img_reg_array_49_52_imag <= _zz_171;
      end
      if(_zz_52)begin
        img_reg_array_50_52_imag <= _zz_171;
      end
      if(_zz_53)begin
        img_reg_array_51_52_imag <= _zz_171;
      end
      if(_zz_54)begin
        img_reg_array_52_52_imag <= _zz_171;
      end
      if(_zz_55)begin
        img_reg_array_53_52_imag <= _zz_171;
      end
      if(_zz_56)begin
        img_reg_array_54_52_imag <= _zz_171;
      end
      if(_zz_57)begin
        img_reg_array_55_52_imag <= _zz_171;
      end
      if(_zz_58)begin
        img_reg_array_56_52_imag <= _zz_171;
      end
      if(_zz_59)begin
        img_reg_array_57_52_imag <= _zz_171;
      end
      if(_zz_60)begin
        img_reg_array_58_52_imag <= _zz_171;
      end
      if(_zz_61)begin
        img_reg_array_59_52_imag <= _zz_171;
      end
      if(_zz_62)begin
        img_reg_array_60_52_imag <= _zz_171;
      end
      if(_zz_63)begin
        img_reg_array_61_52_imag <= _zz_171;
      end
      if(_zz_64)begin
        img_reg_array_62_52_imag <= _zz_171;
      end
      if(_zz_65)begin
        img_reg_array_63_52_imag <= _zz_171;
      end
      if(_zz_2)begin
        img_reg_array_0_53_real <= _zz_172;
      end
      if(_zz_3)begin
        img_reg_array_1_53_real <= _zz_172;
      end
      if(_zz_4)begin
        img_reg_array_2_53_real <= _zz_172;
      end
      if(_zz_5)begin
        img_reg_array_3_53_real <= _zz_172;
      end
      if(_zz_6)begin
        img_reg_array_4_53_real <= _zz_172;
      end
      if(_zz_7)begin
        img_reg_array_5_53_real <= _zz_172;
      end
      if(_zz_8)begin
        img_reg_array_6_53_real <= _zz_172;
      end
      if(_zz_9)begin
        img_reg_array_7_53_real <= _zz_172;
      end
      if(_zz_10)begin
        img_reg_array_8_53_real <= _zz_172;
      end
      if(_zz_11)begin
        img_reg_array_9_53_real <= _zz_172;
      end
      if(_zz_12)begin
        img_reg_array_10_53_real <= _zz_172;
      end
      if(_zz_13)begin
        img_reg_array_11_53_real <= _zz_172;
      end
      if(_zz_14)begin
        img_reg_array_12_53_real <= _zz_172;
      end
      if(_zz_15)begin
        img_reg_array_13_53_real <= _zz_172;
      end
      if(_zz_16)begin
        img_reg_array_14_53_real <= _zz_172;
      end
      if(_zz_17)begin
        img_reg_array_15_53_real <= _zz_172;
      end
      if(_zz_18)begin
        img_reg_array_16_53_real <= _zz_172;
      end
      if(_zz_19)begin
        img_reg_array_17_53_real <= _zz_172;
      end
      if(_zz_20)begin
        img_reg_array_18_53_real <= _zz_172;
      end
      if(_zz_21)begin
        img_reg_array_19_53_real <= _zz_172;
      end
      if(_zz_22)begin
        img_reg_array_20_53_real <= _zz_172;
      end
      if(_zz_23)begin
        img_reg_array_21_53_real <= _zz_172;
      end
      if(_zz_24)begin
        img_reg_array_22_53_real <= _zz_172;
      end
      if(_zz_25)begin
        img_reg_array_23_53_real <= _zz_172;
      end
      if(_zz_26)begin
        img_reg_array_24_53_real <= _zz_172;
      end
      if(_zz_27)begin
        img_reg_array_25_53_real <= _zz_172;
      end
      if(_zz_28)begin
        img_reg_array_26_53_real <= _zz_172;
      end
      if(_zz_29)begin
        img_reg_array_27_53_real <= _zz_172;
      end
      if(_zz_30)begin
        img_reg_array_28_53_real <= _zz_172;
      end
      if(_zz_31)begin
        img_reg_array_29_53_real <= _zz_172;
      end
      if(_zz_32)begin
        img_reg_array_30_53_real <= _zz_172;
      end
      if(_zz_33)begin
        img_reg_array_31_53_real <= _zz_172;
      end
      if(_zz_34)begin
        img_reg_array_32_53_real <= _zz_172;
      end
      if(_zz_35)begin
        img_reg_array_33_53_real <= _zz_172;
      end
      if(_zz_36)begin
        img_reg_array_34_53_real <= _zz_172;
      end
      if(_zz_37)begin
        img_reg_array_35_53_real <= _zz_172;
      end
      if(_zz_38)begin
        img_reg_array_36_53_real <= _zz_172;
      end
      if(_zz_39)begin
        img_reg_array_37_53_real <= _zz_172;
      end
      if(_zz_40)begin
        img_reg_array_38_53_real <= _zz_172;
      end
      if(_zz_41)begin
        img_reg_array_39_53_real <= _zz_172;
      end
      if(_zz_42)begin
        img_reg_array_40_53_real <= _zz_172;
      end
      if(_zz_43)begin
        img_reg_array_41_53_real <= _zz_172;
      end
      if(_zz_44)begin
        img_reg_array_42_53_real <= _zz_172;
      end
      if(_zz_45)begin
        img_reg_array_43_53_real <= _zz_172;
      end
      if(_zz_46)begin
        img_reg_array_44_53_real <= _zz_172;
      end
      if(_zz_47)begin
        img_reg_array_45_53_real <= _zz_172;
      end
      if(_zz_48)begin
        img_reg_array_46_53_real <= _zz_172;
      end
      if(_zz_49)begin
        img_reg_array_47_53_real <= _zz_172;
      end
      if(_zz_50)begin
        img_reg_array_48_53_real <= _zz_172;
      end
      if(_zz_51)begin
        img_reg_array_49_53_real <= _zz_172;
      end
      if(_zz_52)begin
        img_reg_array_50_53_real <= _zz_172;
      end
      if(_zz_53)begin
        img_reg_array_51_53_real <= _zz_172;
      end
      if(_zz_54)begin
        img_reg_array_52_53_real <= _zz_172;
      end
      if(_zz_55)begin
        img_reg_array_53_53_real <= _zz_172;
      end
      if(_zz_56)begin
        img_reg_array_54_53_real <= _zz_172;
      end
      if(_zz_57)begin
        img_reg_array_55_53_real <= _zz_172;
      end
      if(_zz_58)begin
        img_reg_array_56_53_real <= _zz_172;
      end
      if(_zz_59)begin
        img_reg_array_57_53_real <= _zz_172;
      end
      if(_zz_60)begin
        img_reg_array_58_53_real <= _zz_172;
      end
      if(_zz_61)begin
        img_reg_array_59_53_real <= _zz_172;
      end
      if(_zz_62)begin
        img_reg_array_60_53_real <= _zz_172;
      end
      if(_zz_63)begin
        img_reg_array_61_53_real <= _zz_172;
      end
      if(_zz_64)begin
        img_reg_array_62_53_real <= _zz_172;
      end
      if(_zz_65)begin
        img_reg_array_63_53_real <= _zz_172;
      end
      if(_zz_2)begin
        img_reg_array_0_53_imag <= _zz_173;
      end
      if(_zz_3)begin
        img_reg_array_1_53_imag <= _zz_173;
      end
      if(_zz_4)begin
        img_reg_array_2_53_imag <= _zz_173;
      end
      if(_zz_5)begin
        img_reg_array_3_53_imag <= _zz_173;
      end
      if(_zz_6)begin
        img_reg_array_4_53_imag <= _zz_173;
      end
      if(_zz_7)begin
        img_reg_array_5_53_imag <= _zz_173;
      end
      if(_zz_8)begin
        img_reg_array_6_53_imag <= _zz_173;
      end
      if(_zz_9)begin
        img_reg_array_7_53_imag <= _zz_173;
      end
      if(_zz_10)begin
        img_reg_array_8_53_imag <= _zz_173;
      end
      if(_zz_11)begin
        img_reg_array_9_53_imag <= _zz_173;
      end
      if(_zz_12)begin
        img_reg_array_10_53_imag <= _zz_173;
      end
      if(_zz_13)begin
        img_reg_array_11_53_imag <= _zz_173;
      end
      if(_zz_14)begin
        img_reg_array_12_53_imag <= _zz_173;
      end
      if(_zz_15)begin
        img_reg_array_13_53_imag <= _zz_173;
      end
      if(_zz_16)begin
        img_reg_array_14_53_imag <= _zz_173;
      end
      if(_zz_17)begin
        img_reg_array_15_53_imag <= _zz_173;
      end
      if(_zz_18)begin
        img_reg_array_16_53_imag <= _zz_173;
      end
      if(_zz_19)begin
        img_reg_array_17_53_imag <= _zz_173;
      end
      if(_zz_20)begin
        img_reg_array_18_53_imag <= _zz_173;
      end
      if(_zz_21)begin
        img_reg_array_19_53_imag <= _zz_173;
      end
      if(_zz_22)begin
        img_reg_array_20_53_imag <= _zz_173;
      end
      if(_zz_23)begin
        img_reg_array_21_53_imag <= _zz_173;
      end
      if(_zz_24)begin
        img_reg_array_22_53_imag <= _zz_173;
      end
      if(_zz_25)begin
        img_reg_array_23_53_imag <= _zz_173;
      end
      if(_zz_26)begin
        img_reg_array_24_53_imag <= _zz_173;
      end
      if(_zz_27)begin
        img_reg_array_25_53_imag <= _zz_173;
      end
      if(_zz_28)begin
        img_reg_array_26_53_imag <= _zz_173;
      end
      if(_zz_29)begin
        img_reg_array_27_53_imag <= _zz_173;
      end
      if(_zz_30)begin
        img_reg_array_28_53_imag <= _zz_173;
      end
      if(_zz_31)begin
        img_reg_array_29_53_imag <= _zz_173;
      end
      if(_zz_32)begin
        img_reg_array_30_53_imag <= _zz_173;
      end
      if(_zz_33)begin
        img_reg_array_31_53_imag <= _zz_173;
      end
      if(_zz_34)begin
        img_reg_array_32_53_imag <= _zz_173;
      end
      if(_zz_35)begin
        img_reg_array_33_53_imag <= _zz_173;
      end
      if(_zz_36)begin
        img_reg_array_34_53_imag <= _zz_173;
      end
      if(_zz_37)begin
        img_reg_array_35_53_imag <= _zz_173;
      end
      if(_zz_38)begin
        img_reg_array_36_53_imag <= _zz_173;
      end
      if(_zz_39)begin
        img_reg_array_37_53_imag <= _zz_173;
      end
      if(_zz_40)begin
        img_reg_array_38_53_imag <= _zz_173;
      end
      if(_zz_41)begin
        img_reg_array_39_53_imag <= _zz_173;
      end
      if(_zz_42)begin
        img_reg_array_40_53_imag <= _zz_173;
      end
      if(_zz_43)begin
        img_reg_array_41_53_imag <= _zz_173;
      end
      if(_zz_44)begin
        img_reg_array_42_53_imag <= _zz_173;
      end
      if(_zz_45)begin
        img_reg_array_43_53_imag <= _zz_173;
      end
      if(_zz_46)begin
        img_reg_array_44_53_imag <= _zz_173;
      end
      if(_zz_47)begin
        img_reg_array_45_53_imag <= _zz_173;
      end
      if(_zz_48)begin
        img_reg_array_46_53_imag <= _zz_173;
      end
      if(_zz_49)begin
        img_reg_array_47_53_imag <= _zz_173;
      end
      if(_zz_50)begin
        img_reg_array_48_53_imag <= _zz_173;
      end
      if(_zz_51)begin
        img_reg_array_49_53_imag <= _zz_173;
      end
      if(_zz_52)begin
        img_reg_array_50_53_imag <= _zz_173;
      end
      if(_zz_53)begin
        img_reg_array_51_53_imag <= _zz_173;
      end
      if(_zz_54)begin
        img_reg_array_52_53_imag <= _zz_173;
      end
      if(_zz_55)begin
        img_reg_array_53_53_imag <= _zz_173;
      end
      if(_zz_56)begin
        img_reg_array_54_53_imag <= _zz_173;
      end
      if(_zz_57)begin
        img_reg_array_55_53_imag <= _zz_173;
      end
      if(_zz_58)begin
        img_reg_array_56_53_imag <= _zz_173;
      end
      if(_zz_59)begin
        img_reg_array_57_53_imag <= _zz_173;
      end
      if(_zz_60)begin
        img_reg_array_58_53_imag <= _zz_173;
      end
      if(_zz_61)begin
        img_reg_array_59_53_imag <= _zz_173;
      end
      if(_zz_62)begin
        img_reg_array_60_53_imag <= _zz_173;
      end
      if(_zz_63)begin
        img_reg_array_61_53_imag <= _zz_173;
      end
      if(_zz_64)begin
        img_reg_array_62_53_imag <= _zz_173;
      end
      if(_zz_65)begin
        img_reg_array_63_53_imag <= _zz_173;
      end
      if(_zz_2)begin
        img_reg_array_0_54_real <= _zz_174;
      end
      if(_zz_3)begin
        img_reg_array_1_54_real <= _zz_174;
      end
      if(_zz_4)begin
        img_reg_array_2_54_real <= _zz_174;
      end
      if(_zz_5)begin
        img_reg_array_3_54_real <= _zz_174;
      end
      if(_zz_6)begin
        img_reg_array_4_54_real <= _zz_174;
      end
      if(_zz_7)begin
        img_reg_array_5_54_real <= _zz_174;
      end
      if(_zz_8)begin
        img_reg_array_6_54_real <= _zz_174;
      end
      if(_zz_9)begin
        img_reg_array_7_54_real <= _zz_174;
      end
      if(_zz_10)begin
        img_reg_array_8_54_real <= _zz_174;
      end
      if(_zz_11)begin
        img_reg_array_9_54_real <= _zz_174;
      end
      if(_zz_12)begin
        img_reg_array_10_54_real <= _zz_174;
      end
      if(_zz_13)begin
        img_reg_array_11_54_real <= _zz_174;
      end
      if(_zz_14)begin
        img_reg_array_12_54_real <= _zz_174;
      end
      if(_zz_15)begin
        img_reg_array_13_54_real <= _zz_174;
      end
      if(_zz_16)begin
        img_reg_array_14_54_real <= _zz_174;
      end
      if(_zz_17)begin
        img_reg_array_15_54_real <= _zz_174;
      end
      if(_zz_18)begin
        img_reg_array_16_54_real <= _zz_174;
      end
      if(_zz_19)begin
        img_reg_array_17_54_real <= _zz_174;
      end
      if(_zz_20)begin
        img_reg_array_18_54_real <= _zz_174;
      end
      if(_zz_21)begin
        img_reg_array_19_54_real <= _zz_174;
      end
      if(_zz_22)begin
        img_reg_array_20_54_real <= _zz_174;
      end
      if(_zz_23)begin
        img_reg_array_21_54_real <= _zz_174;
      end
      if(_zz_24)begin
        img_reg_array_22_54_real <= _zz_174;
      end
      if(_zz_25)begin
        img_reg_array_23_54_real <= _zz_174;
      end
      if(_zz_26)begin
        img_reg_array_24_54_real <= _zz_174;
      end
      if(_zz_27)begin
        img_reg_array_25_54_real <= _zz_174;
      end
      if(_zz_28)begin
        img_reg_array_26_54_real <= _zz_174;
      end
      if(_zz_29)begin
        img_reg_array_27_54_real <= _zz_174;
      end
      if(_zz_30)begin
        img_reg_array_28_54_real <= _zz_174;
      end
      if(_zz_31)begin
        img_reg_array_29_54_real <= _zz_174;
      end
      if(_zz_32)begin
        img_reg_array_30_54_real <= _zz_174;
      end
      if(_zz_33)begin
        img_reg_array_31_54_real <= _zz_174;
      end
      if(_zz_34)begin
        img_reg_array_32_54_real <= _zz_174;
      end
      if(_zz_35)begin
        img_reg_array_33_54_real <= _zz_174;
      end
      if(_zz_36)begin
        img_reg_array_34_54_real <= _zz_174;
      end
      if(_zz_37)begin
        img_reg_array_35_54_real <= _zz_174;
      end
      if(_zz_38)begin
        img_reg_array_36_54_real <= _zz_174;
      end
      if(_zz_39)begin
        img_reg_array_37_54_real <= _zz_174;
      end
      if(_zz_40)begin
        img_reg_array_38_54_real <= _zz_174;
      end
      if(_zz_41)begin
        img_reg_array_39_54_real <= _zz_174;
      end
      if(_zz_42)begin
        img_reg_array_40_54_real <= _zz_174;
      end
      if(_zz_43)begin
        img_reg_array_41_54_real <= _zz_174;
      end
      if(_zz_44)begin
        img_reg_array_42_54_real <= _zz_174;
      end
      if(_zz_45)begin
        img_reg_array_43_54_real <= _zz_174;
      end
      if(_zz_46)begin
        img_reg_array_44_54_real <= _zz_174;
      end
      if(_zz_47)begin
        img_reg_array_45_54_real <= _zz_174;
      end
      if(_zz_48)begin
        img_reg_array_46_54_real <= _zz_174;
      end
      if(_zz_49)begin
        img_reg_array_47_54_real <= _zz_174;
      end
      if(_zz_50)begin
        img_reg_array_48_54_real <= _zz_174;
      end
      if(_zz_51)begin
        img_reg_array_49_54_real <= _zz_174;
      end
      if(_zz_52)begin
        img_reg_array_50_54_real <= _zz_174;
      end
      if(_zz_53)begin
        img_reg_array_51_54_real <= _zz_174;
      end
      if(_zz_54)begin
        img_reg_array_52_54_real <= _zz_174;
      end
      if(_zz_55)begin
        img_reg_array_53_54_real <= _zz_174;
      end
      if(_zz_56)begin
        img_reg_array_54_54_real <= _zz_174;
      end
      if(_zz_57)begin
        img_reg_array_55_54_real <= _zz_174;
      end
      if(_zz_58)begin
        img_reg_array_56_54_real <= _zz_174;
      end
      if(_zz_59)begin
        img_reg_array_57_54_real <= _zz_174;
      end
      if(_zz_60)begin
        img_reg_array_58_54_real <= _zz_174;
      end
      if(_zz_61)begin
        img_reg_array_59_54_real <= _zz_174;
      end
      if(_zz_62)begin
        img_reg_array_60_54_real <= _zz_174;
      end
      if(_zz_63)begin
        img_reg_array_61_54_real <= _zz_174;
      end
      if(_zz_64)begin
        img_reg_array_62_54_real <= _zz_174;
      end
      if(_zz_65)begin
        img_reg_array_63_54_real <= _zz_174;
      end
      if(_zz_2)begin
        img_reg_array_0_54_imag <= _zz_175;
      end
      if(_zz_3)begin
        img_reg_array_1_54_imag <= _zz_175;
      end
      if(_zz_4)begin
        img_reg_array_2_54_imag <= _zz_175;
      end
      if(_zz_5)begin
        img_reg_array_3_54_imag <= _zz_175;
      end
      if(_zz_6)begin
        img_reg_array_4_54_imag <= _zz_175;
      end
      if(_zz_7)begin
        img_reg_array_5_54_imag <= _zz_175;
      end
      if(_zz_8)begin
        img_reg_array_6_54_imag <= _zz_175;
      end
      if(_zz_9)begin
        img_reg_array_7_54_imag <= _zz_175;
      end
      if(_zz_10)begin
        img_reg_array_8_54_imag <= _zz_175;
      end
      if(_zz_11)begin
        img_reg_array_9_54_imag <= _zz_175;
      end
      if(_zz_12)begin
        img_reg_array_10_54_imag <= _zz_175;
      end
      if(_zz_13)begin
        img_reg_array_11_54_imag <= _zz_175;
      end
      if(_zz_14)begin
        img_reg_array_12_54_imag <= _zz_175;
      end
      if(_zz_15)begin
        img_reg_array_13_54_imag <= _zz_175;
      end
      if(_zz_16)begin
        img_reg_array_14_54_imag <= _zz_175;
      end
      if(_zz_17)begin
        img_reg_array_15_54_imag <= _zz_175;
      end
      if(_zz_18)begin
        img_reg_array_16_54_imag <= _zz_175;
      end
      if(_zz_19)begin
        img_reg_array_17_54_imag <= _zz_175;
      end
      if(_zz_20)begin
        img_reg_array_18_54_imag <= _zz_175;
      end
      if(_zz_21)begin
        img_reg_array_19_54_imag <= _zz_175;
      end
      if(_zz_22)begin
        img_reg_array_20_54_imag <= _zz_175;
      end
      if(_zz_23)begin
        img_reg_array_21_54_imag <= _zz_175;
      end
      if(_zz_24)begin
        img_reg_array_22_54_imag <= _zz_175;
      end
      if(_zz_25)begin
        img_reg_array_23_54_imag <= _zz_175;
      end
      if(_zz_26)begin
        img_reg_array_24_54_imag <= _zz_175;
      end
      if(_zz_27)begin
        img_reg_array_25_54_imag <= _zz_175;
      end
      if(_zz_28)begin
        img_reg_array_26_54_imag <= _zz_175;
      end
      if(_zz_29)begin
        img_reg_array_27_54_imag <= _zz_175;
      end
      if(_zz_30)begin
        img_reg_array_28_54_imag <= _zz_175;
      end
      if(_zz_31)begin
        img_reg_array_29_54_imag <= _zz_175;
      end
      if(_zz_32)begin
        img_reg_array_30_54_imag <= _zz_175;
      end
      if(_zz_33)begin
        img_reg_array_31_54_imag <= _zz_175;
      end
      if(_zz_34)begin
        img_reg_array_32_54_imag <= _zz_175;
      end
      if(_zz_35)begin
        img_reg_array_33_54_imag <= _zz_175;
      end
      if(_zz_36)begin
        img_reg_array_34_54_imag <= _zz_175;
      end
      if(_zz_37)begin
        img_reg_array_35_54_imag <= _zz_175;
      end
      if(_zz_38)begin
        img_reg_array_36_54_imag <= _zz_175;
      end
      if(_zz_39)begin
        img_reg_array_37_54_imag <= _zz_175;
      end
      if(_zz_40)begin
        img_reg_array_38_54_imag <= _zz_175;
      end
      if(_zz_41)begin
        img_reg_array_39_54_imag <= _zz_175;
      end
      if(_zz_42)begin
        img_reg_array_40_54_imag <= _zz_175;
      end
      if(_zz_43)begin
        img_reg_array_41_54_imag <= _zz_175;
      end
      if(_zz_44)begin
        img_reg_array_42_54_imag <= _zz_175;
      end
      if(_zz_45)begin
        img_reg_array_43_54_imag <= _zz_175;
      end
      if(_zz_46)begin
        img_reg_array_44_54_imag <= _zz_175;
      end
      if(_zz_47)begin
        img_reg_array_45_54_imag <= _zz_175;
      end
      if(_zz_48)begin
        img_reg_array_46_54_imag <= _zz_175;
      end
      if(_zz_49)begin
        img_reg_array_47_54_imag <= _zz_175;
      end
      if(_zz_50)begin
        img_reg_array_48_54_imag <= _zz_175;
      end
      if(_zz_51)begin
        img_reg_array_49_54_imag <= _zz_175;
      end
      if(_zz_52)begin
        img_reg_array_50_54_imag <= _zz_175;
      end
      if(_zz_53)begin
        img_reg_array_51_54_imag <= _zz_175;
      end
      if(_zz_54)begin
        img_reg_array_52_54_imag <= _zz_175;
      end
      if(_zz_55)begin
        img_reg_array_53_54_imag <= _zz_175;
      end
      if(_zz_56)begin
        img_reg_array_54_54_imag <= _zz_175;
      end
      if(_zz_57)begin
        img_reg_array_55_54_imag <= _zz_175;
      end
      if(_zz_58)begin
        img_reg_array_56_54_imag <= _zz_175;
      end
      if(_zz_59)begin
        img_reg_array_57_54_imag <= _zz_175;
      end
      if(_zz_60)begin
        img_reg_array_58_54_imag <= _zz_175;
      end
      if(_zz_61)begin
        img_reg_array_59_54_imag <= _zz_175;
      end
      if(_zz_62)begin
        img_reg_array_60_54_imag <= _zz_175;
      end
      if(_zz_63)begin
        img_reg_array_61_54_imag <= _zz_175;
      end
      if(_zz_64)begin
        img_reg_array_62_54_imag <= _zz_175;
      end
      if(_zz_65)begin
        img_reg_array_63_54_imag <= _zz_175;
      end
      if(_zz_2)begin
        img_reg_array_0_55_real <= _zz_176;
      end
      if(_zz_3)begin
        img_reg_array_1_55_real <= _zz_176;
      end
      if(_zz_4)begin
        img_reg_array_2_55_real <= _zz_176;
      end
      if(_zz_5)begin
        img_reg_array_3_55_real <= _zz_176;
      end
      if(_zz_6)begin
        img_reg_array_4_55_real <= _zz_176;
      end
      if(_zz_7)begin
        img_reg_array_5_55_real <= _zz_176;
      end
      if(_zz_8)begin
        img_reg_array_6_55_real <= _zz_176;
      end
      if(_zz_9)begin
        img_reg_array_7_55_real <= _zz_176;
      end
      if(_zz_10)begin
        img_reg_array_8_55_real <= _zz_176;
      end
      if(_zz_11)begin
        img_reg_array_9_55_real <= _zz_176;
      end
      if(_zz_12)begin
        img_reg_array_10_55_real <= _zz_176;
      end
      if(_zz_13)begin
        img_reg_array_11_55_real <= _zz_176;
      end
      if(_zz_14)begin
        img_reg_array_12_55_real <= _zz_176;
      end
      if(_zz_15)begin
        img_reg_array_13_55_real <= _zz_176;
      end
      if(_zz_16)begin
        img_reg_array_14_55_real <= _zz_176;
      end
      if(_zz_17)begin
        img_reg_array_15_55_real <= _zz_176;
      end
      if(_zz_18)begin
        img_reg_array_16_55_real <= _zz_176;
      end
      if(_zz_19)begin
        img_reg_array_17_55_real <= _zz_176;
      end
      if(_zz_20)begin
        img_reg_array_18_55_real <= _zz_176;
      end
      if(_zz_21)begin
        img_reg_array_19_55_real <= _zz_176;
      end
      if(_zz_22)begin
        img_reg_array_20_55_real <= _zz_176;
      end
      if(_zz_23)begin
        img_reg_array_21_55_real <= _zz_176;
      end
      if(_zz_24)begin
        img_reg_array_22_55_real <= _zz_176;
      end
      if(_zz_25)begin
        img_reg_array_23_55_real <= _zz_176;
      end
      if(_zz_26)begin
        img_reg_array_24_55_real <= _zz_176;
      end
      if(_zz_27)begin
        img_reg_array_25_55_real <= _zz_176;
      end
      if(_zz_28)begin
        img_reg_array_26_55_real <= _zz_176;
      end
      if(_zz_29)begin
        img_reg_array_27_55_real <= _zz_176;
      end
      if(_zz_30)begin
        img_reg_array_28_55_real <= _zz_176;
      end
      if(_zz_31)begin
        img_reg_array_29_55_real <= _zz_176;
      end
      if(_zz_32)begin
        img_reg_array_30_55_real <= _zz_176;
      end
      if(_zz_33)begin
        img_reg_array_31_55_real <= _zz_176;
      end
      if(_zz_34)begin
        img_reg_array_32_55_real <= _zz_176;
      end
      if(_zz_35)begin
        img_reg_array_33_55_real <= _zz_176;
      end
      if(_zz_36)begin
        img_reg_array_34_55_real <= _zz_176;
      end
      if(_zz_37)begin
        img_reg_array_35_55_real <= _zz_176;
      end
      if(_zz_38)begin
        img_reg_array_36_55_real <= _zz_176;
      end
      if(_zz_39)begin
        img_reg_array_37_55_real <= _zz_176;
      end
      if(_zz_40)begin
        img_reg_array_38_55_real <= _zz_176;
      end
      if(_zz_41)begin
        img_reg_array_39_55_real <= _zz_176;
      end
      if(_zz_42)begin
        img_reg_array_40_55_real <= _zz_176;
      end
      if(_zz_43)begin
        img_reg_array_41_55_real <= _zz_176;
      end
      if(_zz_44)begin
        img_reg_array_42_55_real <= _zz_176;
      end
      if(_zz_45)begin
        img_reg_array_43_55_real <= _zz_176;
      end
      if(_zz_46)begin
        img_reg_array_44_55_real <= _zz_176;
      end
      if(_zz_47)begin
        img_reg_array_45_55_real <= _zz_176;
      end
      if(_zz_48)begin
        img_reg_array_46_55_real <= _zz_176;
      end
      if(_zz_49)begin
        img_reg_array_47_55_real <= _zz_176;
      end
      if(_zz_50)begin
        img_reg_array_48_55_real <= _zz_176;
      end
      if(_zz_51)begin
        img_reg_array_49_55_real <= _zz_176;
      end
      if(_zz_52)begin
        img_reg_array_50_55_real <= _zz_176;
      end
      if(_zz_53)begin
        img_reg_array_51_55_real <= _zz_176;
      end
      if(_zz_54)begin
        img_reg_array_52_55_real <= _zz_176;
      end
      if(_zz_55)begin
        img_reg_array_53_55_real <= _zz_176;
      end
      if(_zz_56)begin
        img_reg_array_54_55_real <= _zz_176;
      end
      if(_zz_57)begin
        img_reg_array_55_55_real <= _zz_176;
      end
      if(_zz_58)begin
        img_reg_array_56_55_real <= _zz_176;
      end
      if(_zz_59)begin
        img_reg_array_57_55_real <= _zz_176;
      end
      if(_zz_60)begin
        img_reg_array_58_55_real <= _zz_176;
      end
      if(_zz_61)begin
        img_reg_array_59_55_real <= _zz_176;
      end
      if(_zz_62)begin
        img_reg_array_60_55_real <= _zz_176;
      end
      if(_zz_63)begin
        img_reg_array_61_55_real <= _zz_176;
      end
      if(_zz_64)begin
        img_reg_array_62_55_real <= _zz_176;
      end
      if(_zz_65)begin
        img_reg_array_63_55_real <= _zz_176;
      end
      if(_zz_2)begin
        img_reg_array_0_55_imag <= _zz_177;
      end
      if(_zz_3)begin
        img_reg_array_1_55_imag <= _zz_177;
      end
      if(_zz_4)begin
        img_reg_array_2_55_imag <= _zz_177;
      end
      if(_zz_5)begin
        img_reg_array_3_55_imag <= _zz_177;
      end
      if(_zz_6)begin
        img_reg_array_4_55_imag <= _zz_177;
      end
      if(_zz_7)begin
        img_reg_array_5_55_imag <= _zz_177;
      end
      if(_zz_8)begin
        img_reg_array_6_55_imag <= _zz_177;
      end
      if(_zz_9)begin
        img_reg_array_7_55_imag <= _zz_177;
      end
      if(_zz_10)begin
        img_reg_array_8_55_imag <= _zz_177;
      end
      if(_zz_11)begin
        img_reg_array_9_55_imag <= _zz_177;
      end
      if(_zz_12)begin
        img_reg_array_10_55_imag <= _zz_177;
      end
      if(_zz_13)begin
        img_reg_array_11_55_imag <= _zz_177;
      end
      if(_zz_14)begin
        img_reg_array_12_55_imag <= _zz_177;
      end
      if(_zz_15)begin
        img_reg_array_13_55_imag <= _zz_177;
      end
      if(_zz_16)begin
        img_reg_array_14_55_imag <= _zz_177;
      end
      if(_zz_17)begin
        img_reg_array_15_55_imag <= _zz_177;
      end
      if(_zz_18)begin
        img_reg_array_16_55_imag <= _zz_177;
      end
      if(_zz_19)begin
        img_reg_array_17_55_imag <= _zz_177;
      end
      if(_zz_20)begin
        img_reg_array_18_55_imag <= _zz_177;
      end
      if(_zz_21)begin
        img_reg_array_19_55_imag <= _zz_177;
      end
      if(_zz_22)begin
        img_reg_array_20_55_imag <= _zz_177;
      end
      if(_zz_23)begin
        img_reg_array_21_55_imag <= _zz_177;
      end
      if(_zz_24)begin
        img_reg_array_22_55_imag <= _zz_177;
      end
      if(_zz_25)begin
        img_reg_array_23_55_imag <= _zz_177;
      end
      if(_zz_26)begin
        img_reg_array_24_55_imag <= _zz_177;
      end
      if(_zz_27)begin
        img_reg_array_25_55_imag <= _zz_177;
      end
      if(_zz_28)begin
        img_reg_array_26_55_imag <= _zz_177;
      end
      if(_zz_29)begin
        img_reg_array_27_55_imag <= _zz_177;
      end
      if(_zz_30)begin
        img_reg_array_28_55_imag <= _zz_177;
      end
      if(_zz_31)begin
        img_reg_array_29_55_imag <= _zz_177;
      end
      if(_zz_32)begin
        img_reg_array_30_55_imag <= _zz_177;
      end
      if(_zz_33)begin
        img_reg_array_31_55_imag <= _zz_177;
      end
      if(_zz_34)begin
        img_reg_array_32_55_imag <= _zz_177;
      end
      if(_zz_35)begin
        img_reg_array_33_55_imag <= _zz_177;
      end
      if(_zz_36)begin
        img_reg_array_34_55_imag <= _zz_177;
      end
      if(_zz_37)begin
        img_reg_array_35_55_imag <= _zz_177;
      end
      if(_zz_38)begin
        img_reg_array_36_55_imag <= _zz_177;
      end
      if(_zz_39)begin
        img_reg_array_37_55_imag <= _zz_177;
      end
      if(_zz_40)begin
        img_reg_array_38_55_imag <= _zz_177;
      end
      if(_zz_41)begin
        img_reg_array_39_55_imag <= _zz_177;
      end
      if(_zz_42)begin
        img_reg_array_40_55_imag <= _zz_177;
      end
      if(_zz_43)begin
        img_reg_array_41_55_imag <= _zz_177;
      end
      if(_zz_44)begin
        img_reg_array_42_55_imag <= _zz_177;
      end
      if(_zz_45)begin
        img_reg_array_43_55_imag <= _zz_177;
      end
      if(_zz_46)begin
        img_reg_array_44_55_imag <= _zz_177;
      end
      if(_zz_47)begin
        img_reg_array_45_55_imag <= _zz_177;
      end
      if(_zz_48)begin
        img_reg_array_46_55_imag <= _zz_177;
      end
      if(_zz_49)begin
        img_reg_array_47_55_imag <= _zz_177;
      end
      if(_zz_50)begin
        img_reg_array_48_55_imag <= _zz_177;
      end
      if(_zz_51)begin
        img_reg_array_49_55_imag <= _zz_177;
      end
      if(_zz_52)begin
        img_reg_array_50_55_imag <= _zz_177;
      end
      if(_zz_53)begin
        img_reg_array_51_55_imag <= _zz_177;
      end
      if(_zz_54)begin
        img_reg_array_52_55_imag <= _zz_177;
      end
      if(_zz_55)begin
        img_reg_array_53_55_imag <= _zz_177;
      end
      if(_zz_56)begin
        img_reg_array_54_55_imag <= _zz_177;
      end
      if(_zz_57)begin
        img_reg_array_55_55_imag <= _zz_177;
      end
      if(_zz_58)begin
        img_reg_array_56_55_imag <= _zz_177;
      end
      if(_zz_59)begin
        img_reg_array_57_55_imag <= _zz_177;
      end
      if(_zz_60)begin
        img_reg_array_58_55_imag <= _zz_177;
      end
      if(_zz_61)begin
        img_reg_array_59_55_imag <= _zz_177;
      end
      if(_zz_62)begin
        img_reg_array_60_55_imag <= _zz_177;
      end
      if(_zz_63)begin
        img_reg_array_61_55_imag <= _zz_177;
      end
      if(_zz_64)begin
        img_reg_array_62_55_imag <= _zz_177;
      end
      if(_zz_65)begin
        img_reg_array_63_55_imag <= _zz_177;
      end
      if(_zz_2)begin
        img_reg_array_0_56_real <= _zz_178;
      end
      if(_zz_3)begin
        img_reg_array_1_56_real <= _zz_178;
      end
      if(_zz_4)begin
        img_reg_array_2_56_real <= _zz_178;
      end
      if(_zz_5)begin
        img_reg_array_3_56_real <= _zz_178;
      end
      if(_zz_6)begin
        img_reg_array_4_56_real <= _zz_178;
      end
      if(_zz_7)begin
        img_reg_array_5_56_real <= _zz_178;
      end
      if(_zz_8)begin
        img_reg_array_6_56_real <= _zz_178;
      end
      if(_zz_9)begin
        img_reg_array_7_56_real <= _zz_178;
      end
      if(_zz_10)begin
        img_reg_array_8_56_real <= _zz_178;
      end
      if(_zz_11)begin
        img_reg_array_9_56_real <= _zz_178;
      end
      if(_zz_12)begin
        img_reg_array_10_56_real <= _zz_178;
      end
      if(_zz_13)begin
        img_reg_array_11_56_real <= _zz_178;
      end
      if(_zz_14)begin
        img_reg_array_12_56_real <= _zz_178;
      end
      if(_zz_15)begin
        img_reg_array_13_56_real <= _zz_178;
      end
      if(_zz_16)begin
        img_reg_array_14_56_real <= _zz_178;
      end
      if(_zz_17)begin
        img_reg_array_15_56_real <= _zz_178;
      end
      if(_zz_18)begin
        img_reg_array_16_56_real <= _zz_178;
      end
      if(_zz_19)begin
        img_reg_array_17_56_real <= _zz_178;
      end
      if(_zz_20)begin
        img_reg_array_18_56_real <= _zz_178;
      end
      if(_zz_21)begin
        img_reg_array_19_56_real <= _zz_178;
      end
      if(_zz_22)begin
        img_reg_array_20_56_real <= _zz_178;
      end
      if(_zz_23)begin
        img_reg_array_21_56_real <= _zz_178;
      end
      if(_zz_24)begin
        img_reg_array_22_56_real <= _zz_178;
      end
      if(_zz_25)begin
        img_reg_array_23_56_real <= _zz_178;
      end
      if(_zz_26)begin
        img_reg_array_24_56_real <= _zz_178;
      end
      if(_zz_27)begin
        img_reg_array_25_56_real <= _zz_178;
      end
      if(_zz_28)begin
        img_reg_array_26_56_real <= _zz_178;
      end
      if(_zz_29)begin
        img_reg_array_27_56_real <= _zz_178;
      end
      if(_zz_30)begin
        img_reg_array_28_56_real <= _zz_178;
      end
      if(_zz_31)begin
        img_reg_array_29_56_real <= _zz_178;
      end
      if(_zz_32)begin
        img_reg_array_30_56_real <= _zz_178;
      end
      if(_zz_33)begin
        img_reg_array_31_56_real <= _zz_178;
      end
      if(_zz_34)begin
        img_reg_array_32_56_real <= _zz_178;
      end
      if(_zz_35)begin
        img_reg_array_33_56_real <= _zz_178;
      end
      if(_zz_36)begin
        img_reg_array_34_56_real <= _zz_178;
      end
      if(_zz_37)begin
        img_reg_array_35_56_real <= _zz_178;
      end
      if(_zz_38)begin
        img_reg_array_36_56_real <= _zz_178;
      end
      if(_zz_39)begin
        img_reg_array_37_56_real <= _zz_178;
      end
      if(_zz_40)begin
        img_reg_array_38_56_real <= _zz_178;
      end
      if(_zz_41)begin
        img_reg_array_39_56_real <= _zz_178;
      end
      if(_zz_42)begin
        img_reg_array_40_56_real <= _zz_178;
      end
      if(_zz_43)begin
        img_reg_array_41_56_real <= _zz_178;
      end
      if(_zz_44)begin
        img_reg_array_42_56_real <= _zz_178;
      end
      if(_zz_45)begin
        img_reg_array_43_56_real <= _zz_178;
      end
      if(_zz_46)begin
        img_reg_array_44_56_real <= _zz_178;
      end
      if(_zz_47)begin
        img_reg_array_45_56_real <= _zz_178;
      end
      if(_zz_48)begin
        img_reg_array_46_56_real <= _zz_178;
      end
      if(_zz_49)begin
        img_reg_array_47_56_real <= _zz_178;
      end
      if(_zz_50)begin
        img_reg_array_48_56_real <= _zz_178;
      end
      if(_zz_51)begin
        img_reg_array_49_56_real <= _zz_178;
      end
      if(_zz_52)begin
        img_reg_array_50_56_real <= _zz_178;
      end
      if(_zz_53)begin
        img_reg_array_51_56_real <= _zz_178;
      end
      if(_zz_54)begin
        img_reg_array_52_56_real <= _zz_178;
      end
      if(_zz_55)begin
        img_reg_array_53_56_real <= _zz_178;
      end
      if(_zz_56)begin
        img_reg_array_54_56_real <= _zz_178;
      end
      if(_zz_57)begin
        img_reg_array_55_56_real <= _zz_178;
      end
      if(_zz_58)begin
        img_reg_array_56_56_real <= _zz_178;
      end
      if(_zz_59)begin
        img_reg_array_57_56_real <= _zz_178;
      end
      if(_zz_60)begin
        img_reg_array_58_56_real <= _zz_178;
      end
      if(_zz_61)begin
        img_reg_array_59_56_real <= _zz_178;
      end
      if(_zz_62)begin
        img_reg_array_60_56_real <= _zz_178;
      end
      if(_zz_63)begin
        img_reg_array_61_56_real <= _zz_178;
      end
      if(_zz_64)begin
        img_reg_array_62_56_real <= _zz_178;
      end
      if(_zz_65)begin
        img_reg_array_63_56_real <= _zz_178;
      end
      if(_zz_2)begin
        img_reg_array_0_56_imag <= _zz_179;
      end
      if(_zz_3)begin
        img_reg_array_1_56_imag <= _zz_179;
      end
      if(_zz_4)begin
        img_reg_array_2_56_imag <= _zz_179;
      end
      if(_zz_5)begin
        img_reg_array_3_56_imag <= _zz_179;
      end
      if(_zz_6)begin
        img_reg_array_4_56_imag <= _zz_179;
      end
      if(_zz_7)begin
        img_reg_array_5_56_imag <= _zz_179;
      end
      if(_zz_8)begin
        img_reg_array_6_56_imag <= _zz_179;
      end
      if(_zz_9)begin
        img_reg_array_7_56_imag <= _zz_179;
      end
      if(_zz_10)begin
        img_reg_array_8_56_imag <= _zz_179;
      end
      if(_zz_11)begin
        img_reg_array_9_56_imag <= _zz_179;
      end
      if(_zz_12)begin
        img_reg_array_10_56_imag <= _zz_179;
      end
      if(_zz_13)begin
        img_reg_array_11_56_imag <= _zz_179;
      end
      if(_zz_14)begin
        img_reg_array_12_56_imag <= _zz_179;
      end
      if(_zz_15)begin
        img_reg_array_13_56_imag <= _zz_179;
      end
      if(_zz_16)begin
        img_reg_array_14_56_imag <= _zz_179;
      end
      if(_zz_17)begin
        img_reg_array_15_56_imag <= _zz_179;
      end
      if(_zz_18)begin
        img_reg_array_16_56_imag <= _zz_179;
      end
      if(_zz_19)begin
        img_reg_array_17_56_imag <= _zz_179;
      end
      if(_zz_20)begin
        img_reg_array_18_56_imag <= _zz_179;
      end
      if(_zz_21)begin
        img_reg_array_19_56_imag <= _zz_179;
      end
      if(_zz_22)begin
        img_reg_array_20_56_imag <= _zz_179;
      end
      if(_zz_23)begin
        img_reg_array_21_56_imag <= _zz_179;
      end
      if(_zz_24)begin
        img_reg_array_22_56_imag <= _zz_179;
      end
      if(_zz_25)begin
        img_reg_array_23_56_imag <= _zz_179;
      end
      if(_zz_26)begin
        img_reg_array_24_56_imag <= _zz_179;
      end
      if(_zz_27)begin
        img_reg_array_25_56_imag <= _zz_179;
      end
      if(_zz_28)begin
        img_reg_array_26_56_imag <= _zz_179;
      end
      if(_zz_29)begin
        img_reg_array_27_56_imag <= _zz_179;
      end
      if(_zz_30)begin
        img_reg_array_28_56_imag <= _zz_179;
      end
      if(_zz_31)begin
        img_reg_array_29_56_imag <= _zz_179;
      end
      if(_zz_32)begin
        img_reg_array_30_56_imag <= _zz_179;
      end
      if(_zz_33)begin
        img_reg_array_31_56_imag <= _zz_179;
      end
      if(_zz_34)begin
        img_reg_array_32_56_imag <= _zz_179;
      end
      if(_zz_35)begin
        img_reg_array_33_56_imag <= _zz_179;
      end
      if(_zz_36)begin
        img_reg_array_34_56_imag <= _zz_179;
      end
      if(_zz_37)begin
        img_reg_array_35_56_imag <= _zz_179;
      end
      if(_zz_38)begin
        img_reg_array_36_56_imag <= _zz_179;
      end
      if(_zz_39)begin
        img_reg_array_37_56_imag <= _zz_179;
      end
      if(_zz_40)begin
        img_reg_array_38_56_imag <= _zz_179;
      end
      if(_zz_41)begin
        img_reg_array_39_56_imag <= _zz_179;
      end
      if(_zz_42)begin
        img_reg_array_40_56_imag <= _zz_179;
      end
      if(_zz_43)begin
        img_reg_array_41_56_imag <= _zz_179;
      end
      if(_zz_44)begin
        img_reg_array_42_56_imag <= _zz_179;
      end
      if(_zz_45)begin
        img_reg_array_43_56_imag <= _zz_179;
      end
      if(_zz_46)begin
        img_reg_array_44_56_imag <= _zz_179;
      end
      if(_zz_47)begin
        img_reg_array_45_56_imag <= _zz_179;
      end
      if(_zz_48)begin
        img_reg_array_46_56_imag <= _zz_179;
      end
      if(_zz_49)begin
        img_reg_array_47_56_imag <= _zz_179;
      end
      if(_zz_50)begin
        img_reg_array_48_56_imag <= _zz_179;
      end
      if(_zz_51)begin
        img_reg_array_49_56_imag <= _zz_179;
      end
      if(_zz_52)begin
        img_reg_array_50_56_imag <= _zz_179;
      end
      if(_zz_53)begin
        img_reg_array_51_56_imag <= _zz_179;
      end
      if(_zz_54)begin
        img_reg_array_52_56_imag <= _zz_179;
      end
      if(_zz_55)begin
        img_reg_array_53_56_imag <= _zz_179;
      end
      if(_zz_56)begin
        img_reg_array_54_56_imag <= _zz_179;
      end
      if(_zz_57)begin
        img_reg_array_55_56_imag <= _zz_179;
      end
      if(_zz_58)begin
        img_reg_array_56_56_imag <= _zz_179;
      end
      if(_zz_59)begin
        img_reg_array_57_56_imag <= _zz_179;
      end
      if(_zz_60)begin
        img_reg_array_58_56_imag <= _zz_179;
      end
      if(_zz_61)begin
        img_reg_array_59_56_imag <= _zz_179;
      end
      if(_zz_62)begin
        img_reg_array_60_56_imag <= _zz_179;
      end
      if(_zz_63)begin
        img_reg_array_61_56_imag <= _zz_179;
      end
      if(_zz_64)begin
        img_reg_array_62_56_imag <= _zz_179;
      end
      if(_zz_65)begin
        img_reg_array_63_56_imag <= _zz_179;
      end
      if(_zz_2)begin
        img_reg_array_0_57_real <= _zz_180;
      end
      if(_zz_3)begin
        img_reg_array_1_57_real <= _zz_180;
      end
      if(_zz_4)begin
        img_reg_array_2_57_real <= _zz_180;
      end
      if(_zz_5)begin
        img_reg_array_3_57_real <= _zz_180;
      end
      if(_zz_6)begin
        img_reg_array_4_57_real <= _zz_180;
      end
      if(_zz_7)begin
        img_reg_array_5_57_real <= _zz_180;
      end
      if(_zz_8)begin
        img_reg_array_6_57_real <= _zz_180;
      end
      if(_zz_9)begin
        img_reg_array_7_57_real <= _zz_180;
      end
      if(_zz_10)begin
        img_reg_array_8_57_real <= _zz_180;
      end
      if(_zz_11)begin
        img_reg_array_9_57_real <= _zz_180;
      end
      if(_zz_12)begin
        img_reg_array_10_57_real <= _zz_180;
      end
      if(_zz_13)begin
        img_reg_array_11_57_real <= _zz_180;
      end
      if(_zz_14)begin
        img_reg_array_12_57_real <= _zz_180;
      end
      if(_zz_15)begin
        img_reg_array_13_57_real <= _zz_180;
      end
      if(_zz_16)begin
        img_reg_array_14_57_real <= _zz_180;
      end
      if(_zz_17)begin
        img_reg_array_15_57_real <= _zz_180;
      end
      if(_zz_18)begin
        img_reg_array_16_57_real <= _zz_180;
      end
      if(_zz_19)begin
        img_reg_array_17_57_real <= _zz_180;
      end
      if(_zz_20)begin
        img_reg_array_18_57_real <= _zz_180;
      end
      if(_zz_21)begin
        img_reg_array_19_57_real <= _zz_180;
      end
      if(_zz_22)begin
        img_reg_array_20_57_real <= _zz_180;
      end
      if(_zz_23)begin
        img_reg_array_21_57_real <= _zz_180;
      end
      if(_zz_24)begin
        img_reg_array_22_57_real <= _zz_180;
      end
      if(_zz_25)begin
        img_reg_array_23_57_real <= _zz_180;
      end
      if(_zz_26)begin
        img_reg_array_24_57_real <= _zz_180;
      end
      if(_zz_27)begin
        img_reg_array_25_57_real <= _zz_180;
      end
      if(_zz_28)begin
        img_reg_array_26_57_real <= _zz_180;
      end
      if(_zz_29)begin
        img_reg_array_27_57_real <= _zz_180;
      end
      if(_zz_30)begin
        img_reg_array_28_57_real <= _zz_180;
      end
      if(_zz_31)begin
        img_reg_array_29_57_real <= _zz_180;
      end
      if(_zz_32)begin
        img_reg_array_30_57_real <= _zz_180;
      end
      if(_zz_33)begin
        img_reg_array_31_57_real <= _zz_180;
      end
      if(_zz_34)begin
        img_reg_array_32_57_real <= _zz_180;
      end
      if(_zz_35)begin
        img_reg_array_33_57_real <= _zz_180;
      end
      if(_zz_36)begin
        img_reg_array_34_57_real <= _zz_180;
      end
      if(_zz_37)begin
        img_reg_array_35_57_real <= _zz_180;
      end
      if(_zz_38)begin
        img_reg_array_36_57_real <= _zz_180;
      end
      if(_zz_39)begin
        img_reg_array_37_57_real <= _zz_180;
      end
      if(_zz_40)begin
        img_reg_array_38_57_real <= _zz_180;
      end
      if(_zz_41)begin
        img_reg_array_39_57_real <= _zz_180;
      end
      if(_zz_42)begin
        img_reg_array_40_57_real <= _zz_180;
      end
      if(_zz_43)begin
        img_reg_array_41_57_real <= _zz_180;
      end
      if(_zz_44)begin
        img_reg_array_42_57_real <= _zz_180;
      end
      if(_zz_45)begin
        img_reg_array_43_57_real <= _zz_180;
      end
      if(_zz_46)begin
        img_reg_array_44_57_real <= _zz_180;
      end
      if(_zz_47)begin
        img_reg_array_45_57_real <= _zz_180;
      end
      if(_zz_48)begin
        img_reg_array_46_57_real <= _zz_180;
      end
      if(_zz_49)begin
        img_reg_array_47_57_real <= _zz_180;
      end
      if(_zz_50)begin
        img_reg_array_48_57_real <= _zz_180;
      end
      if(_zz_51)begin
        img_reg_array_49_57_real <= _zz_180;
      end
      if(_zz_52)begin
        img_reg_array_50_57_real <= _zz_180;
      end
      if(_zz_53)begin
        img_reg_array_51_57_real <= _zz_180;
      end
      if(_zz_54)begin
        img_reg_array_52_57_real <= _zz_180;
      end
      if(_zz_55)begin
        img_reg_array_53_57_real <= _zz_180;
      end
      if(_zz_56)begin
        img_reg_array_54_57_real <= _zz_180;
      end
      if(_zz_57)begin
        img_reg_array_55_57_real <= _zz_180;
      end
      if(_zz_58)begin
        img_reg_array_56_57_real <= _zz_180;
      end
      if(_zz_59)begin
        img_reg_array_57_57_real <= _zz_180;
      end
      if(_zz_60)begin
        img_reg_array_58_57_real <= _zz_180;
      end
      if(_zz_61)begin
        img_reg_array_59_57_real <= _zz_180;
      end
      if(_zz_62)begin
        img_reg_array_60_57_real <= _zz_180;
      end
      if(_zz_63)begin
        img_reg_array_61_57_real <= _zz_180;
      end
      if(_zz_64)begin
        img_reg_array_62_57_real <= _zz_180;
      end
      if(_zz_65)begin
        img_reg_array_63_57_real <= _zz_180;
      end
      if(_zz_2)begin
        img_reg_array_0_57_imag <= _zz_181;
      end
      if(_zz_3)begin
        img_reg_array_1_57_imag <= _zz_181;
      end
      if(_zz_4)begin
        img_reg_array_2_57_imag <= _zz_181;
      end
      if(_zz_5)begin
        img_reg_array_3_57_imag <= _zz_181;
      end
      if(_zz_6)begin
        img_reg_array_4_57_imag <= _zz_181;
      end
      if(_zz_7)begin
        img_reg_array_5_57_imag <= _zz_181;
      end
      if(_zz_8)begin
        img_reg_array_6_57_imag <= _zz_181;
      end
      if(_zz_9)begin
        img_reg_array_7_57_imag <= _zz_181;
      end
      if(_zz_10)begin
        img_reg_array_8_57_imag <= _zz_181;
      end
      if(_zz_11)begin
        img_reg_array_9_57_imag <= _zz_181;
      end
      if(_zz_12)begin
        img_reg_array_10_57_imag <= _zz_181;
      end
      if(_zz_13)begin
        img_reg_array_11_57_imag <= _zz_181;
      end
      if(_zz_14)begin
        img_reg_array_12_57_imag <= _zz_181;
      end
      if(_zz_15)begin
        img_reg_array_13_57_imag <= _zz_181;
      end
      if(_zz_16)begin
        img_reg_array_14_57_imag <= _zz_181;
      end
      if(_zz_17)begin
        img_reg_array_15_57_imag <= _zz_181;
      end
      if(_zz_18)begin
        img_reg_array_16_57_imag <= _zz_181;
      end
      if(_zz_19)begin
        img_reg_array_17_57_imag <= _zz_181;
      end
      if(_zz_20)begin
        img_reg_array_18_57_imag <= _zz_181;
      end
      if(_zz_21)begin
        img_reg_array_19_57_imag <= _zz_181;
      end
      if(_zz_22)begin
        img_reg_array_20_57_imag <= _zz_181;
      end
      if(_zz_23)begin
        img_reg_array_21_57_imag <= _zz_181;
      end
      if(_zz_24)begin
        img_reg_array_22_57_imag <= _zz_181;
      end
      if(_zz_25)begin
        img_reg_array_23_57_imag <= _zz_181;
      end
      if(_zz_26)begin
        img_reg_array_24_57_imag <= _zz_181;
      end
      if(_zz_27)begin
        img_reg_array_25_57_imag <= _zz_181;
      end
      if(_zz_28)begin
        img_reg_array_26_57_imag <= _zz_181;
      end
      if(_zz_29)begin
        img_reg_array_27_57_imag <= _zz_181;
      end
      if(_zz_30)begin
        img_reg_array_28_57_imag <= _zz_181;
      end
      if(_zz_31)begin
        img_reg_array_29_57_imag <= _zz_181;
      end
      if(_zz_32)begin
        img_reg_array_30_57_imag <= _zz_181;
      end
      if(_zz_33)begin
        img_reg_array_31_57_imag <= _zz_181;
      end
      if(_zz_34)begin
        img_reg_array_32_57_imag <= _zz_181;
      end
      if(_zz_35)begin
        img_reg_array_33_57_imag <= _zz_181;
      end
      if(_zz_36)begin
        img_reg_array_34_57_imag <= _zz_181;
      end
      if(_zz_37)begin
        img_reg_array_35_57_imag <= _zz_181;
      end
      if(_zz_38)begin
        img_reg_array_36_57_imag <= _zz_181;
      end
      if(_zz_39)begin
        img_reg_array_37_57_imag <= _zz_181;
      end
      if(_zz_40)begin
        img_reg_array_38_57_imag <= _zz_181;
      end
      if(_zz_41)begin
        img_reg_array_39_57_imag <= _zz_181;
      end
      if(_zz_42)begin
        img_reg_array_40_57_imag <= _zz_181;
      end
      if(_zz_43)begin
        img_reg_array_41_57_imag <= _zz_181;
      end
      if(_zz_44)begin
        img_reg_array_42_57_imag <= _zz_181;
      end
      if(_zz_45)begin
        img_reg_array_43_57_imag <= _zz_181;
      end
      if(_zz_46)begin
        img_reg_array_44_57_imag <= _zz_181;
      end
      if(_zz_47)begin
        img_reg_array_45_57_imag <= _zz_181;
      end
      if(_zz_48)begin
        img_reg_array_46_57_imag <= _zz_181;
      end
      if(_zz_49)begin
        img_reg_array_47_57_imag <= _zz_181;
      end
      if(_zz_50)begin
        img_reg_array_48_57_imag <= _zz_181;
      end
      if(_zz_51)begin
        img_reg_array_49_57_imag <= _zz_181;
      end
      if(_zz_52)begin
        img_reg_array_50_57_imag <= _zz_181;
      end
      if(_zz_53)begin
        img_reg_array_51_57_imag <= _zz_181;
      end
      if(_zz_54)begin
        img_reg_array_52_57_imag <= _zz_181;
      end
      if(_zz_55)begin
        img_reg_array_53_57_imag <= _zz_181;
      end
      if(_zz_56)begin
        img_reg_array_54_57_imag <= _zz_181;
      end
      if(_zz_57)begin
        img_reg_array_55_57_imag <= _zz_181;
      end
      if(_zz_58)begin
        img_reg_array_56_57_imag <= _zz_181;
      end
      if(_zz_59)begin
        img_reg_array_57_57_imag <= _zz_181;
      end
      if(_zz_60)begin
        img_reg_array_58_57_imag <= _zz_181;
      end
      if(_zz_61)begin
        img_reg_array_59_57_imag <= _zz_181;
      end
      if(_zz_62)begin
        img_reg_array_60_57_imag <= _zz_181;
      end
      if(_zz_63)begin
        img_reg_array_61_57_imag <= _zz_181;
      end
      if(_zz_64)begin
        img_reg_array_62_57_imag <= _zz_181;
      end
      if(_zz_65)begin
        img_reg_array_63_57_imag <= _zz_181;
      end
      if(_zz_2)begin
        img_reg_array_0_58_real <= _zz_182;
      end
      if(_zz_3)begin
        img_reg_array_1_58_real <= _zz_182;
      end
      if(_zz_4)begin
        img_reg_array_2_58_real <= _zz_182;
      end
      if(_zz_5)begin
        img_reg_array_3_58_real <= _zz_182;
      end
      if(_zz_6)begin
        img_reg_array_4_58_real <= _zz_182;
      end
      if(_zz_7)begin
        img_reg_array_5_58_real <= _zz_182;
      end
      if(_zz_8)begin
        img_reg_array_6_58_real <= _zz_182;
      end
      if(_zz_9)begin
        img_reg_array_7_58_real <= _zz_182;
      end
      if(_zz_10)begin
        img_reg_array_8_58_real <= _zz_182;
      end
      if(_zz_11)begin
        img_reg_array_9_58_real <= _zz_182;
      end
      if(_zz_12)begin
        img_reg_array_10_58_real <= _zz_182;
      end
      if(_zz_13)begin
        img_reg_array_11_58_real <= _zz_182;
      end
      if(_zz_14)begin
        img_reg_array_12_58_real <= _zz_182;
      end
      if(_zz_15)begin
        img_reg_array_13_58_real <= _zz_182;
      end
      if(_zz_16)begin
        img_reg_array_14_58_real <= _zz_182;
      end
      if(_zz_17)begin
        img_reg_array_15_58_real <= _zz_182;
      end
      if(_zz_18)begin
        img_reg_array_16_58_real <= _zz_182;
      end
      if(_zz_19)begin
        img_reg_array_17_58_real <= _zz_182;
      end
      if(_zz_20)begin
        img_reg_array_18_58_real <= _zz_182;
      end
      if(_zz_21)begin
        img_reg_array_19_58_real <= _zz_182;
      end
      if(_zz_22)begin
        img_reg_array_20_58_real <= _zz_182;
      end
      if(_zz_23)begin
        img_reg_array_21_58_real <= _zz_182;
      end
      if(_zz_24)begin
        img_reg_array_22_58_real <= _zz_182;
      end
      if(_zz_25)begin
        img_reg_array_23_58_real <= _zz_182;
      end
      if(_zz_26)begin
        img_reg_array_24_58_real <= _zz_182;
      end
      if(_zz_27)begin
        img_reg_array_25_58_real <= _zz_182;
      end
      if(_zz_28)begin
        img_reg_array_26_58_real <= _zz_182;
      end
      if(_zz_29)begin
        img_reg_array_27_58_real <= _zz_182;
      end
      if(_zz_30)begin
        img_reg_array_28_58_real <= _zz_182;
      end
      if(_zz_31)begin
        img_reg_array_29_58_real <= _zz_182;
      end
      if(_zz_32)begin
        img_reg_array_30_58_real <= _zz_182;
      end
      if(_zz_33)begin
        img_reg_array_31_58_real <= _zz_182;
      end
      if(_zz_34)begin
        img_reg_array_32_58_real <= _zz_182;
      end
      if(_zz_35)begin
        img_reg_array_33_58_real <= _zz_182;
      end
      if(_zz_36)begin
        img_reg_array_34_58_real <= _zz_182;
      end
      if(_zz_37)begin
        img_reg_array_35_58_real <= _zz_182;
      end
      if(_zz_38)begin
        img_reg_array_36_58_real <= _zz_182;
      end
      if(_zz_39)begin
        img_reg_array_37_58_real <= _zz_182;
      end
      if(_zz_40)begin
        img_reg_array_38_58_real <= _zz_182;
      end
      if(_zz_41)begin
        img_reg_array_39_58_real <= _zz_182;
      end
      if(_zz_42)begin
        img_reg_array_40_58_real <= _zz_182;
      end
      if(_zz_43)begin
        img_reg_array_41_58_real <= _zz_182;
      end
      if(_zz_44)begin
        img_reg_array_42_58_real <= _zz_182;
      end
      if(_zz_45)begin
        img_reg_array_43_58_real <= _zz_182;
      end
      if(_zz_46)begin
        img_reg_array_44_58_real <= _zz_182;
      end
      if(_zz_47)begin
        img_reg_array_45_58_real <= _zz_182;
      end
      if(_zz_48)begin
        img_reg_array_46_58_real <= _zz_182;
      end
      if(_zz_49)begin
        img_reg_array_47_58_real <= _zz_182;
      end
      if(_zz_50)begin
        img_reg_array_48_58_real <= _zz_182;
      end
      if(_zz_51)begin
        img_reg_array_49_58_real <= _zz_182;
      end
      if(_zz_52)begin
        img_reg_array_50_58_real <= _zz_182;
      end
      if(_zz_53)begin
        img_reg_array_51_58_real <= _zz_182;
      end
      if(_zz_54)begin
        img_reg_array_52_58_real <= _zz_182;
      end
      if(_zz_55)begin
        img_reg_array_53_58_real <= _zz_182;
      end
      if(_zz_56)begin
        img_reg_array_54_58_real <= _zz_182;
      end
      if(_zz_57)begin
        img_reg_array_55_58_real <= _zz_182;
      end
      if(_zz_58)begin
        img_reg_array_56_58_real <= _zz_182;
      end
      if(_zz_59)begin
        img_reg_array_57_58_real <= _zz_182;
      end
      if(_zz_60)begin
        img_reg_array_58_58_real <= _zz_182;
      end
      if(_zz_61)begin
        img_reg_array_59_58_real <= _zz_182;
      end
      if(_zz_62)begin
        img_reg_array_60_58_real <= _zz_182;
      end
      if(_zz_63)begin
        img_reg_array_61_58_real <= _zz_182;
      end
      if(_zz_64)begin
        img_reg_array_62_58_real <= _zz_182;
      end
      if(_zz_65)begin
        img_reg_array_63_58_real <= _zz_182;
      end
      if(_zz_2)begin
        img_reg_array_0_58_imag <= _zz_183;
      end
      if(_zz_3)begin
        img_reg_array_1_58_imag <= _zz_183;
      end
      if(_zz_4)begin
        img_reg_array_2_58_imag <= _zz_183;
      end
      if(_zz_5)begin
        img_reg_array_3_58_imag <= _zz_183;
      end
      if(_zz_6)begin
        img_reg_array_4_58_imag <= _zz_183;
      end
      if(_zz_7)begin
        img_reg_array_5_58_imag <= _zz_183;
      end
      if(_zz_8)begin
        img_reg_array_6_58_imag <= _zz_183;
      end
      if(_zz_9)begin
        img_reg_array_7_58_imag <= _zz_183;
      end
      if(_zz_10)begin
        img_reg_array_8_58_imag <= _zz_183;
      end
      if(_zz_11)begin
        img_reg_array_9_58_imag <= _zz_183;
      end
      if(_zz_12)begin
        img_reg_array_10_58_imag <= _zz_183;
      end
      if(_zz_13)begin
        img_reg_array_11_58_imag <= _zz_183;
      end
      if(_zz_14)begin
        img_reg_array_12_58_imag <= _zz_183;
      end
      if(_zz_15)begin
        img_reg_array_13_58_imag <= _zz_183;
      end
      if(_zz_16)begin
        img_reg_array_14_58_imag <= _zz_183;
      end
      if(_zz_17)begin
        img_reg_array_15_58_imag <= _zz_183;
      end
      if(_zz_18)begin
        img_reg_array_16_58_imag <= _zz_183;
      end
      if(_zz_19)begin
        img_reg_array_17_58_imag <= _zz_183;
      end
      if(_zz_20)begin
        img_reg_array_18_58_imag <= _zz_183;
      end
      if(_zz_21)begin
        img_reg_array_19_58_imag <= _zz_183;
      end
      if(_zz_22)begin
        img_reg_array_20_58_imag <= _zz_183;
      end
      if(_zz_23)begin
        img_reg_array_21_58_imag <= _zz_183;
      end
      if(_zz_24)begin
        img_reg_array_22_58_imag <= _zz_183;
      end
      if(_zz_25)begin
        img_reg_array_23_58_imag <= _zz_183;
      end
      if(_zz_26)begin
        img_reg_array_24_58_imag <= _zz_183;
      end
      if(_zz_27)begin
        img_reg_array_25_58_imag <= _zz_183;
      end
      if(_zz_28)begin
        img_reg_array_26_58_imag <= _zz_183;
      end
      if(_zz_29)begin
        img_reg_array_27_58_imag <= _zz_183;
      end
      if(_zz_30)begin
        img_reg_array_28_58_imag <= _zz_183;
      end
      if(_zz_31)begin
        img_reg_array_29_58_imag <= _zz_183;
      end
      if(_zz_32)begin
        img_reg_array_30_58_imag <= _zz_183;
      end
      if(_zz_33)begin
        img_reg_array_31_58_imag <= _zz_183;
      end
      if(_zz_34)begin
        img_reg_array_32_58_imag <= _zz_183;
      end
      if(_zz_35)begin
        img_reg_array_33_58_imag <= _zz_183;
      end
      if(_zz_36)begin
        img_reg_array_34_58_imag <= _zz_183;
      end
      if(_zz_37)begin
        img_reg_array_35_58_imag <= _zz_183;
      end
      if(_zz_38)begin
        img_reg_array_36_58_imag <= _zz_183;
      end
      if(_zz_39)begin
        img_reg_array_37_58_imag <= _zz_183;
      end
      if(_zz_40)begin
        img_reg_array_38_58_imag <= _zz_183;
      end
      if(_zz_41)begin
        img_reg_array_39_58_imag <= _zz_183;
      end
      if(_zz_42)begin
        img_reg_array_40_58_imag <= _zz_183;
      end
      if(_zz_43)begin
        img_reg_array_41_58_imag <= _zz_183;
      end
      if(_zz_44)begin
        img_reg_array_42_58_imag <= _zz_183;
      end
      if(_zz_45)begin
        img_reg_array_43_58_imag <= _zz_183;
      end
      if(_zz_46)begin
        img_reg_array_44_58_imag <= _zz_183;
      end
      if(_zz_47)begin
        img_reg_array_45_58_imag <= _zz_183;
      end
      if(_zz_48)begin
        img_reg_array_46_58_imag <= _zz_183;
      end
      if(_zz_49)begin
        img_reg_array_47_58_imag <= _zz_183;
      end
      if(_zz_50)begin
        img_reg_array_48_58_imag <= _zz_183;
      end
      if(_zz_51)begin
        img_reg_array_49_58_imag <= _zz_183;
      end
      if(_zz_52)begin
        img_reg_array_50_58_imag <= _zz_183;
      end
      if(_zz_53)begin
        img_reg_array_51_58_imag <= _zz_183;
      end
      if(_zz_54)begin
        img_reg_array_52_58_imag <= _zz_183;
      end
      if(_zz_55)begin
        img_reg_array_53_58_imag <= _zz_183;
      end
      if(_zz_56)begin
        img_reg_array_54_58_imag <= _zz_183;
      end
      if(_zz_57)begin
        img_reg_array_55_58_imag <= _zz_183;
      end
      if(_zz_58)begin
        img_reg_array_56_58_imag <= _zz_183;
      end
      if(_zz_59)begin
        img_reg_array_57_58_imag <= _zz_183;
      end
      if(_zz_60)begin
        img_reg_array_58_58_imag <= _zz_183;
      end
      if(_zz_61)begin
        img_reg_array_59_58_imag <= _zz_183;
      end
      if(_zz_62)begin
        img_reg_array_60_58_imag <= _zz_183;
      end
      if(_zz_63)begin
        img_reg_array_61_58_imag <= _zz_183;
      end
      if(_zz_64)begin
        img_reg_array_62_58_imag <= _zz_183;
      end
      if(_zz_65)begin
        img_reg_array_63_58_imag <= _zz_183;
      end
      if(_zz_2)begin
        img_reg_array_0_59_real <= _zz_184;
      end
      if(_zz_3)begin
        img_reg_array_1_59_real <= _zz_184;
      end
      if(_zz_4)begin
        img_reg_array_2_59_real <= _zz_184;
      end
      if(_zz_5)begin
        img_reg_array_3_59_real <= _zz_184;
      end
      if(_zz_6)begin
        img_reg_array_4_59_real <= _zz_184;
      end
      if(_zz_7)begin
        img_reg_array_5_59_real <= _zz_184;
      end
      if(_zz_8)begin
        img_reg_array_6_59_real <= _zz_184;
      end
      if(_zz_9)begin
        img_reg_array_7_59_real <= _zz_184;
      end
      if(_zz_10)begin
        img_reg_array_8_59_real <= _zz_184;
      end
      if(_zz_11)begin
        img_reg_array_9_59_real <= _zz_184;
      end
      if(_zz_12)begin
        img_reg_array_10_59_real <= _zz_184;
      end
      if(_zz_13)begin
        img_reg_array_11_59_real <= _zz_184;
      end
      if(_zz_14)begin
        img_reg_array_12_59_real <= _zz_184;
      end
      if(_zz_15)begin
        img_reg_array_13_59_real <= _zz_184;
      end
      if(_zz_16)begin
        img_reg_array_14_59_real <= _zz_184;
      end
      if(_zz_17)begin
        img_reg_array_15_59_real <= _zz_184;
      end
      if(_zz_18)begin
        img_reg_array_16_59_real <= _zz_184;
      end
      if(_zz_19)begin
        img_reg_array_17_59_real <= _zz_184;
      end
      if(_zz_20)begin
        img_reg_array_18_59_real <= _zz_184;
      end
      if(_zz_21)begin
        img_reg_array_19_59_real <= _zz_184;
      end
      if(_zz_22)begin
        img_reg_array_20_59_real <= _zz_184;
      end
      if(_zz_23)begin
        img_reg_array_21_59_real <= _zz_184;
      end
      if(_zz_24)begin
        img_reg_array_22_59_real <= _zz_184;
      end
      if(_zz_25)begin
        img_reg_array_23_59_real <= _zz_184;
      end
      if(_zz_26)begin
        img_reg_array_24_59_real <= _zz_184;
      end
      if(_zz_27)begin
        img_reg_array_25_59_real <= _zz_184;
      end
      if(_zz_28)begin
        img_reg_array_26_59_real <= _zz_184;
      end
      if(_zz_29)begin
        img_reg_array_27_59_real <= _zz_184;
      end
      if(_zz_30)begin
        img_reg_array_28_59_real <= _zz_184;
      end
      if(_zz_31)begin
        img_reg_array_29_59_real <= _zz_184;
      end
      if(_zz_32)begin
        img_reg_array_30_59_real <= _zz_184;
      end
      if(_zz_33)begin
        img_reg_array_31_59_real <= _zz_184;
      end
      if(_zz_34)begin
        img_reg_array_32_59_real <= _zz_184;
      end
      if(_zz_35)begin
        img_reg_array_33_59_real <= _zz_184;
      end
      if(_zz_36)begin
        img_reg_array_34_59_real <= _zz_184;
      end
      if(_zz_37)begin
        img_reg_array_35_59_real <= _zz_184;
      end
      if(_zz_38)begin
        img_reg_array_36_59_real <= _zz_184;
      end
      if(_zz_39)begin
        img_reg_array_37_59_real <= _zz_184;
      end
      if(_zz_40)begin
        img_reg_array_38_59_real <= _zz_184;
      end
      if(_zz_41)begin
        img_reg_array_39_59_real <= _zz_184;
      end
      if(_zz_42)begin
        img_reg_array_40_59_real <= _zz_184;
      end
      if(_zz_43)begin
        img_reg_array_41_59_real <= _zz_184;
      end
      if(_zz_44)begin
        img_reg_array_42_59_real <= _zz_184;
      end
      if(_zz_45)begin
        img_reg_array_43_59_real <= _zz_184;
      end
      if(_zz_46)begin
        img_reg_array_44_59_real <= _zz_184;
      end
      if(_zz_47)begin
        img_reg_array_45_59_real <= _zz_184;
      end
      if(_zz_48)begin
        img_reg_array_46_59_real <= _zz_184;
      end
      if(_zz_49)begin
        img_reg_array_47_59_real <= _zz_184;
      end
      if(_zz_50)begin
        img_reg_array_48_59_real <= _zz_184;
      end
      if(_zz_51)begin
        img_reg_array_49_59_real <= _zz_184;
      end
      if(_zz_52)begin
        img_reg_array_50_59_real <= _zz_184;
      end
      if(_zz_53)begin
        img_reg_array_51_59_real <= _zz_184;
      end
      if(_zz_54)begin
        img_reg_array_52_59_real <= _zz_184;
      end
      if(_zz_55)begin
        img_reg_array_53_59_real <= _zz_184;
      end
      if(_zz_56)begin
        img_reg_array_54_59_real <= _zz_184;
      end
      if(_zz_57)begin
        img_reg_array_55_59_real <= _zz_184;
      end
      if(_zz_58)begin
        img_reg_array_56_59_real <= _zz_184;
      end
      if(_zz_59)begin
        img_reg_array_57_59_real <= _zz_184;
      end
      if(_zz_60)begin
        img_reg_array_58_59_real <= _zz_184;
      end
      if(_zz_61)begin
        img_reg_array_59_59_real <= _zz_184;
      end
      if(_zz_62)begin
        img_reg_array_60_59_real <= _zz_184;
      end
      if(_zz_63)begin
        img_reg_array_61_59_real <= _zz_184;
      end
      if(_zz_64)begin
        img_reg_array_62_59_real <= _zz_184;
      end
      if(_zz_65)begin
        img_reg_array_63_59_real <= _zz_184;
      end
      if(_zz_2)begin
        img_reg_array_0_59_imag <= _zz_185;
      end
      if(_zz_3)begin
        img_reg_array_1_59_imag <= _zz_185;
      end
      if(_zz_4)begin
        img_reg_array_2_59_imag <= _zz_185;
      end
      if(_zz_5)begin
        img_reg_array_3_59_imag <= _zz_185;
      end
      if(_zz_6)begin
        img_reg_array_4_59_imag <= _zz_185;
      end
      if(_zz_7)begin
        img_reg_array_5_59_imag <= _zz_185;
      end
      if(_zz_8)begin
        img_reg_array_6_59_imag <= _zz_185;
      end
      if(_zz_9)begin
        img_reg_array_7_59_imag <= _zz_185;
      end
      if(_zz_10)begin
        img_reg_array_8_59_imag <= _zz_185;
      end
      if(_zz_11)begin
        img_reg_array_9_59_imag <= _zz_185;
      end
      if(_zz_12)begin
        img_reg_array_10_59_imag <= _zz_185;
      end
      if(_zz_13)begin
        img_reg_array_11_59_imag <= _zz_185;
      end
      if(_zz_14)begin
        img_reg_array_12_59_imag <= _zz_185;
      end
      if(_zz_15)begin
        img_reg_array_13_59_imag <= _zz_185;
      end
      if(_zz_16)begin
        img_reg_array_14_59_imag <= _zz_185;
      end
      if(_zz_17)begin
        img_reg_array_15_59_imag <= _zz_185;
      end
      if(_zz_18)begin
        img_reg_array_16_59_imag <= _zz_185;
      end
      if(_zz_19)begin
        img_reg_array_17_59_imag <= _zz_185;
      end
      if(_zz_20)begin
        img_reg_array_18_59_imag <= _zz_185;
      end
      if(_zz_21)begin
        img_reg_array_19_59_imag <= _zz_185;
      end
      if(_zz_22)begin
        img_reg_array_20_59_imag <= _zz_185;
      end
      if(_zz_23)begin
        img_reg_array_21_59_imag <= _zz_185;
      end
      if(_zz_24)begin
        img_reg_array_22_59_imag <= _zz_185;
      end
      if(_zz_25)begin
        img_reg_array_23_59_imag <= _zz_185;
      end
      if(_zz_26)begin
        img_reg_array_24_59_imag <= _zz_185;
      end
      if(_zz_27)begin
        img_reg_array_25_59_imag <= _zz_185;
      end
      if(_zz_28)begin
        img_reg_array_26_59_imag <= _zz_185;
      end
      if(_zz_29)begin
        img_reg_array_27_59_imag <= _zz_185;
      end
      if(_zz_30)begin
        img_reg_array_28_59_imag <= _zz_185;
      end
      if(_zz_31)begin
        img_reg_array_29_59_imag <= _zz_185;
      end
      if(_zz_32)begin
        img_reg_array_30_59_imag <= _zz_185;
      end
      if(_zz_33)begin
        img_reg_array_31_59_imag <= _zz_185;
      end
      if(_zz_34)begin
        img_reg_array_32_59_imag <= _zz_185;
      end
      if(_zz_35)begin
        img_reg_array_33_59_imag <= _zz_185;
      end
      if(_zz_36)begin
        img_reg_array_34_59_imag <= _zz_185;
      end
      if(_zz_37)begin
        img_reg_array_35_59_imag <= _zz_185;
      end
      if(_zz_38)begin
        img_reg_array_36_59_imag <= _zz_185;
      end
      if(_zz_39)begin
        img_reg_array_37_59_imag <= _zz_185;
      end
      if(_zz_40)begin
        img_reg_array_38_59_imag <= _zz_185;
      end
      if(_zz_41)begin
        img_reg_array_39_59_imag <= _zz_185;
      end
      if(_zz_42)begin
        img_reg_array_40_59_imag <= _zz_185;
      end
      if(_zz_43)begin
        img_reg_array_41_59_imag <= _zz_185;
      end
      if(_zz_44)begin
        img_reg_array_42_59_imag <= _zz_185;
      end
      if(_zz_45)begin
        img_reg_array_43_59_imag <= _zz_185;
      end
      if(_zz_46)begin
        img_reg_array_44_59_imag <= _zz_185;
      end
      if(_zz_47)begin
        img_reg_array_45_59_imag <= _zz_185;
      end
      if(_zz_48)begin
        img_reg_array_46_59_imag <= _zz_185;
      end
      if(_zz_49)begin
        img_reg_array_47_59_imag <= _zz_185;
      end
      if(_zz_50)begin
        img_reg_array_48_59_imag <= _zz_185;
      end
      if(_zz_51)begin
        img_reg_array_49_59_imag <= _zz_185;
      end
      if(_zz_52)begin
        img_reg_array_50_59_imag <= _zz_185;
      end
      if(_zz_53)begin
        img_reg_array_51_59_imag <= _zz_185;
      end
      if(_zz_54)begin
        img_reg_array_52_59_imag <= _zz_185;
      end
      if(_zz_55)begin
        img_reg_array_53_59_imag <= _zz_185;
      end
      if(_zz_56)begin
        img_reg_array_54_59_imag <= _zz_185;
      end
      if(_zz_57)begin
        img_reg_array_55_59_imag <= _zz_185;
      end
      if(_zz_58)begin
        img_reg_array_56_59_imag <= _zz_185;
      end
      if(_zz_59)begin
        img_reg_array_57_59_imag <= _zz_185;
      end
      if(_zz_60)begin
        img_reg_array_58_59_imag <= _zz_185;
      end
      if(_zz_61)begin
        img_reg_array_59_59_imag <= _zz_185;
      end
      if(_zz_62)begin
        img_reg_array_60_59_imag <= _zz_185;
      end
      if(_zz_63)begin
        img_reg_array_61_59_imag <= _zz_185;
      end
      if(_zz_64)begin
        img_reg_array_62_59_imag <= _zz_185;
      end
      if(_zz_65)begin
        img_reg_array_63_59_imag <= _zz_185;
      end
      if(_zz_2)begin
        img_reg_array_0_60_real <= _zz_186;
      end
      if(_zz_3)begin
        img_reg_array_1_60_real <= _zz_186;
      end
      if(_zz_4)begin
        img_reg_array_2_60_real <= _zz_186;
      end
      if(_zz_5)begin
        img_reg_array_3_60_real <= _zz_186;
      end
      if(_zz_6)begin
        img_reg_array_4_60_real <= _zz_186;
      end
      if(_zz_7)begin
        img_reg_array_5_60_real <= _zz_186;
      end
      if(_zz_8)begin
        img_reg_array_6_60_real <= _zz_186;
      end
      if(_zz_9)begin
        img_reg_array_7_60_real <= _zz_186;
      end
      if(_zz_10)begin
        img_reg_array_8_60_real <= _zz_186;
      end
      if(_zz_11)begin
        img_reg_array_9_60_real <= _zz_186;
      end
      if(_zz_12)begin
        img_reg_array_10_60_real <= _zz_186;
      end
      if(_zz_13)begin
        img_reg_array_11_60_real <= _zz_186;
      end
      if(_zz_14)begin
        img_reg_array_12_60_real <= _zz_186;
      end
      if(_zz_15)begin
        img_reg_array_13_60_real <= _zz_186;
      end
      if(_zz_16)begin
        img_reg_array_14_60_real <= _zz_186;
      end
      if(_zz_17)begin
        img_reg_array_15_60_real <= _zz_186;
      end
      if(_zz_18)begin
        img_reg_array_16_60_real <= _zz_186;
      end
      if(_zz_19)begin
        img_reg_array_17_60_real <= _zz_186;
      end
      if(_zz_20)begin
        img_reg_array_18_60_real <= _zz_186;
      end
      if(_zz_21)begin
        img_reg_array_19_60_real <= _zz_186;
      end
      if(_zz_22)begin
        img_reg_array_20_60_real <= _zz_186;
      end
      if(_zz_23)begin
        img_reg_array_21_60_real <= _zz_186;
      end
      if(_zz_24)begin
        img_reg_array_22_60_real <= _zz_186;
      end
      if(_zz_25)begin
        img_reg_array_23_60_real <= _zz_186;
      end
      if(_zz_26)begin
        img_reg_array_24_60_real <= _zz_186;
      end
      if(_zz_27)begin
        img_reg_array_25_60_real <= _zz_186;
      end
      if(_zz_28)begin
        img_reg_array_26_60_real <= _zz_186;
      end
      if(_zz_29)begin
        img_reg_array_27_60_real <= _zz_186;
      end
      if(_zz_30)begin
        img_reg_array_28_60_real <= _zz_186;
      end
      if(_zz_31)begin
        img_reg_array_29_60_real <= _zz_186;
      end
      if(_zz_32)begin
        img_reg_array_30_60_real <= _zz_186;
      end
      if(_zz_33)begin
        img_reg_array_31_60_real <= _zz_186;
      end
      if(_zz_34)begin
        img_reg_array_32_60_real <= _zz_186;
      end
      if(_zz_35)begin
        img_reg_array_33_60_real <= _zz_186;
      end
      if(_zz_36)begin
        img_reg_array_34_60_real <= _zz_186;
      end
      if(_zz_37)begin
        img_reg_array_35_60_real <= _zz_186;
      end
      if(_zz_38)begin
        img_reg_array_36_60_real <= _zz_186;
      end
      if(_zz_39)begin
        img_reg_array_37_60_real <= _zz_186;
      end
      if(_zz_40)begin
        img_reg_array_38_60_real <= _zz_186;
      end
      if(_zz_41)begin
        img_reg_array_39_60_real <= _zz_186;
      end
      if(_zz_42)begin
        img_reg_array_40_60_real <= _zz_186;
      end
      if(_zz_43)begin
        img_reg_array_41_60_real <= _zz_186;
      end
      if(_zz_44)begin
        img_reg_array_42_60_real <= _zz_186;
      end
      if(_zz_45)begin
        img_reg_array_43_60_real <= _zz_186;
      end
      if(_zz_46)begin
        img_reg_array_44_60_real <= _zz_186;
      end
      if(_zz_47)begin
        img_reg_array_45_60_real <= _zz_186;
      end
      if(_zz_48)begin
        img_reg_array_46_60_real <= _zz_186;
      end
      if(_zz_49)begin
        img_reg_array_47_60_real <= _zz_186;
      end
      if(_zz_50)begin
        img_reg_array_48_60_real <= _zz_186;
      end
      if(_zz_51)begin
        img_reg_array_49_60_real <= _zz_186;
      end
      if(_zz_52)begin
        img_reg_array_50_60_real <= _zz_186;
      end
      if(_zz_53)begin
        img_reg_array_51_60_real <= _zz_186;
      end
      if(_zz_54)begin
        img_reg_array_52_60_real <= _zz_186;
      end
      if(_zz_55)begin
        img_reg_array_53_60_real <= _zz_186;
      end
      if(_zz_56)begin
        img_reg_array_54_60_real <= _zz_186;
      end
      if(_zz_57)begin
        img_reg_array_55_60_real <= _zz_186;
      end
      if(_zz_58)begin
        img_reg_array_56_60_real <= _zz_186;
      end
      if(_zz_59)begin
        img_reg_array_57_60_real <= _zz_186;
      end
      if(_zz_60)begin
        img_reg_array_58_60_real <= _zz_186;
      end
      if(_zz_61)begin
        img_reg_array_59_60_real <= _zz_186;
      end
      if(_zz_62)begin
        img_reg_array_60_60_real <= _zz_186;
      end
      if(_zz_63)begin
        img_reg_array_61_60_real <= _zz_186;
      end
      if(_zz_64)begin
        img_reg_array_62_60_real <= _zz_186;
      end
      if(_zz_65)begin
        img_reg_array_63_60_real <= _zz_186;
      end
      if(_zz_2)begin
        img_reg_array_0_60_imag <= _zz_187;
      end
      if(_zz_3)begin
        img_reg_array_1_60_imag <= _zz_187;
      end
      if(_zz_4)begin
        img_reg_array_2_60_imag <= _zz_187;
      end
      if(_zz_5)begin
        img_reg_array_3_60_imag <= _zz_187;
      end
      if(_zz_6)begin
        img_reg_array_4_60_imag <= _zz_187;
      end
      if(_zz_7)begin
        img_reg_array_5_60_imag <= _zz_187;
      end
      if(_zz_8)begin
        img_reg_array_6_60_imag <= _zz_187;
      end
      if(_zz_9)begin
        img_reg_array_7_60_imag <= _zz_187;
      end
      if(_zz_10)begin
        img_reg_array_8_60_imag <= _zz_187;
      end
      if(_zz_11)begin
        img_reg_array_9_60_imag <= _zz_187;
      end
      if(_zz_12)begin
        img_reg_array_10_60_imag <= _zz_187;
      end
      if(_zz_13)begin
        img_reg_array_11_60_imag <= _zz_187;
      end
      if(_zz_14)begin
        img_reg_array_12_60_imag <= _zz_187;
      end
      if(_zz_15)begin
        img_reg_array_13_60_imag <= _zz_187;
      end
      if(_zz_16)begin
        img_reg_array_14_60_imag <= _zz_187;
      end
      if(_zz_17)begin
        img_reg_array_15_60_imag <= _zz_187;
      end
      if(_zz_18)begin
        img_reg_array_16_60_imag <= _zz_187;
      end
      if(_zz_19)begin
        img_reg_array_17_60_imag <= _zz_187;
      end
      if(_zz_20)begin
        img_reg_array_18_60_imag <= _zz_187;
      end
      if(_zz_21)begin
        img_reg_array_19_60_imag <= _zz_187;
      end
      if(_zz_22)begin
        img_reg_array_20_60_imag <= _zz_187;
      end
      if(_zz_23)begin
        img_reg_array_21_60_imag <= _zz_187;
      end
      if(_zz_24)begin
        img_reg_array_22_60_imag <= _zz_187;
      end
      if(_zz_25)begin
        img_reg_array_23_60_imag <= _zz_187;
      end
      if(_zz_26)begin
        img_reg_array_24_60_imag <= _zz_187;
      end
      if(_zz_27)begin
        img_reg_array_25_60_imag <= _zz_187;
      end
      if(_zz_28)begin
        img_reg_array_26_60_imag <= _zz_187;
      end
      if(_zz_29)begin
        img_reg_array_27_60_imag <= _zz_187;
      end
      if(_zz_30)begin
        img_reg_array_28_60_imag <= _zz_187;
      end
      if(_zz_31)begin
        img_reg_array_29_60_imag <= _zz_187;
      end
      if(_zz_32)begin
        img_reg_array_30_60_imag <= _zz_187;
      end
      if(_zz_33)begin
        img_reg_array_31_60_imag <= _zz_187;
      end
      if(_zz_34)begin
        img_reg_array_32_60_imag <= _zz_187;
      end
      if(_zz_35)begin
        img_reg_array_33_60_imag <= _zz_187;
      end
      if(_zz_36)begin
        img_reg_array_34_60_imag <= _zz_187;
      end
      if(_zz_37)begin
        img_reg_array_35_60_imag <= _zz_187;
      end
      if(_zz_38)begin
        img_reg_array_36_60_imag <= _zz_187;
      end
      if(_zz_39)begin
        img_reg_array_37_60_imag <= _zz_187;
      end
      if(_zz_40)begin
        img_reg_array_38_60_imag <= _zz_187;
      end
      if(_zz_41)begin
        img_reg_array_39_60_imag <= _zz_187;
      end
      if(_zz_42)begin
        img_reg_array_40_60_imag <= _zz_187;
      end
      if(_zz_43)begin
        img_reg_array_41_60_imag <= _zz_187;
      end
      if(_zz_44)begin
        img_reg_array_42_60_imag <= _zz_187;
      end
      if(_zz_45)begin
        img_reg_array_43_60_imag <= _zz_187;
      end
      if(_zz_46)begin
        img_reg_array_44_60_imag <= _zz_187;
      end
      if(_zz_47)begin
        img_reg_array_45_60_imag <= _zz_187;
      end
      if(_zz_48)begin
        img_reg_array_46_60_imag <= _zz_187;
      end
      if(_zz_49)begin
        img_reg_array_47_60_imag <= _zz_187;
      end
      if(_zz_50)begin
        img_reg_array_48_60_imag <= _zz_187;
      end
      if(_zz_51)begin
        img_reg_array_49_60_imag <= _zz_187;
      end
      if(_zz_52)begin
        img_reg_array_50_60_imag <= _zz_187;
      end
      if(_zz_53)begin
        img_reg_array_51_60_imag <= _zz_187;
      end
      if(_zz_54)begin
        img_reg_array_52_60_imag <= _zz_187;
      end
      if(_zz_55)begin
        img_reg_array_53_60_imag <= _zz_187;
      end
      if(_zz_56)begin
        img_reg_array_54_60_imag <= _zz_187;
      end
      if(_zz_57)begin
        img_reg_array_55_60_imag <= _zz_187;
      end
      if(_zz_58)begin
        img_reg_array_56_60_imag <= _zz_187;
      end
      if(_zz_59)begin
        img_reg_array_57_60_imag <= _zz_187;
      end
      if(_zz_60)begin
        img_reg_array_58_60_imag <= _zz_187;
      end
      if(_zz_61)begin
        img_reg_array_59_60_imag <= _zz_187;
      end
      if(_zz_62)begin
        img_reg_array_60_60_imag <= _zz_187;
      end
      if(_zz_63)begin
        img_reg_array_61_60_imag <= _zz_187;
      end
      if(_zz_64)begin
        img_reg_array_62_60_imag <= _zz_187;
      end
      if(_zz_65)begin
        img_reg_array_63_60_imag <= _zz_187;
      end
      if(_zz_2)begin
        img_reg_array_0_61_real <= _zz_188;
      end
      if(_zz_3)begin
        img_reg_array_1_61_real <= _zz_188;
      end
      if(_zz_4)begin
        img_reg_array_2_61_real <= _zz_188;
      end
      if(_zz_5)begin
        img_reg_array_3_61_real <= _zz_188;
      end
      if(_zz_6)begin
        img_reg_array_4_61_real <= _zz_188;
      end
      if(_zz_7)begin
        img_reg_array_5_61_real <= _zz_188;
      end
      if(_zz_8)begin
        img_reg_array_6_61_real <= _zz_188;
      end
      if(_zz_9)begin
        img_reg_array_7_61_real <= _zz_188;
      end
      if(_zz_10)begin
        img_reg_array_8_61_real <= _zz_188;
      end
      if(_zz_11)begin
        img_reg_array_9_61_real <= _zz_188;
      end
      if(_zz_12)begin
        img_reg_array_10_61_real <= _zz_188;
      end
      if(_zz_13)begin
        img_reg_array_11_61_real <= _zz_188;
      end
      if(_zz_14)begin
        img_reg_array_12_61_real <= _zz_188;
      end
      if(_zz_15)begin
        img_reg_array_13_61_real <= _zz_188;
      end
      if(_zz_16)begin
        img_reg_array_14_61_real <= _zz_188;
      end
      if(_zz_17)begin
        img_reg_array_15_61_real <= _zz_188;
      end
      if(_zz_18)begin
        img_reg_array_16_61_real <= _zz_188;
      end
      if(_zz_19)begin
        img_reg_array_17_61_real <= _zz_188;
      end
      if(_zz_20)begin
        img_reg_array_18_61_real <= _zz_188;
      end
      if(_zz_21)begin
        img_reg_array_19_61_real <= _zz_188;
      end
      if(_zz_22)begin
        img_reg_array_20_61_real <= _zz_188;
      end
      if(_zz_23)begin
        img_reg_array_21_61_real <= _zz_188;
      end
      if(_zz_24)begin
        img_reg_array_22_61_real <= _zz_188;
      end
      if(_zz_25)begin
        img_reg_array_23_61_real <= _zz_188;
      end
      if(_zz_26)begin
        img_reg_array_24_61_real <= _zz_188;
      end
      if(_zz_27)begin
        img_reg_array_25_61_real <= _zz_188;
      end
      if(_zz_28)begin
        img_reg_array_26_61_real <= _zz_188;
      end
      if(_zz_29)begin
        img_reg_array_27_61_real <= _zz_188;
      end
      if(_zz_30)begin
        img_reg_array_28_61_real <= _zz_188;
      end
      if(_zz_31)begin
        img_reg_array_29_61_real <= _zz_188;
      end
      if(_zz_32)begin
        img_reg_array_30_61_real <= _zz_188;
      end
      if(_zz_33)begin
        img_reg_array_31_61_real <= _zz_188;
      end
      if(_zz_34)begin
        img_reg_array_32_61_real <= _zz_188;
      end
      if(_zz_35)begin
        img_reg_array_33_61_real <= _zz_188;
      end
      if(_zz_36)begin
        img_reg_array_34_61_real <= _zz_188;
      end
      if(_zz_37)begin
        img_reg_array_35_61_real <= _zz_188;
      end
      if(_zz_38)begin
        img_reg_array_36_61_real <= _zz_188;
      end
      if(_zz_39)begin
        img_reg_array_37_61_real <= _zz_188;
      end
      if(_zz_40)begin
        img_reg_array_38_61_real <= _zz_188;
      end
      if(_zz_41)begin
        img_reg_array_39_61_real <= _zz_188;
      end
      if(_zz_42)begin
        img_reg_array_40_61_real <= _zz_188;
      end
      if(_zz_43)begin
        img_reg_array_41_61_real <= _zz_188;
      end
      if(_zz_44)begin
        img_reg_array_42_61_real <= _zz_188;
      end
      if(_zz_45)begin
        img_reg_array_43_61_real <= _zz_188;
      end
      if(_zz_46)begin
        img_reg_array_44_61_real <= _zz_188;
      end
      if(_zz_47)begin
        img_reg_array_45_61_real <= _zz_188;
      end
      if(_zz_48)begin
        img_reg_array_46_61_real <= _zz_188;
      end
      if(_zz_49)begin
        img_reg_array_47_61_real <= _zz_188;
      end
      if(_zz_50)begin
        img_reg_array_48_61_real <= _zz_188;
      end
      if(_zz_51)begin
        img_reg_array_49_61_real <= _zz_188;
      end
      if(_zz_52)begin
        img_reg_array_50_61_real <= _zz_188;
      end
      if(_zz_53)begin
        img_reg_array_51_61_real <= _zz_188;
      end
      if(_zz_54)begin
        img_reg_array_52_61_real <= _zz_188;
      end
      if(_zz_55)begin
        img_reg_array_53_61_real <= _zz_188;
      end
      if(_zz_56)begin
        img_reg_array_54_61_real <= _zz_188;
      end
      if(_zz_57)begin
        img_reg_array_55_61_real <= _zz_188;
      end
      if(_zz_58)begin
        img_reg_array_56_61_real <= _zz_188;
      end
      if(_zz_59)begin
        img_reg_array_57_61_real <= _zz_188;
      end
      if(_zz_60)begin
        img_reg_array_58_61_real <= _zz_188;
      end
      if(_zz_61)begin
        img_reg_array_59_61_real <= _zz_188;
      end
      if(_zz_62)begin
        img_reg_array_60_61_real <= _zz_188;
      end
      if(_zz_63)begin
        img_reg_array_61_61_real <= _zz_188;
      end
      if(_zz_64)begin
        img_reg_array_62_61_real <= _zz_188;
      end
      if(_zz_65)begin
        img_reg_array_63_61_real <= _zz_188;
      end
      if(_zz_2)begin
        img_reg_array_0_61_imag <= _zz_189;
      end
      if(_zz_3)begin
        img_reg_array_1_61_imag <= _zz_189;
      end
      if(_zz_4)begin
        img_reg_array_2_61_imag <= _zz_189;
      end
      if(_zz_5)begin
        img_reg_array_3_61_imag <= _zz_189;
      end
      if(_zz_6)begin
        img_reg_array_4_61_imag <= _zz_189;
      end
      if(_zz_7)begin
        img_reg_array_5_61_imag <= _zz_189;
      end
      if(_zz_8)begin
        img_reg_array_6_61_imag <= _zz_189;
      end
      if(_zz_9)begin
        img_reg_array_7_61_imag <= _zz_189;
      end
      if(_zz_10)begin
        img_reg_array_8_61_imag <= _zz_189;
      end
      if(_zz_11)begin
        img_reg_array_9_61_imag <= _zz_189;
      end
      if(_zz_12)begin
        img_reg_array_10_61_imag <= _zz_189;
      end
      if(_zz_13)begin
        img_reg_array_11_61_imag <= _zz_189;
      end
      if(_zz_14)begin
        img_reg_array_12_61_imag <= _zz_189;
      end
      if(_zz_15)begin
        img_reg_array_13_61_imag <= _zz_189;
      end
      if(_zz_16)begin
        img_reg_array_14_61_imag <= _zz_189;
      end
      if(_zz_17)begin
        img_reg_array_15_61_imag <= _zz_189;
      end
      if(_zz_18)begin
        img_reg_array_16_61_imag <= _zz_189;
      end
      if(_zz_19)begin
        img_reg_array_17_61_imag <= _zz_189;
      end
      if(_zz_20)begin
        img_reg_array_18_61_imag <= _zz_189;
      end
      if(_zz_21)begin
        img_reg_array_19_61_imag <= _zz_189;
      end
      if(_zz_22)begin
        img_reg_array_20_61_imag <= _zz_189;
      end
      if(_zz_23)begin
        img_reg_array_21_61_imag <= _zz_189;
      end
      if(_zz_24)begin
        img_reg_array_22_61_imag <= _zz_189;
      end
      if(_zz_25)begin
        img_reg_array_23_61_imag <= _zz_189;
      end
      if(_zz_26)begin
        img_reg_array_24_61_imag <= _zz_189;
      end
      if(_zz_27)begin
        img_reg_array_25_61_imag <= _zz_189;
      end
      if(_zz_28)begin
        img_reg_array_26_61_imag <= _zz_189;
      end
      if(_zz_29)begin
        img_reg_array_27_61_imag <= _zz_189;
      end
      if(_zz_30)begin
        img_reg_array_28_61_imag <= _zz_189;
      end
      if(_zz_31)begin
        img_reg_array_29_61_imag <= _zz_189;
      end
      if(_zz_32)begin
        img_reg_array_30_61_imag <= _zz_189;
      end
      if(_zz_33)begin
        img_reg_array_31_61_imag <= _zz_189;
      end
      if(_zz_34)begin
        img_reg_array_32_61_imag <= _zz_189;
      end
      if(_zz_35)begin
        img_reg_array_33_61_imag <= _zz_189;
      end
      if(_zz_36)begin
        img_reg_array_34_61_imag <= _zz_189;
      end
      if(_zz_37)begin
        img_reg_array_35_61_imag <= _zz_189;
      end
      if(_zz_38)begin
        img_reg_array_36_61_imag <= _zz_189;
      end
      if(_zz_39)begin
        img_reg_array_37_61_imag <= _zz_189;
      end
      if(_zz_40)begin
        img_reg_array_38_61_imag <= _zz_189;
      end
      if(_zz_41)begin
        img_reg_array_39_61_imag <= _zz_189;
      end
      if(_zz_42)begin
        img_reg_array_40_61_imag <= _zz_189;
      end
      if(_zz_43)begin
        img_reg_array_41_61_imag <= _zz_189;
      end
      if(_zz_44)begin
        img_reg_array_42_61_imag <= _zz_189;
      end
      if(_zz_45)begin
        img_reg_array_43_61_imag <= _zz_189;
      end
      if(_zz_46)begin
        img_reg_array_44_61_imag <= _zz_189;
      end
      if(_zz_47)begin
        img_reg_array_45_61_imag <= _zz_189;
      end
      if(_zz_48)begin
        img_reg_array_46_61_imag <= _zz_189;
      end
      if(_zz_49)begin
        img_reg_array_47_61_imag <= _zz_189;
      end
      if(_zz_50)begin
        img_reg_array_48_61_imag <= _zz_189;
      end
      if(_zz_51)begin
        img_reg_array_49_61_imag <= _zz_189;
      end
      if(_zz_52)begin
        img_reg_array_50_61_imag <= _zz_189;
      end
      if(_zz_53)begin
        img_reg_array_51_61_imag <= _zz_189;
      end
      if(_zz_54)begin
        img_reg_array_52_61_imag <= _zz_189;
      end
      if(_zz_55)begin
        img_reg_array_53_61_imag <= _zz_189;
      end
      if(_zz_56)begin
        img_reg_array_54_61_imag <= _zz_189;
      end
      if(_zz_57)begin
        img_reg_array_55_61_imag <= _zz_189;
      end
      if(_zz_58)begin
        img_reg_array_56_61_imag <= _zz_189;
      end
      if(_zz_59)begin
        img_reg_array_57_61_imag <= _zz_189;
      end
      if(_zz_60)begin
        img_reg_array_58_61_imag <= _zz_189;
      end
      if(_zz_61)begin
        img_reg_array_59_61_imag <= _zz_189;
      end
      if(_zz_62)begin
        img_reg_array_60_61_imag <= _zz_189;
      end
      if(_zz_63)begin
        img_reg_array_61_61_imag <= _zz_189;
      end
      if(_zz_64)begin
        img_reg_array_62_61_imag <= _zz_189;
      end
      if(_zz_65)begin
        img_reg_array_63_61_imag <= _zz_189;
      end
      if(_zz_2)begin
        img_reg_array_0_62_real <= _zz_190;
      end
      if(_zz_3)begin
        img_reg_array_1_62_real <= _zz_190;
      end
      if(_zz_4)begin
        img_reg_array_2_62_real <= _zz_190;
      end
      if(_zz_5)begin
        img_reg_array_3_62_real <= _zz_190;
      end
      if(_zz_6)begin
        img_reg_array_4_62_real <= _zz_190;
      end
      if(_zz_7)begin
        img_reg_array_5_62_real <= _zz_190;
      end
      if(_zz_8)begin
        img_reg_array_6_62_real <= _zz_190;
      end
      if(_zz_9)begin
        img_reg_array_7_62_real <= _zz_190;
      end
      if(_zz_10)begin
        img_reg_array_8_62_real <= _zz_190;
      end
      if(_zz_11)begin
        img_reg_array_9_62_real <= _zz_190;
      end
      if(_zz_12)begin
        img_reg_array_10_62_real <= _zz_190;
      end
      if(_zz_13)begin
        img_reg_array_11_62_real <= _zz_190;
      end
      if(_zz_14)begin
        img_reg_array_12_62_real <= _zz_190;
      end
      if(_zz_15)begin
        img_reg_array_13_62_real <= _zz_190;
      end
      if(_zz_16)begin
        img_reg_array_14_62_real <= _zz_190;
      end
      if(_zz_17)begin
        img_reg_array_15_62_real <= _zz_190;
      end
      if(_zz_18)begin
        img_reg_array_16_62_real <= _zz_190;
      end
      if(_zz_19)begin
        img_reg_array_17_62_real <= _zz_190;
      end
      if(_zz_20)begin
        img_reg_array_18_62_real <= _zz_190;
      end
      if(_zz_21)begin
        img_reg_array_19_62_real <= _zz_190;
      end
      if(_zz_22)begin
        img_reg_array_20_62_real <= _zz_190;
      end
      if(_zz_23)begin
        img_reg_array_21_62_real <= _zz_190;
      end
      if(_zz_24)begin
        img_reg_array_22_62_real <= _zz_190;
      end
      if(_zz_25)begin
        img_reg_array_23_62_real <= _zz_190;
      end
      if(_zz_26)begin
        img_reg_array_24_62_real <= _zz_190;
      end
      if(_zz_27)begin
        img_reg_array_25_62_real <= _zz_190;
      end
      if(_zz_28)begin
        img_reg_array_26_62_real <= _zz_190;
      end
      if(_zz_29)begin
        img_reg_array_27_62_real <= _zz_190;
      end
      if(_zz_30)begin
        img_reg_array_28_62_real <= _zz_190;
      end
      if(_zz_31)begin
        img_reg_array_29_62_real <= _zz_190;
      end
      if(_zz_32)begin
        img_reg_array_30_62_real <= _zz_190;
      end
      if(_zz_33)begin
        img_reg_array_31_62_real <= _zz_190;
      end
      if(_zz_34)begin
        img_reg_array_32_62_real <= _zz_190;
      end
      if(_zz_35)begin
        img_reg_array_33_62_real <= _zz_190;
      end
      if(_zz_36)begin
        img_reg_array_34_62_real <= _zz_190;
      end
      if(_zz_37)begin
        img_reg_array_35_62_real <= _zz_190;
      end
      if(_zz_38)begin
        img_reg_array_36_62_real <= _zz_190;
      end
      if(_zz_39)begin
        img_reg_array_37_62_real <= _zz_190;
      end
      if(_zz_40)begin
        img_reg_array_38_62_real <= _zz_190;
      end
      if(_zz_41)begin
        img_reg_array_39_62_real <= _zz_190;
      end
      if(_zz_42)begin
        img_reg_array_40_62_real <= _zz_190;
      end
      if(_zz_43)begin
        img_reg_array_41_62_real <= _zz_190;
      end
      if(_zz_44)begin
        img_reg_array_42_62_real <= _zz_190;
      end
      if(_zz_45)begin
        img_reg_array_43_62_real <= _zz_190;
      end
      if(_zz_46)begin
        img_reg_array_44_62_real <= _zz_190;
      end
      if(_zz_47)begin
        img_reg_array_45_62_real <= _zz_190;
      end
      if(_zz_48)begin
        img_reg_array_46_62_real <= _zz_190;
      end
      if(_zz_49)begin
        img_reg_array_47_62_real <= _zz_190;
      end
      if(_zz_50)begin
        img_reg_array_48_62_real <= _zz_190;
      end
      if(_zz_51)begin
        img_reg_array_49_62_real <= _zz_190;
      end
      if(_zz_52)begin
        img_reg_array_50_62_real <= _zz_190;
      end
      if(_zz_53)begin
        img_reg_array_51_62_real <= _zz_190;
      end
      if(_zz_54)begin
        img_reg_array_52_62_real <= _zz_190;
      end
      if(_zz_55)begin
        img_reg_array_53_62_real <= _zz_190;
      end
      if(_zz_56)begin
        img_reg_array_54_62_real <= _zz_190;
      end
      if(_zz_57)begin
        img_reg_array_55_62_real <= _zz_190;
      end
      if(_zz_58)begin
        img_reg_array_56_62_real <= _zz_190;
      end
      if(_zz_59)begin
        img_reg_array_57_62_real <= _zz_190;
      end
      if(_zz_60)begin
        img_reg_array_58_62_real <= _zz_190;
      end
      if(_zz_61)begin
        img_reg_array_59_62_real <= _zz_190;
      end
      if(_zz_62)begin
        img_reg_array_60_62_real <= _zz_190;
      end
      if(_zz_63)begin
        img_reg_array_61_62_real <= _zz_190;
      end
      if(_zz_64)begin
        img_reg_array_62_62_real <= _zz_190;
      end
      if(_zz_65)begin
        img_reg_array_63_62_real <= _zz_190;
      end
      if(_zz_2)begin
        img_reg_array_0_62_imag <= _zz_191;
      end
      if(_zz_3)begin
        img_reg_array_1_62_imag <= _zz_191;
      end
      if(_zz_4)begin
        img_reg_array_2_62_imag <= _zz_191;
      end
      if(_zz_5)begin
        img_reg_array_3_62_imag <= _zz_191;
      end
      if(_zz_6)begin
        img_reg_array_4_62_imag <= _zz_191;
      end
      if(_zz_7)begin
        img_reg_array_5_62_imag <= _zz_191;
      end
      if(_zz_8)begin
        img_reg_array_6_62_imag <= _zz_191;
      end
      if(_zz_9)begin
        img_reg_array_7_62_imag <= _zz_191;
      end
      if(_zz_10)begin
        img_reg_array_8_62_imag <= _zz_191;
      end
      if(_zz_11)begin
        img_reg_array_9_62_imag <= _zz_191;
      end
      if(_zz_12)begin
        img_reg_array_10_62_imag <= _zz_191;
      end
      if(_zz_13)begin
        img_reg_array_11_62_imag <= _zz_191;
      end
      if(_zz_14)begin
        img_reg_array_12_62_imag <= _zz_191;
      end
      if(_zz_15)begin
        img_reg_array_13_62_imag <= _zz_191;
      end
      if(_zz_16)begin
        img_reg_array_14_62_imag <= _zz_191;
      end
      if(_zz_17)begin
        img_reg_array_15_62_imag <= _zz_191;
      end
      if(_zz_18)begin
        img_reg_array_16_62_imag <= _zz_191;
      end
      if(_zz_19)begin
        img_reg_array_17_62_imag <= _zz_191;
      end
      if(_zz_20)begin
        img_reg_array_18_62_imag <= _zz_191;
      end
      if(_zz_21)begin
        img_reg_array_19_62_imag <= _zz_191;
      end
      if(_zz_22)begin
        img_reg_array_20_62_imag <= _zz_191;
      end
      if(_zz_23)begin
        img_reg_array_21_62_imag <= _zz_191;
      end
      if(_zz_24)begin
        img_reg_array_22_62_imag <= _zz_191;
      end
      if(_zz_25)begin
        img_reg_array_23_62_imag <= _zz_191;
      end
      if(_zz_26)begin
        img_reg_array_24_62_imag <= _zz_191;
      end
      if(_zz_27)begin
        img_reg_array_25_62_imag <= _zz_191;
      end
      if(_zz_28)begin
        img_reg_array_26_62_imag <= _zz_191;
      end
      if(_zz_29)begin
        img_reg_array_27_62_imag <= _zz_191;
      end
      if(_zz_30)begin
        img_reg_array_28_62_imag <= _zz_191;
      end
      if(_zz_31)begin
        img_reg_array_29_62_imag <= _zz_191;
      end
      if(_zz_32)begin
        img_reg_array_30_62_imag <= _zz_191;
      end
      if(_zz_33)begin
        img_reg_array_31_62_imag <= _zz_191;
      end
      if(_zz_34)begin
        img_reg_array_32_62_imag <= _zz_191;
      end
      if(_zz_35)begin
        img_reg_array_33_62_imag <= _zz_191;
      end
      if(_zz_36)begin
        img_reg_array_34_62_imag <= _zz_191;
      end
      if(_zz_37)begin
        img_reg_array_35_62_imag <= _zz_191;
      end
      if(_zz_38)begin
        img_reg_array_36_62_imag <= _zz_191;
      end
      if(_zz_39)begin
        img_reg_array_37_62_imag <= _zz_191;
      end
      if(_zz_40)begin
        img_reg_array_38_62_imag <= _zz_191;
      end
      if(_zz_41)begin
        img_reg_array_39_62_imag <= _zz_191;
      end
      if(_zz_42)begin
        img_reg_array_40_62_imag <= _zz_191;
      end
      if(_zz_43)begin
        img_reg_array_41_62_imag <= _zz_191;
      end
      if(_zz_44)begin
        img_reg_array_42_62_imag <= _zz_191;
      end
      if(_zz_45)begin
        img_reg_array_43_62_imag <= _zz_191;
      end
      if(_zz_46)begin
        img_reg_array_44_62_imag <= _zz_191;
      end
      if(_zz_47)begin
        img_reg_array_45_62_imag <= _zz_191;
      end
      if(_zz_48)begin
        img_reg_array_46_62_imag <= _zz_191;
      end
      if(_zz_49)begin
        img_reg_array_47_62_imag <= _zz_191;
      end
      if(_zz_50)begin
        img_reg_array_48_62_imag <= _zz_191;
      end
      if(_zz_51)begin
        img_reg_array_49_62_imag <= _zz_191;
      end
      if(_zz_52)begin
        img_reg_array_50_62_imag <= _zz_191;
      end
      if(_zz_53)begin
        img_reg_array_51_62_imag <= _zz_191;
      end
      if(_zz_54)begin
        img_reg_array_52_62_imag <= _zz_191;
      end
      if(_zz_55)begin
        img_reg_array_53_62_imag <= _zz_191;
      end
      if(_zz_56)begin
        img_reg_array_54_62_imag <= _zz_191;
      end
      if(_zz_57)begin
        img_reg_array_55_62_imag <= _zz_191;
      end
      if(_zz_58)begin
        img_reg_array_56_62_imag <= _zz_191;
      end
      if(_zz_59)begin
        img_reg_array_57_62_imag <= _zz_191;
      end
      if(_zz_60)begin
        img_reg_array_58_62_imag <= _zz_191;
      end
      if(_zz_61)begin
        img_reg_array_59_62_imag <= _zz_191;
      end
      if(_zz_62)begin
        img_reg_array_60_62_imag <= _zz_191;
      end
      if(_zz_63)begin
        img_reg_array_61_62_imag <= _zz_191;
      end
      if(_zz_64)begin
        img_reg_array_62_62_imag <= _zz_191;
      end
      if(_zz_65)begin
        img_reg_array_63_62_imag <= _zz_191;
      end
      if(_zz_2)begin
        img_reg_array_0_63_real <= _zz_192;
      end
      if(_zz_3)begin
        img_reg_array_1_63_real <= _zz_192;
      end
      if(_zz_4)begin
        img_reg_array_2_63_real <= _zz_192;
      end
      if(_zz_5)begin
        img_reg_array_3_63_real <= _zz_192;
      end
      if(_zz_6)begin
        img_reg_array_4_63_real <= _zz_192;
      end
      if(_zz_7)begin
        img_reg_array_5_63_real <= _zz_192;
      end
      if(_zz_8)begin
        img_reg_array_6_63_real <= _zz_192;
      end
      if(_zz_9)begin
        img_reg_array_7_63_real <= _zz_192;
      end
      if(_zz_10)begin
        img_reg_array_8_63_real <= _zz_192;
      end
      if(_zz_11)begin
        img_reg_array_9_63_real <= _zz_192;
      end
      if(_zz_12)begin
        img_reg_array_10_63_real <= _zz_192;
      end
      if(_zz_13)begin
        img_reg_array_11_63_real <= _zz_192;
      end
      if(_zz_14)begin
        img_reg_array_12_63_real <= _zz_192;
      end
      if(_zz_15)begin
        img_reg_array_13_63_real <= _zz_192;
      end
      if(_zz_16)begin
        img_reg_array_14_63_real <= _zz_192;
      end
      if(_zz_17)begin
        img_reg_array_15_63_real <= _zz_192;
      end
      if(_zz_18)begin
        img_reg_array_16_63_real <= _zz_192;
      end
      if(_zz_19)begin
        img_reg_array_17_63_real <= _zz_192;
      end
      if(_zz_20)begin
        img_reg_array_18_63_real <= _zz_192;
      end
      if(_zz_21)begin
        img_reg_array_19_63_real <= _zz_192;
      end
      if(_zz_22)begin
        img_reg_array_20_63_real <= _zz_192;
      end
      if(_zz_23)begin
        img_reg_array_21_63_real <= _zz_192;
      end
      if(_zz_24)begin
        img_reg_array_22_63_real <= _zz_192;
      end
      if(_zz_25)begin
        img_reg_array_23_63_real <= _zz_192;
      end
      if(_zz_26)begin
        img_reg_array_24_63_real <= _zz_192;
      end
      if(_zz_27)begin
        img_reg_array_25_63_real <= _zz_192;
      end
      if(_zz_28)begin
        img_reg_array_26_63_real <= _zz_192;
      end
      if(_zz_29)begin
        img_reg_array_27_63_real <= _zz_192;
      end
      if(_zz_30)begin
        img_reg_array_28_63_real <= _zz_192;
      end
      if(_zz_31)begin
        img_reg_array_29_63_real <= _zz_192;
      end
      if(_zz_32)begin
        img_reg_array_30_63_real <= _zz_192;
      end
      if(_zz_33)begin
        img_reg_array_31_63_real <= _zz_192;
      end
      if(_zz_34)begin
        img_reg_array_32_63_real <= _zz_192;
      end
      if(_zz_35)begin
        img_reg_array_33_63_real <= _zz_192;
      end
      if(_zz_36)begin
        img_reg_array_34_63_real <= _zz_192;
      end
      if(_zz_37)begin
        img_reg_array_35_63_real <= _zz_192;
      end
      if(_zz_38)begin
        img_reg_array_36_63_real <= _zz_192;
      end
      if(_zz_39)begin
        img_reg_array_37_63_real <= _zz_192;
      end
      if(_zz_40)begin
        img_reg_array_38_63_real <= _zz_192;
      end
      if(_zz_41)begin
        img_reg_array_39_63_real <= _zz_192;
      end
      if(_zz_42)begin
        img_reg_array_40_63_real <= _zz_192;
      end
      if(_zz_43)begin
        img_reg_array_41_63_real <= _zz_192;
      end
      if(_zz_44)begin
        img_reg_array_42_63_real <= _zz_192;
      end
      if(_zz_45)begin
        img_reg_array_43_63_real <= _zz_192;
      end
      if(_zz_46)begin
        img_reg_array_44_63_real <= _zz_192;
      end
      if(_zz_47)begin
        img_reg_array_45_63_real <= _zz_192;
      end
      if(_zz_48)begin
        img_reg_array_46_63_real <= _zz_192;
      end
      if(_zz_49)begin
        img_reg_array_47_63_real <= _zz_192;
      end
      if(_zz_50)begin
        img_reg_array_48_63_real <= _zz_192;
      end
      if(_zz_51)begin
        img_reg_array_49_63_real <= _zz_192;
      end
      if(_zz_52)begin
        img_reg_array_50_63_real <= _zz_192;
      end
      if(_zz_53)begin
        img_reg_array_51_63_real <= _zz_192;
      end
      if(_zz_54)begin
        img_reg_array_52_63_real <= _zz_192;
      end
      if(_zz_55)begin
        img_reg_array_53_63_real <= _zz_192;
      end
      if(_zz_56)begin
        img_reg_array_54_63_real <= _zz_192;
      end
      if(_zz_57)begin
        img_reg_array_55_63_real <= _zz_192;
      end
      if(_zz_58)begin
        img_reg_array_56_63_real <= _zz_192;
      end
      if(_zz_59)begin
        img_reg_array_57_63_real <= _zz_192;
      end
      if(_zz_60)begin
        img_reg_array_58_63_real <= _zz_192;
      end
      if(_zz_61)begin
        img_reg_array_59_63_real <= _zz_192;
      end
      if(_zz_62)begin
        img_reg_array_60_63_real <= _zz_192;
      end
      if(_zz_63)begin
        img_reg_array_61_63_real <= _zz_192;
      end
      if(_zz_64)begin
        img_reg_array_62_63_real <= _zz_192;
      end
      if(_zz_65)begin
        img_reg_array_63_63_real <= _zz_192;
      end
      if(_zz_2)begin
        img_reg_array_0_63_imag <= _zz_193;
      end
      if(_zz_3)begin
        img_reg_array_1_63_imag <= _zz_193;
      end
      if(_zz_4)begin
        img_reg_array_2_63_imag <= _zz_193;
      end
      if(_zz_5)begin
        img_reg_array_3_63_imag <= _zz_193;
      end
      if(_zz_6)begin
        img_reg_array_4_63_imag <= _zz_193;
      end
      if(_zz_7)begin
        img_reg_array_5_63_imag <= _zz_193;
      end
      if(_zz_8)begin
        img_reg_array_6_63_imag <= _zz_193;
      end
      if(_zz_9)begin
        img_reg_array_7_63_imag <= _zz_193;
      end
      if(_zz_10)begin
        img_reg_array_8_63_imag <= _zz_193;
      end
      if(_zz_11)begin
        img_reg_array_9_63_imag <= _zz_193;
      end
      if(_zz_12)begin
        img_reg_array_10_63_imag <= _zz_193;
      end
      if(_zz_13)begin
        img_reg_array_11_63_imag <= _zz_193;
      end
      if(_zz_14)begin
        img_reg_array_12_63_imag <= _zz_193;
      end
      if(_zz_15)begin
        img_reg_array_13_63_imag <= _zz_193;
      end
      if(_zz_16)begin
        img_reg_array_14_63_imag <= _zz_193;
      end
      if(_zz_17)begin
        img_reg_array_15_63_imag <= _zz_193;
      end
      if(_zz_18)begin
        img_reg_array_16_63_imag <= _zz_193;
      end
      if(_zz_19)begin
        img_reg_array_17_63_imag <= _zz_193;
      end
      if(_zz_20)begin
        img_reg_array_18_63_imag <= _zz_193;
      end
      if(_zz_21)begin
        img_reg_array_19_63_imag <= _zz_193;
      end
      if(_zz_22)begin
        img_reg_array_20_63_imag <= _zz_193;
      end
      if(_zz_23)begin
        img_reg_array_21_63_imag <= _zz_193;
      end
      if(_zz_24)begin
        img_reg_array_22_63_imag <= _zz_193;
      end
      if(_zz_25)begin
        img_reg_array_23_63_imag <= _zz_193;
      end
      if(_zz_26)begin
        img_reg_array_24_63_imag <= _zz_193;
      end
      if(_zz_27)begin
        img_reg_array_25_63_imag <= _zz_193;
      end
      if(_zz_28)begin
        img_reg_array_26_63_imag <= _zz_193;
      end
      if(_zz_29)begin
        img_reg_array_27_63_imag <= _zz_193;
      end
      if(_zz_30)begin
        img_reg_array_28_63_imag <= _zz_193;
      end
      if(_zz_31)begin
        img_reg_array_29_63_imag <= _zz_193;
      end
      if(_zz_32)begin
        img_reg_array_30_63_imag <= _zz_193;
      end
      if(_zz_33)begin
        img_reg_array_31_63_imag <= _zz_193;
      end
      if(_zz_34)begin
        img_reg_array_32_63_imag <= _zz_193;
      end
      if(_zz_35)begin
        img_reg_array_33_63_imag <= _zz_193;
      end
      if(_zz_36)begin
        img_reg_array_34_63_imag <= _zz_193;
      end
      if(_zz_37)begin
        img_reg_array_35_63_imag <= _zz_193;
      end
      if(_zz_38)begin
        img_reg_array_36_63_imag <= _zz_193;
      end
      if(_zz_39)begin
        img_reg_array_37_63_imag <= _zz_193;
      end
      if(_zz_40)begin
        img_reg_array_38_63_imag <= _zz_193;
      end
      if(_zz_41)begin
        img_reg_array_39_63_imag <= _zz_193;
      end
      if(_zz_42)begin
        img_reg_array_40_63_imag <= _zz_193;
      end
      if(_zz_43)begin
        img_reg_array_41_63_imag <= _zz_193;
      end
      if(_zz_44)begin
        img_reg_array_42_63_imag <= _zz_193;
      end
      if(_zz_45)begin
        img_reg_array_43_63_imag <= _zz_193;
      end
      if(_zz_46)begin
        img_reg_array_44_63_imag <= _zz_193;
      end
      if(_zz_47)begin
        img_reg_array_45_63_imag <= _zz_193;
      end
      if(_zz_48)begin
        img_reg_array_46_63_imag <= _zz_193;
      end
      if(_zz_49)begin
        img_reg_array_47_63_imag <= _zz_193;
      end
      if(_zz_50)begin
        img_reg_array_48_63_imag <= _zz_193;
      end
      if(_zz_51)begin
        img_reg_array_49_63_imag <= _zz_193;
      end
      if(_zz_52)begin
        img_reg_array_50_63_imag <= _zz_193;
      end
      if(_zz_53)begin
        img_reg_array_51_63_imag <= _zz_193;
      end
      if(_zz_54)begin
        img_reg_array_52_63_imag <= _zz_193;
      end
      if(_zz_55)begin
        img_reg_array_53_63_imag <= _zz_193;
      end
      if(_zz_56)begin
        img_reg_array_54_63_imag <= _zz_193;
      end
      if(_zz_57)begin
        img_reg_array_55_63_imag <= _zz_193;
      end
      if(_zz_58)begin
        img_reg_array_56_63_imag <= _zz_193;
      end
      if(_zz_59)begin
        img_reg_array_57_63_imag <= _zz_193;
      end
      if(_zz_60)begin
        img_reg_array_58_63_imag <= _zz_193;
      end
      if(_zz_61)begin
        img_reg_array_59_63_imag <= _zz_193;
      end
      if(_zz_62)begin
        img_reg_array_60_63_imag <= _zz_193;
      end
      if(_zz_63)begin
        img_reg_array_61_63_imag <= _zz_193;
      end
      if(_zz_64)begin
        img_reg_array_62_63_imag <= _zz_193;
      end
      if(_zz_65)begin
        img_reg_array_63_63_imag <= _zz_193;
      end
    end
    col_addr <= null_cnt_value;
    myFFT_3_fft_col_out_regNext_payload_0_real <= myFFT_3_fft_col_out_payload_0_real;
    myFFT_3_fft_col_out_regNext_payload_0_imag <= myFFT_3_fft_col_out_payload_0_imag;
    myFFT_3_fft_col_out_regNext_payload_1_real <= myFFT_3_fft_col_out_payload_1_real;
    myFFT_3_fft_col_out_regNext_payload_1_imag <= myFFT_3_fft_col_out_payload_1_imag;
    myFFT_3_fft_col_out_regNext_payload_2_real <= myFFT_3_fft_col_out_payload_2_real;
    myFFT_3_fft_col_out_regNext_payload_2_imag <= myFFT_3_fft_col_out_payload_2_imag;
    myFFT_3_fft_col_out_regNext_payload_3_real <= myFFT_3_fft_col_out_payload_3_real;
    myFFT_3_fft_col_out_regNext_payload_3_imag <= myFFT_3_fft_col_out_payload_3_imag;
    myFFT_3_fft_col_out_regNext_payload_4_real <= myFFT_3_fft_col_out_payload_4_real;
    myFFT_3_fft_col_out_regNext_payload_4_imag <= myFFT_3_fft_col_out_payload_4_imag;
    myFFT_3_fft_col_out_regNext_payload_5_real <= myFFT_3_fft_col_out_payload_5_real;
    myFFT_3_fft_col_out_regNext_payload_5_imag <= myFFT_3_fft_col_out_payload_5_imag;
    myFFT_3_fft_col_out_regNext_payload_6_real <= myFFT_3_fft_col_out_payload_6_real;
    myFFT_3_fft_col_out_regNext_payload_6_imag <= myFFT_3_fft_col_out_payload_6_imag;
    myFFT_3_fft_col_out_regNext_payload_7_real <= myFFT_3_fft_col_out_payload_7_real;
    myFFT_3_fft_col_out_regNext_payload_7_imag <= myFFT_3_fft_col_out_payload_7_imag;
    myFFT_3_fft_col_out_regNext_payload_8_real <= myFFT_3_fft_col_out_payload_8_real;
    myFFT_3_fft_col_out_regNext_payload_8_imag <= myFFT_3_fft_col_out_payload_8_imag;
    myFFT_3_fft_col_out_regNext_payload_9_real <= myFFT_3_fft_col_out_payload_9_real;
    myFFT_3_fft_col_out_regNext_payload_9_imag <= myFFT_3_fft_col_out_payload_9_imag;
    myFFT_3_fft_col_out_regNext_payload_10_real <= myFFT_3_fft_col_out_payload_10_real;
    myFFT_3_fft_col_out_regNext_payload_10_imag <= myFFT_3_fft_col_out_payload_10_imag;
    myFFT_3_fft_col_out_regNext_payload_11_real <= myFFT_3_fft_col_out_payload_11_real;
    myFFT_3_fft_col_out_regNext_payload_11_imag <= myFFT_3_fft_col_out_payload_11_imag;
    myFFT_3_fft_col_out_regNext_payload_12_real <= myFFT_3_fft_col_out_payload_12_real;
    myFFT_3_fft_col_out_regNext_payload_12_imag <= myFFT_3_fft_col_out_payload_12_imag;
    myFFT_3_fft_col_out_regNext_payload_13_real <= myFFT_3_fft_col_out_payload_13_real;
    myFFT_3_fft_col_out_regNext_payload_13_imag <= myFFT_3_fft_col_out_payload_13_imag;
    myFFT_3_fft_col_out_regNext_payload_14_real <= myFFT_3_fft_col_out_payload_14_real;
    myFFT_3_fft_col_out_regNext_payload_14_imag <= myFFT_3_fft_col_out_payload_14_imag;
    myFFT_3_fft_col_out_regNext_payload_15_real <= myFFT_3_fft_col_out_payload_15_real;
    myFFT_3_fft_col_out_regNext_payload_15_imag <= myFFT_3_fft_col_out_payload_15_imag;
    myFFT_3_fft_col_out_regNext_payload_16_real <= myFFT_3_fft_col_out_payload_16_real;
    myFFT_3_fft_col_out_regNext_payload_16_imag <= myFFT_3_fft_col_out_payload_16_imag;
    myFFT_3_fft_col_out_regNext_payload_17_real <= myFFT_3_fft_col_out_payload_17_real;
    myFFT_3_fft_col_out_regNext_payload_17_imag <= myFFT_3_fft_col_out_payload_17_imag;
    myFFT_3_fft_col_out_regNext_payload_18_real <= myFFT_3_fft_col_out_payload_18_real;
    myFFT_3_fft_col_out_regNext_payload_18_imag <= myFFT_3_fft_col_out_payload_18_imag;
    myFFT_3_fft_col_out_regNext_payload_19_real <= myFFT_3_fft_col_out_payload_19_real;
    myFFT_3_fft_col_out_regNext_payload_19_imag <= myFFT_3_fft_col_out_payload_19_imag;
    myFFT_3_fft_col_out_regNext_payload_20_real <= myFFT_3_fft_col_out_payload_20_real;
    myFFT_3_fft_col_out_regNext_payload_20_imag <= myFFT_3_fft_col_out_payload_20_imag;
    myFFT_3_fft_col_out_regNext_payload_21_real <= myFFT_3_fft_col_out_payload_21_real;
    myFFT_3_fft_col_out_regNext_payload_21_imag <= myFFT_3_fft_col_out_payload_21_imag;
    myFFT_3_fft_col_out_regNext_payload_22_real <= myFFT_3_fft_col_out_payload_22_real;
    myFFT_3_fft_col_out_regNext_payload_22_imag <= myFFT_3_fft_col_out_payload_22_imag;
    myFFT_3_fft_col_out_regNext_payload_23_real <= myFFT_3_fft_col_out_payload_23_real;
    myFFT_3_fft_col_out_regNext_payload_23_imag <= myFFT_3_fft_col_out_payload_23_imag;
    myFFT_3_fft_col_out_regNext_payload_24_real <= myFFT_3_fft_col_out_payload_24_real;
    myFFT_3_fft_col_out_regNext_payload_24_imag <= myFFT_3_fft_col_out_payload_24_imag;
    myFFT_3_fft_col_out_regNext_payload_25_real <= myFFT_3_fft_col_out_payload_25_real;
    myFFT_3_fft_col_out_regNext_payload_25_imag <= myFFT_3_fft_col_out_payload_25_imag;
    myFFT_3_fft_col_out_regNext_payload_26_real <= myFFT_3_fft_col_out_payload_26_real;
    myFFT_3_fft_col_out_regNext_payload_26_imag <= myFFT_3_fft_col_out_payload_26_imag;
    myFFT_3_fft_col_out_regNext_payload_27_real <= myFFT_3_fft_col_out_payload_27_real;
    myFFT_3_fft_col_out_regNext_payload_27_imag <= myFFT_3_fft_col_out_payload_27_imag;
    myFFT_3_fft_col_out_regNext_payload_28_real <= myFFT_3_fft_col_out_payload_28_real;
    myFFT_3_fft_col_out_regNext_payload_28_imag <= myFFT_3_fft_col_out_payload_28_imag;
    myFFT_3_fft_col_out_regNext_payload_29_real <= myFFT_3_fft_col_out_payload_29_real;
    myFFT_3_fft_col_out_regNext_payload_29_imag <= myFFT_3_fft_col_out_payload_29_imag;
    myFFT_3_fft_col_out_regNext_payload_30_real <= myFFT_3_fft_col_out_payload_30_real;
    myFFT_3_fft_col_out_regNext_payload_30_imag <= myFFT_3_fft_col_out_payload_30_imag;
    myFFT_3_fft_col_out_regNext_payload_31_real <= myFFT_3_fft_col_out_payload_31_real;
    myFFT_3_fft_col_out_regNext_payload_31_imag <= myFFT_3_fft_col_out_payload_31_imag;
    myFFT_3_fft_col_out_regNext_payload_32_real <= myFFT_3_fft_col_out_payload_32_real;
    myFFT_3_fft_col_out_regNext_payload_32_imag <= myFFT_3_fft_col_out_payload_32_imag;
    myFFT_3_fft_col_out_regNext_payload_33_real <= myFFT_3_fft_col_out_payload_33_real;
    myFFT_3_fft_col_out_regNext_payload_33_imag <= myFFT_3_fft_col_out_payload_33_imag;
    myFFT_3_fft_col_out_regNext_payload_34_real <= myFFT_3_fft_col_out_payload_34_real;
    myFFT_3_fft_col_out_regNext_payload_34_imag <= myFFT_3_fft_col_out_payload_34_imag;
    myFFT_3_fft_col_out_regNext_payload_35_real <= myFFT_3_fft_col_out_payload_35_real;
    myFFT_3_fft_col_out_regNext_payload_35_imag <= myFFT_3_fft_col_out_payload_35_imag;
    myFFT_3_fft_col_out_regNext_payload_36_real <= myFFT_3_fft_col_out_payload_36_real;
    myFFT_3_fft_col_out_regNext_payload_36_imag <= myFFT_3_fft_col_out_payload_36_imag;
    myFFT_3_fft_col_out_regNext_payload_37_real <= myFFT_3_fft_col_out_payload_37_real;
    myFFT_3_fft_col_out_regNext_payload_37_imag <= myFFT_3_fft_col_out_payload_37_imag;
    myFFT_3_fft_col_out_regNext_payload_38_real <= myFFT_3_fft_col_out_payload_38_real;
    myFFT_3_fft_col_out_regNext_payload_38_imag <= myFFT_3_fft_col_out_payload_38_imag;
    myFFT_3_fft_col_out_regNext_payload_39_real <= myFFT_3_fft_col_out_payload_39_real;
    myFFT_3_fft_col_out_regNext_payload_39_imag <= myFFT_3_fft_col_out_payload_39_imag;
    myFFT_3_fft_col_out_regNext_payload_40_real <= myFFT_3_fft_col_out_payload_40_real;
    myFFT_3_fft_col_out_regNext_payload_40_imag <= myFFT_3_fft_col_out_payload_40_imag;
    myFFT_3_fft_col_out_regNext_payload_41_real <= myFFT_3_fft_col_out_payload_41_real;
    myFFT_3_fft_col_out_regNext_payload_41_imag <= myFFT_3_fft_col_out_payload_41_imag;
    myFFT_3_fft_col_out_regNext_payload_42_real <= myFFT_3_fft_col_out_payload_42_real;
    myFFT_3_fft_col_out_regNext_payload_42_imag <= myFFT_3_fft_col_out_payload_42_imag;
    myFFT_3_fft_col_out_regNext_payload_43_real <= myFFT_3_fft_col_out_payload_43_real;
    myFFT_3_fft_col_out_regNext_payload_43_imag <= myFFT_3_fft_col_out_payload_43_imag;
    myFFT_3_fft_col_out_regNext_payload_44_real <= myFFT_3_fft_col_out_payload_44_real;
    myFFT_3_fft_col_out_regNext_payload_44_imag <= myFFT_3_fft_col_out_payload_44_imag;
    myFFT_3_fft_col_out_regNext_payload_45_real <= myFFT_3_fft_col_out_payload_45_real;
    myFFT_3_fft_col_out_regNext_payload_45_imag <= myFFT_3_fft_col_out_payload_45_imag;
    myFFT_3_fft_col_out_regNext_payload_46_real <= myFFT_3_fft_col_out_payload_46_real;
    myFFT_3_fft_col_out_regNext_payload_46_imag <= myFFT_3_fft_col_out_payload_46_imag;
    myFFT_3_fft_col_out_regNext_payload_47_real <= myFFT_3_fft_col_out_payload_47_real;
    myFFT_3_fft_col_out_regNext_payload_47_imag <= myFFT_3_fft_col_out_payload_47_imag;
    myFFT_3_fft_col_out_regNext_payload_48_real <= myFFT_3_fft_col_out_payload_48_real;
    myFFT_3_fft_col_out_regNext_payload_48_imag <= myFFT_3_fft_col_out_payload_48_imag;
    myFFT_3_fft_col_out_regNext_payload_49_real <= myFFT_3_fft_col_out_payload_49_real;
    myFFT_3_fft_col_out_regNext_payload_49_imag <= myFFT_3_fft_col_out_payload_49_imag;
    myFFT_3_fft_col_out_regNext_payload_50_real <= myFFT_3_fft_col_out_payload_50_real;
    myFFT_3_fft_col_out_regNext_payload_50_imag <= myFFT_3_fft_col_out_payload_50_imag;
    myFFT_3_fft_col_out_regNext_payload_51_real <= myFFT_3_fft_col_out_payload_51_real;
    myFFT_3_fft_col_out_regNext_payload_51_imag <= myFFT_3_fft_col_out_payload_51_imag;
    myFFT_3_fft_col_out_regNext_payload_52_real <= myFFT_3_fft_col_out_payload_52_real;
    myFFT_3_fft_col_out_regNext_payload_52_imag <= myFFT_3_fft_col_out_payload_52_imag;
    myFFT_3_fft_col_out_regNext_payload_53_real <= myFFT_3_fft_col_out_payload_53_real;
    myFFT_3_fft_col_out_regNext_payload_53_imag <= myFFT_3_fft_col_out_payload_53_imag;
    myFFT_3_fft_col_out_regNext_payload_54_real <= myFFT_3_fft_col_out_payload_54_real;
    myFFT_3_fft_col_out_regNext_payload_54_imag <= myFFT_3_fft_col_out_payload_54_imag;
    myFFT_3_fft_col_out_regNext_payload_55_real <= myFFT_3_fft_col_out_payload_55_real;
    myFFT_3_fft_col_out_regNext_payload_55_imag <= myFFT_3_fft_col_out_payload_55_imag;
    myFFT_3_fft_col_out_regNext_payload_56_real <= myFFT_3_fft_col_out_payload_56_real;
    myFFT_3_fft_col_out_regNext_payload_56_imag <= myFFT_3_fft_col_out_payload_56_imag;
    myFFT_3_fft_col_out_regNext_payload_57_real <= myFFT_3_fft_col_out_payload_57_real;
    myFFT_3_fft_col_out_regNext_payload_57_imag <= myFFT_3_fft_col_out_payload_57_imag;
    myFFT_3_fft_col_out_regNext_payload_58_real <= myFFT_3_fft_col_out_payload_58_real;
    myFFT_3_fft_col_out_regNext_payload_58_imag <= myFFT_3_fft_col_out_payload_58_imag;
    myFFT_3_fft_col_out_regNext_payload_59_real <= myFFT_3_fft_col_out_payload_59_real;
    myFFT_3_fft_col_out_regNext_payload_59_imag <= myFFT_3_fft_col_out_payload_59_imag;
    myFFT_3_fft_col_out_regNext_payload_60_real <= myFFT_3_fft_col_out_payload_60_real;
    myFFT_3_fft_col_out_regNext_payload_60_imag <= myFFT_3_fft_col_out_payload_60_imag;
    myFFT_3_fft_col_out_regNext_payload_61_real <= myFFT_3_fft_col_out_payload_61_real;
    myFFT_3_fft_col_out_regNext_payload_61_imag <= myFFT_3_fft_col_out_payload_61_imag;
    myFFT_3_fft_col_out_regNext_payload_62_real <= myFFT_3_fft_col_out_payload_62_real;
    myFFT_3_fft_col_out_regNext_payload_62_imag <= myFFT_3_fft_col_out_payload_62_imag;
    myFFT_3_fft_col_out_regNext_payload_63_real <= myFFT_3_fft_col_out_payload_63_real;
    myFFT_3_fft_col_out_regNext_payload_63_imag <= myFFT_3_fft_col_out_payload_63_imag;
  end


endmodule

module MyFFT_1 (
  input               io_data_in_valid,
  input      [17:0]   io_data_in_payload_0_real,
  input      [17:0]   io_data_in_payload_0_imag,
  input      [17:0]   io_data_in_payload_1_real,
  input      [17:0]   io_data_in_payload_1_imag,
  input      [17:0]   io_data_in_payload_2_real,
  input      [17:0]   io_data_in_payload_2_imag,
  input      [17:0]   io_data_in_payload_3_real,
  input      [17:0]   io_data_in_payload_3_imag,
  input      [17:0]   io_data_in_payload_4_real,
  input      [17:0]   io_data_in_payload_4_imag,
  input      [17:0]   io_data_in_payload_5_real,
  input      [17:0]   io_data_in_payload_5_imag,
  input      [17:0]   io_data_in_payload_6_real,
  input      [17:0]   io_data_in_payload_6_imag,
  input      [17:0]   io_data_in_payload_7_real,
  input      [17:0]   io_data_in_payload_7_imag,
  input      [17:0]   io_data_in_payload_8_real,
  input      [17:0]   io_data_in_payload_8_imag,
  input      [17:0]   io_data_in_payload_9_real,
  input      [17:0]   io_data_in_payload_9_imag,
  input      [17:0]   io_data_in_payload_10_real,
  input      [17:0]   io_data_in_payload_10_imag,
  input      [17:0]   io_data_in_payload_11_real,
  input      [17:0]   io_data_in_payload_11_imag,
  input      [17:0]   io_data_in_payload_12_real,
  input      [17:0]   io_data_in_payload_12_imag,
  input      [17:0]   io_data_in_payload_13_real,
  input      [17:0]   io_data_in_payload_13_imag,
  input      [17:0]   io_data_in_payload_14_real,
  input      [17:0]   io_data_in_payload_14_imag,
  input      [17:0]   io_data_in_payload_15_real,
  input      [17:0]   io_data_in_payload_15_imag,
  input      [17:0]   io_data_in_payload_16_real,
  input      [17:0]   io_data_in_payload_16_imag,
  input      [17:0]   io_data_in_payload_17_real,
  input      [17:0]   io_data_in_payload_17_imag,
  input      [17:0]   io_data_in_payload_18_real,
  input      [17:0]   io_data_in_payload_18_imag,
  input      [17:0]   io_data_in_payload_19_real,
  input      [17:0]   io_data_in_payload_19_imag,
  input      [17:0]   io_data_in_payload_20_real,
  input      [17:0]   io_data_in_payload_20_imag,
  input      [17:0]   io_data_in_payload_21_real,
  input      [17:0]   io_data_in_payload_21_imag,
  input      [17:0]   io_data_in_payload_22_real,
  input      [17:0]   io_data_in_payload_22_imag,
  input      [17:0]   io_data_in_payload_23_real,
  input      [17:0]   io_data_in_payload_23_imag,
  input      [17:0]   io_data_in_payload_24_real,
  input      [17:0]   io_data_in_payload_24_imag,
  input      [17:0]   io_data_in_payload_25_real,
  input      [17:0]   io_data_in_payload_25_imag,
  input      [17:0]   io_data_in_payload_26_real,
  input      [17:0]   io_data_in_payload_26_imag,
  input      [17:0]   io_data_in_payload_27_real,
  input      [17:0]   io_data_in_payload_27_imag,
  input      [17:0]   io_data_in_payload_28_real,
  input      [17:0]   io_data_in_payload_28_imag,
  input      [17:0]   io_data_in_payload_29_real,
  input      [17:0]   io_data_in_payload_29_imag,
  input      [17:0]   io_data_in_payload_30_real,
  input      [17:0]   io_data_in_payload_30_imag,
  input      [17:0]   io_data_in_payload_31_real,
  input      [17:0]   io_data_in_payload_31_imag,
  input      [17:0]   io_data_in_payload_32_real,
  input      [17:0]   io_data_in_payload_32_imag,
  input      [17:0]   io_data_in_payload_33_real,
  input      [17:0]   io_data_in_payload_33_imag,
  input      [17:0]   io_data_in_payload_34_real,
  input      [17:0]   io_data_in_payload_34_imag,
  input      [17:0]   io_data_in_payload_35_real,
  input      [17:0]   io_data_in_payload_35_imag,
  input      [17:0]   io_data_in_payload_36_real,
  input      [17:0]   io_data_in_payload_36_imag,
  input      [17:0]   io_data_in_payload_37_real,
  input      [17:0]   io_data_in_payload_37_imag,
  input      [17:0]   io_data_in_payload_38_real,
  input      [17:0]   io_data_in_payload_38_imag,
  input      [17:0]   io_data_in_payload_39_real,
  input      [17:0]   io_data_in_payload_39_imag,
  input      [17:0]   io_data_in_payload_40_real,
  input      [17:0]   io_data_in_payload_40_imag,
  input      [17:0]   io_data_in_payload_41_real,
  input      [17:0]   io_data_in_payload_41_imag,
  input      [17:0]   io_data_in_payload_42_real,
  input      [17:0]   io_data_in_payload_42_imag,
  input      [17:0]   io_data_in_payload_43_real,
  input      [17:0]   io_data_in_payload_43_imag,
  input      [17:0]   io_data_in_payload_44_real,
  input      [17:0]   io_data_in_payload_44_imag,
  input      [17:0]   io_data_in_payload_45_real,
  input      [17:0]   io_data_in_payload_45_imag,
  input      [17:0]   io_data_in_payload_46_real,
  input      [17:0]   io_data_in_payload_46_imag,
  input      [17:0]   io_data_in_payload_47_real,
  input      [17:0]   io_data_in_payload_47_imag,
  input      [17:0]   io_data_in_payload_48_real,
  input      [17:0]   io_data_in_payload_48_imag,
  input      [17:0]   io_data_in_payload_49_real,
  input      [17:0]   io_data_in_payload_49_imag,
  input      [17:0]   io_data_in_payload_50_real,
  input      [17:0]   io_data_in_payload_50_imag,
  input      [17:0]   io_data_in_payload_51_real,
  input      [17:0]   io_data_in_payload_51_imag,
  input      [17:0]   io_data_in_payload_52_real,
  input      [17:0]   io_data_in_payload_52_imag,
  input      [17:0]   io_data_in_payload_53_real,
  input      [17:0]   io_data_in_payload_53_imag,
  input      [17:0]   io_data_in_payload_54_real,
  input      [17:0]   io_data_in_payload_54_imag,
  input      [17:0]   io_data_in_payload_55_real,
  input      [17:0]   io_data_in_payload_55_imag,
  input      [17:0]   io_data_in_payload_56_real,
  input      [17:0]   io_data_in_payload_56_imag,
  input      [17:0]   io_data_in_payload_57_real,
  input      [17:0]   io_data_in_payload_57_imag,
  input      [17:0]   io_data_in_payload_58_real,
  input      [17:0]   io_data_in_payload_58_imag,
  input      [17:0]   io_data_in_payload_59_real,
  input      [17:0]   io_data_in_payload_59_imag,
  input      [17:0]   io_data_in_payload_60_real,
  input      [17:0]   io_data_in_payload_60_imag,
  input      [17:0]   io_data_in_payload_61_real,
  input      [17:0]   io_data_in_payload_61_imag,
  input      [17:0]   io_data_in_payload_62_real,
  input      [17:0]   io_data_in_payload_62_imag,
  input      [17:0]   io_data_in_payload_63_real,
  input      [17:0]   io_data_in_payload_63_imag,
  output              fft_col_out_valid,
  output     [17:0]   fft_col_out_payload_0_real,
  output     [17:0]   fft_col_out_payload_0_imag,
  output     [17:0]   fft_col_out_payload_1_real,
  output     [17:0]   fft_col_out_payload_1_imag,
  output     [17:0]   fft_col_out_payload_2_real,
  output     [17:0]   fft_col_out_payload_2_imag,
  output     [17:0]   fft_col_out_payload_3_real,
  output     [17:0]   fft_col_out_payload_3_imag,
  output     [17:0]   fft_col_out_payload_4_real,
  output     [17:0]   fft_col_out_payload_4_imag,
  output     [17:0]   fft_col_out_payload_5_real,
  output     [17:0]   fft_col_out_payload_5_imag,
  output     [17:0]   fft_col_out_payload_6_real,
  output     [17:0]   fft_col_out_payload_6_imag,
  output     [17:0]   fft_col_out_payload_7_real,
  output     [17:0]   fft_col_out_payload_7_imag,
  output     [17:0]   fft_col_out_payload_8_real,
  output     [17:0]   fft_col_out_payload_8_imag,
  output     [17:0]   fft_col_out_payload_9_real,
  output     [17:0]   fft_col_out_payload_9_imag,
  output     [17:0]   fft_col_out_payload_10_real,
  output     [17:0]   fft_col_out_payload_10_imag,
  output     [17:0]   fft_col_out_payload_11_real,
  output     [17:0]   fft_col_out_payload_11_imag,
  output     [17:0]   fft_col_out_payload_12_real,
  output     [17:0]   fft_col_out_payload_12_imag,
  output     [17:0]   fft_col_out_payload_13_real,
  output     [17:0]   fft_col_out_payload_13_imag,
  output     [17:0]   fft_col_out_payload_14_real,
  output     [17:0]   fft_col_out_payload_14_imag,
  output     [17:0]   fft_col_out_payload_15_real,
  output     [17:0]   fft_col_out_payload_15_imag,
  output     [17:0]   fft_col_out_payload_16_real,
  output     [17:0]   fft_col_out_payload_16_imag,
  output     [17:0]   fft_col_out_payload_17_real,
  output     [17:0]   fft_col_out_payload_17_imag,
  output     [17:0]   fft_col_out_payload_18_real,
  output     [17:0]   fft_col_out_payload_18_imag,
  output     [17:0]   fft_col_out_payload_19_real,
  output     [17:0]   fft_col_out_payload_19_imag,
  output     [17:0]   fft_col_out_payload_20_real,
  output     [17:0]   fft_col_out_payload_20_imag,
  output     [17:0]   fft_col_out_payload_21_real,
  output     [17:0]   fft_col_out_payload_21_imag,
  output     [17:0]   fft_col_out_payload_22_real,
  output     [17:0]   fft_col_out_payload_22_imag,
  output     [17:0]   fft_col_out_payload_23_real,
  output     [17:0]   fft_col_out_payload_23_imag,
  output     [17:0]   fft_col_out_payload_24_real,
  output     [17:0]   fft_col_out_payload_24_imag,
  output     [17:0]   fft_col_out_payload_25_real,
  output     [17:0]   fft_col_out_payload_25_imag,
  output     [17:0]   fft_col_out_payload_26_real,
  output     [17:0]   fft_col_out_payload_26_imag,
  output     [17:0]   fft_col_out_payload_27_real,
  output     [17:0]   fft_col_out_payload_27_imag,
  output     [17:0]   fft_col_out_payload_28_real,
  output     [17:0]   fft_col_out_payload_28_imag,
  output     [17:0]   fft_col_out_payload_29_real,
  output     [17:0]   fft_col_out_payload_29_imag,
  output     [17:0]   fft_col_out_payload_30_real,
  output     [17:0]   fft_col_out_payload_30_imag,
  output     [17:0]   fft_col_out_payload_31_real,
  output     [17:0]   fft_col_out_payload_31_imag,
  output     [17:0]   fft_col_out_payload_32_real,
  output     [17:0]   fft_col_out_payload_32_imag,
  output     [17:0]   fft_col_out_payload_33_real,
  output     [17:0]   fft_col_out_payload_33_imag,
  output     [17:0]   fft_col_out_payload_34_real,
  output     [17:0]   fft_col_out_payload_34_imag,
  output     [17:0]   fft_col_out_payload_35_real,
  output     [17:0]   fft_col_out_payload_35_imag,
  output     [17:0]   fft_col_out_payload_36_real,
  output     [17:0]   fft_col_out_payload_36_imag,
  output     [17:0]   fft_col_out_payload_37_real,
  output     [17:0]   fft_col_out_payload_37_imag,
  output     [17:0]   fft_col_out_payload_38_real,
  output     [17:0]   fft_col_out_payload_38_imag,
  output     [17:0]   fft_col_out_payload_39_real,
  output     [17:0]   fft_col_out_payload_39_imag,
  output     [17:0]   fft_col_out_payload_40_real,
  output     [17:0]   fft_col_out_payload_40_imag,
  output     [17:0]   fft_col_out_payload_41_real,
  output     [17:0]   fft_col_out_payload_41_imag,
  output     [17:0]   fft_col_out_payload_42_real,
  output     [17:0]   fft_col_out_payload_42_imag,
  output     [17:0]   fft_col_out_payload_43_real,
  output     [17:0]   fft_col_out_payload_43_imag,
  output     [17:0]   fft_col_out_payload_44_real,
  output     [17:0]   fft_col_out_payload_44_imag,
  output     [17:0]   fft_col_out_payload_45_real,
  output     [17:0]   fft_col_out_payload_45_imag,
  output     [17:0]   fft_col_out_payload_46_real,
  output     [17:0]   fft_col_out_payload_46_imag,
  output     [17:0]   fft_col_out_payload_47_real,
  output     [17:0]   fft_col_out_payload_47_imag,
  output     [17:0]   fft_col_out_payload_48_real,
  output     [17:0]   fft_col_out_payload_48_imag,
  output     [17:0]   fft_col_out_payload_49_real,
  output     [17:0]   fft_col_out_payload_49_imag,
  output     [17:0]   fft_col_out_payload_50_real,
  output     [17:0]   fft_col_out_payload_50_imag,
  output     [17:0]   fft_col_out_payload_51_real,
  output     [17:0]   fft_col_out_payload_51_imag,
  output     [17:0]   fft_col_out_payload_52_real,
  output     [17:0]   fft_col_out_payload_52_imag,
  output     [17:0]   fft_col_out_payload_53_real,
  output     [17:0]   fft_col_out_payload_53_imag,
  output     [17:0]   fft_col_out_payload_54_real,
  output     [17:0]   fft_col_out_payload_54_imag,
  output     [17:0]   fft_col_out_payload_55_real,
  output     [17:0]   fft_col_out_payload_55_imag,
  output     [17:0]   fft_col_out_payload_56_real,
  output     [17:0]   fft_col_out_payload_56_imag,
  output     [17:0]   fft_col_out_payload_57_real,
  output     [17:0]   fft_col_out_payload_57_imag,
  output     [17:0]   fft_col_out_payload_58_real,
  output     [17:0]   fft_col_out_payload_58_imag,
  output     [17:0]   fft_col_out_payload_59_real,
  output     [17:0]   fft_col_out_payload_59_imag,
  output     [17:0]   fft_col_out_payload_60_real,
  output     [17:0]   fft_col_out_payload_60_imag,
  output     [17:0]   fft_col_out_payload_61_real,
  output     [17:0]   fft_col_out_payload_61_imag,
  output     [17:0]   fft_col_out_payload_62_real,
  output     [17:0]   fft_col_out_payload_62_imag,
  output     [17:0]   fft_col_out_payload_63_real,
  output     [17:0]   fft_col_out_payload_63_imag,
  input               clk,
  input               reset
);
  wire       [35:0]   _zz_961;
  wire       [35:0]   _zz_962;
  wire       [35:0]   _zz_963;
  wire       [35:0]   _zz_964;
  wire       [35:0]   _zz_965;
  wire       [35:0]   _zz_966;
  wire       [35:0]   _zz_967;
  wire       [35:0]   _zz_968;
  wire       [35:0]   _zz_969;
  wire       [35:0]   _zz_970;
  wire       [35:0]   _zz_971;
  wire       [35:0]   _zz_972;
  wire       [35:0]   _zz_973;
  wire       [35:0]   _zz_974;
  wire       [35:0]   _zz_975;
  wire       [35:0]   _zz_976;
  wire       [35:0]   _zz_977;
  wire       [35:0]   _zz_978;
  wire       [35:0]   _zz_979;
  wire       [35:0]   _zz_980;
  wire       [35:0]   _zz_981;
  wire       [35:0]   _zz_982;
  wire       [35:0]   _zz_983;
  wire       [35:0]   _zz_984;
  wire       [35:0]   _zz_985;
  wire       [35:0]   _zz_986;
  wire       [35:0]   _zz_987;
  wire       [35:0]   _zz_988;
  wire       [35:0]   _zz_989;
  wire       [35:0]   _zz_990;
  wire       [35:0]   _zz_991;
  wire       [35:0]   _zz_992;
  wire       [35:0]   _zz_993;
  wire       [35:0]   _zz_994;
  wire       [35:0]   _zz_995;
  wire       [35:0]   _zz_996;
  wire       [35:0]   _zz_997;
  wire       [35:0]   _zz_998;
  wire       [35:0]   _zz_999;
  wire       [35:0]   _zz_1000;
  wire       [35:0]   _zz_1001;
  wire       [35:0]   _zz_1002;
  wire       [35:0]   _zz_1003;
  wire       [35:0]   _zz_1004;
  wire       [35:0]   _zz_1005;
  wire       [35:0]   _zz_1006;
  wire       [35:0]   _zz_1007;
  wire       [35:0]   _zz_1008;
  wire       [35:0]   _zz_1009;
  wire       [35:0]   _zz_1010;
  wire       [35:0]   _zz_1011;
  wire       [35:0]   _zz_1012;
  wire       [35:0]   _zz_1013;
  wire       [35:0]   _zz_1014;
  wire       [35:0]   _zz_1015;
  wire       [35:0]   _zz_1016;
  wire       [35:0]   _zz_1017;
  wire       [35:0]   _zz_1018;
  wire       [35:0]   _zz_1019;
  wire       [35:0]   _zz_1020;
  wire       [35:0]   _zz_1021;
  wire       [35:0]   _zz_1022;
  wire       [35:0]   _zz_1023;
  wire       [35:0]   _zz_1024;
  wire       [35:0]   _zz_1025;
  wire       [35:0]   _zz_1026;
  wire       [35:0]   _zz_1027;
  wire       [35:0]   _zz_1028;
  wire       [35:0]   _zz_1029;
  wire       [35:0]   _zz_1030;
  wire       [35:0]   _zz_1031;
  wire       [35:0]   _zz_1032;
  wire       [35:0]   _zz_1033;
  wire       [35:0]   _zz_1034;
  wire       [35:0]   _zz_1035;
  wire       [35:0]   _zz_1036;
  wire       [35:0]   _zz_1037;
  wire       [35:0]   _zz_1038;
  wire       [35:0]   _zz_1039;
  wire       [35:0]   _zz_1040;
  wire       [35:0]   _zz_1041;
  wire       [35:0]   _zz_1042;
  wire       [35:0]   _zz_1043;
  wire       [35:0]   _zz_1044;
  wire       [35:0]   _zz_1045;
  wire       [35:0]   _zz_1046;
  wire       [35:0]   _zz_1047;
  wire       [35:0]   _zz_1048;
  wire       [35:0]   _zz_1049;
  wire       [35:0]   _zz_1050;
  wire       [35:0]   _zz_1051;
  wire       [35:0]   _zz_1052;
  wire       [35:0]   _zz_1053;
  wire       [35:0]   _zz_1054;
  wire       [35:0]   _zz_1055;
  wire       [35:0]   _zz_1056;
  wire       [35:0]   _zz_1057;
  wire       [35:0]   _zz_1058;
  wire       [35:0]   _zz_1059;
  wire       [35:0]   _zz_1060;
  wire       [35:0]   _zz_1061;
  wire       [35:0]   _zz_1062;
  wire       [35:0]   _zz_1063;
  wire       [35:0]   _zz_1064;
  wire       [35:0]   _zz_1065;
  wire       [35:0]   _zz_1066;
  wire       [35:0]   _zz_1067;
  wire       [35:0]   _zz_1068;
  wire       [35:0]   _zz_1069;
  wire       [35:0]   _zz_1070;
  wire       [35:0]   _zz_1071;
  wire       [35:0]   _zz_1072;
  wire       [35:0]   _zz_1073;
  wire       [35:0]   _zz_1074;
  wire       [35:0]   _zz_1075;
  wire       [35:0]   _zz_1076;
  wire       [35:0]   _zz_1077;
  wire       [35:0]   _zz_1078;
  wire       [35:0]   _zz_1079;
  wire       [35:0]   _zz_1080;
  wire       [35:0]   _zz_1081;
  wire       [35:0]   _zz_1082;
  wire       [35:0]   _zz_1083;
  wire       [35:0]   _zz_1084;
  wire       [35:0]   _zz_1085;
  wire       [35:0]   _zz_1086;
  wire       [35:0]   _zz_1087;
  wire       [35:0]   _zz_1088;
  wire       [35:0]   _zz_1089;
  wire       [35:0]   _zz_1090;
  wire       [35:0]   _zz_1091;
  wire       [35:0]   _zz_1092;
  wire       [35:0]   _zz_1093;
  wire       [35:0]   _zz_1094;
  wire       [35:0]   _zz_1095;
  wire       [35:0]   _zz_1096;
  wire       [35:0]   _zz_1097;
  wire       [35:0]   _zz_1098;
  wire       [35:0]   _zz_1099;
  wire       [35:0]   _zz_1100;
  wire       [35:0]   _zz_1101;
  wire       [35:0]   _zz_1102;
  wire       [35:0]   _zz_1103;
  wire       [35:0]   _zz_1104;
  wire       [35:0]   _zz_1105;
  wire       [35:0]   _zz_1106;
  wire       [35:0]   _zz_1107;
  wire       [35:0]   _zz_1108;
  wire       [35:0]   _zz_1109;
  wire       [35:0]   _zz_1110;
  wire       [35:0]   _zz_1111;
  wire       [35:0]   _zz_1112;
  wire       [35:0]   _zz_1113;
  wire       [35:0]   _zz_1114;
  wire       [35:0]   _zz_1115;
  wire       [35:0]   _zz_1116;
  wire       [35:0]   _zz_1117;
  wire       [35:0]   _zz_1118;
  wire       [35:0]   _zz_1119;
  wire       [35:0]   _zz_1120;
  wire       [35:0]   _zz_1121;
  wire       [35:0]   _zz_1122;
  wire       [35:0]   _zz_1123;
  wire       [35:0]   _zz_1124;
  wire       [35:0]   _zz_1125;
  wire       [35:0]   _zz_1126;
  wire       [35:0]   _zz_1127;
  wire       [35:0]   _zz_1128;
  wire       [35:0]   _zz_1129;
  wire       [35:0]   _zz_1130;
  wire       [35:0]   _zz_1131;
  wire       [35:0]   _zz_1132;
  wire       [35:0]   _zz_1133;
  wire       [35:0]   _zz_1134;
  wire       [35:0]   _zz_1135;
  wire       [35:0]   _zz_1136;
  wire       [35:0]   _zz_1137;
  wire       [35:0]   _zz_1138;
  wire       [35:0]   _zz_1139;
  wire       [35:0]   _zz_1140;
  wire       [35:0]   _zz_1141;
  wire       [35:0]   _zz_1142;
  wire       [35:0]   _zz_1143;
  wire       [35:0]   _zz_1144;
  wire       [35:0]   _zz_1145;
  wire       [35:0]   _zz_1146;
  wire       [35:0]   _zz_1147;
  wire       [35:0]   _zz_1148;
  wire       [35:0]   _zz_1149;
  wire       [35:0]   _zz_1150;
  wire       [35:0]   _zz_1151;
  wire       [35:0]   _zz_1152;
  wire       [35:0]   _zz_1153;
  wire       [35:0]   _zz_1154;
  wire       [35:0]   _zz_1155;
  wire       [35:0]   _zz_1156;
  wire       [35:0]   _zz_1157;
  wire       [35:0]   _zz_1158;
  wire       [35:0]   _zz_1159;
  wire       [35:0]   _zz_1160;
  wire       [35:0]   _zz_1161;
  wire       [35:0]   _zz_1162;
  wire       [35:0]   _zz_1163;
  wire       [35:0]   _zz_1164;
  wire       [35:0]   _zz_1165;
  wire       [35:0]   _zz_1166;
  wire       [35:0]   _zz_1167;
  wire       [35:0]   _zz_1168;
  wire       [35:0]   _zz_1169;
  wire       [35:0]   _zz_1170;
  wire       [35:0]   _zz_1171;
  wire       [35:0]   _zz_1172;
  wire       [35:0]   _zz_1173;
  wire       [35:0]   _zz_1174;
  wire       [35:0]   _zz_1175;
  wire       [35:0]   _zz_1176;
  wire       [35:0]   _zz_1177;
  wire       [35:0]   _zz_1178;
  wire       [35:0]   _zz_1179;
  wire       [35:0]   _zz_1180;
  wire       [35:0]   _zz_1181;
  wire       [35:0]   _zz_1182;
  wire       [35:0]   _zz_1183;
  wire       [35:0]   _zz_1184;
  wire       [35:0]   _zz_1185;
  wire       [35:0]   _zz_1186;
  wire       [35:0]   _zz_1187;
  wire       [35:0]   _zz_1188;
  wire       [35:0]   _zz_1189;
  wire       [35:0]   _zz_1190;
  wire       [35:0]   _zz_1191;
  wire       [35:0]   _zz_1192;
  wire       [35:0]   _zz_1193;
  wire       [35:0]   _zz_1194;
  wire       [35:0]   _zz_1195;
  wire       [35:0]   _zz_1196;
  wire       [35:0]   _zz_1197;
  wire       [35:0]   _zz_1198;
  wire       [35:0]   _zz_1199;
  wire       [35:0]   _zz_1200;
  wire       [35:0]   _zz_1201;
  wire       [35:0]   _zz_1202;
  wire       [35:0]   _zz_1203;
  wire       [35:0]   _zz_1204;
  wire       [35:0]   _zz_1205;
  wire       [35:0]   _zz_1206;
  wire       [35:0]   _zz_1207;
  wire       [35:0]   _zz_1208;
  wire       [35:0]   _zz_1209;
  wire       [35:0]   _zz_1210;
  wire       [35:0]   _zz_1211;
  wire       [35:0]   _zz_1212;
  wire       [35:0]   _zz_1213;
  wire       [35:0]   _zz_1214;
  wire       [35:0]   _zz_1215;
  wire       [35:0]   _zz_1216;
  wire       [35:0]   _zz_1217;
  wire       [35:0]   _zz_1218;
  wire       [35:0]   _zz_1219;
  wire       [35:0]   _zz_1220;
  wire       [35:0]   _zz_1221;
  wire       [35:0]   _zz_1222;
  wire       [35:0]   _zz_1223;
  wire       [35:0]   _zz_1224;
  wire       [35:0]   _zz_1225;
  wire       [35:0]   _zz_1226;
  wire       [35:0]   _zz_1227;
  wire       [35:0]   _zz_1228;
  wire       [35:0]   _zz_1229;
  wire       [35:0]   _zz_1230;
  wire       [35:0]   _zz_1231;
  wire       [35:0]   _zz_1232;
  wire       [35:0]   _zz_1233;
  wire       [35:0]   _zz_1234;
  wire       [35:0]   _zz_1235;
  wire       [35:0]   _zz_1236;
  wire       [35:0]   _zz_1237;
  wire       [35:0]   _zz_1238;
  wire       [35:0]   _zz_1239;
  wire       [35:0]   _zz_1240;
  wire       [35:0]   _zz_1241;
  wire       [35:0]   _zz_1242;
  wire       [35:0]   _zz_1243;
  wire       [35:0]   _zz_1244;
  wire       [35:0]   _zz_1245;
  wire       [35:0]   _zz_1246;
  wire       [35:0]   _zz_1247;
  wire       [35:0]   _zz_1248;
  wire       [35:0]   _zz_1249;
  wire       [35:0]   _zz_1250;
  wire       [35:0]   _zz_1251;
  wire       [35:0]   _zz_1252;
  wire       [35:0]   _zz_1253;
  wire       [35:0]   _zz_1254;
  wire       [35:0]   _zz_1255;
  wire       [35:0]   _zz_1256;
  wire       [35:0]   _zz_1257;
  wire       [35:0]   _zz_1258;
  wire       [35:0]   _zz_1259;
  wire       [35:0]   _zz_1260;
  wire       [35:0]   _zz_1261;
  wire       [35:0]   _zz_1262;
  wire       [35:0]   _zz_1263;
  wire       [35:0]   _zz_1264;
  wire       [35:0]   _zz_1265;
  wire       [35:0]   _zz_1266;
  wire       [35:0]   _zz_1267;
  wire       [35:0]   _zz_1268;
  wire       [35:0]   _zz_1269;
  wire       [35:0]   _zz_1270;
  wire       [35:0]   _zz_1271;
  wire       [35:0]   _zz_1272;
  wire       [35:0]   _zz_1273;
  wire       [35:0]   _zz_1274;
  wire       [35:0]   _zz_1275;
  wire       [35:0]   _zz_1276;
  wire       [35:0]   _zz_1277;
  wire       [35:0]   _zz_1278;
  wire       [35:0]   _zz_1279;
  wire       [35:0]   _zz_1280;
  wire       [35:0]   _zz_1281;
  wire       [35:0]   _zz_1282;
  wire       [35:0]   _zz_1283;
  wire       [35:0]   _zz_1284;
  wire       [35:0]   _zz_1285;
  wire       [35:0]   _zz_1286;
  wire       [35:0]   _zz_1287;
  wire       [35:0]   _zz_1288;
  wire       [35:0]   _zz_1289;
  wire       [35:0]   _zz_1290;
  wire       [35:0]   _zz_1291;
  wire       [35:0]   _zz_1292;
  wire       [35:0]   _zz_1293;
  wire       [35:0]   _zz_1294;
  wire       [35:0]   _zz_1295;
  wire       [35:0]   _zz_1296;
  wire       [35:0]   _zz_1297;
  wire       [35:0]   _zz_1298;
  wire       [35:0]   _zz_1299;
  wire       [35:0]   _zz_1300;
  wire       [35:0]   _zz_1301;
  wire       [35:0]   _zz_1302;
  wire       [35:0]   _zz_1303;
  wire       [35:0]   _zz_1304;
  wire       [35:0]   _zz_1305;
  wire       [35:0]   _zz_1306;
  wire       [35:0]   _zz_1307;
  wire       [35:0]   _zz_1308;
  wire       [35:0]   _zz_1309;
  wire       [35:0]   _zz_1310;
  wire       [35:0]   _zz_1311;
  wire       [35:0]   _zz_1312;
  wire       [35:0]   _zz_1313;
  wire       [35:0]   _zz_1314;
  wire       [35:0]   _zz_1315;
  wire       [35:0]   _zz_1316;
  wire       [35:0]   _zz_1317;
  wire       [35:0]   _zz_1318;
  wire       [35:0]   _zz_1319;
  wire       [35:0]   _zz_1320;
  wire       [35:0]   _zz_1321;
  wire       [35:0]   _zz_1322;
  wire       [35:0]   _zz_1323;
  wire       [35:0]   _zz_1324;
  wire       [35:0]   _zz_1325;
  wire       [35:0]   _zz_1326;
  wire       [35:0]   _zz_1327;
  wire       [35:0]   _zz_1328;
  wire       [35:0]   _zz_1329;
  wire       [35:0]   _zz_1330;
  wire       [35:0]   _zz_1331;
  wire       [35:0]   _zz_1332;
  wire       [35:0]   _zz_1333;
  wire       [35:0]   _zz_1334;
  wire       [35:0]   _zz_1335;
  wire       [35:0]   _zz_1336;
  wire       [35:0]   _zz_1337;
  wire       [35:0]   _zz_1338;
  wire       [35:0]   _zz_1339;
  wire       [35:0]   _zz_1340;
  wire       [35:0]   _zz_1341;
  wire       [35:0]   _zz_1342;
  wire       [35:0]   _zz_1343;
  wire       [35:0]   _zz_1344;
  wire       [35:0]   _zz_1345;
  wire       [35:0]   _zz_1346;
  wire       [35:0]   _zz_1347;
  wire       [35:0]   _zz_1348;
  wire       [35:0]   _zz_1349;
  wire       [35:0]   _zz_1350;
  wire       [35:0]   _zz_1351;
  wire       [35:0]   _zz_1352;
  wire       [35:0]   _zz_1353;
  wire       [35:0]   _zz_1354;
  wire       [35:0]   _zz_1355;
  wire       [35:0]   _zz_1356;
  wire       [35:0]   _zz_1357;
  wire       [35:0]   _zz_1358;
  wire       [35:0]   _zz_1359;
  wire       [35:0]   _zz_1360;
  wire       [35:0]   _zz_1361;
  wire       [35:0]   _zz_1362;
  wire       [35:0]   _zz_1363;
  wire       [35:0]   _zz_1364;
  wire       [35:0]   _zz_1365;
  wire       [35:0]   _zz_1366;
  wire       [35:0]   _zz_1367;
  wire       [35:0]   _zz_1368;
  wire       [35:0]   _zz_1369;
  wire       [35:0]   _zz_1370;
  wire       [35:0]   _zz_1371;
  wire       [35:0]   _zz_1372;
  wire       [35:0]   _zz_1373;
  wire       [35:0]   _zz_1374;
  wire       [35:0]   _zz_1375;
  wire       [35:0]   _zz_1376;
  wire       [35:0]   _zz_1377;
  wire       [35:0]   _zz_1378;
  wire       [35:0]   _zz_1379;
  wire       [35:0]   _zz_1380;
  wire       [35:0]   _zz_1381;
  wire       [35:0]   _zz_1382;
  wire       [35:0]   _zz_1383;
  wire       [35:0]   _zz_1384;
  wire       [35:0]   _zz_1385;
  wire       [35:0]   _zz_1386;
  wire       [35:0]   _zz_1387;
  wire       [35:0]   _zz_1388;
  wire       [35:0]   _zz_1389;
  wire       [35:0]   _zz_1390;
  wire       [35:0]   _zz_1391;
  wire       [35:0]   _zz_1392;
  wire       [35:0]   _zz_1393;
  wire       [35:0]   _zz_1394;
  wire       [35:0]   _zz_1395;
  wire       [35:0]   _zz_1396;
  wire       [35:0]   _zz_1397;
  wire       [35:0]   _zz_1398;
  wire       [35:0]   _zz_1399;
  wire       [35:0]   _zz_1400;
  wire       [35:0]   _zz_1401;
  wire       [35:0]   _zz_1402;
  wire       [35:0]   _zz_1403;
  wire       [35:0]   _zz_1404;
  wire       [35:0]   _zz_1405;
  wire       [35:0]   _zz_1406;
  wire       [35:0]   _zz_1407;
  wire       [35:0]   _zz_1408;
  wire       [35:0]   _zz_1409;
  wire       [35:0]   _zz_1410;
  wire       [35:0]   _zz_1411;
  wire       [35:0]   _zz_1412;
  wire       [35:0]   _zz_1413;
  wire       [35:0]   _zz_1414;
  wire       [35:0]   _zz_1415;
  wire       [35:0]   _zz_1416;
  wire       [35:0]   _zz_1417;
  wire       [35:0]   _zz_1418;
  wire       [35:0]   _zz_1419;
  wire       [35:0]   _zz_1420;
  wire       [35:0]   _zz_1421;
  wire       [35:0]   _zz_1422;
  wire       [35:0]   _zz_1423;
  wire       [35:0]   _zz_1424;
  wire       [35:0]   _zz_1425;
  wire       [35:0]   _zz_1426;
  wire       [35:0]   _zz_1427;
  wire       [35:0]   _zz_1428;
  wire       [35:0]   _zz_1429;
  wire       [35:0]   _zz_1430;
  wire       [35:0]   _zz_1431;
  wire       [35:0]   _zz_1432;
  wire       [35:0]   _zz_1433;
  wire       [35:0]   _zz_1434;
  wire       [35:0]   _zz_1435;
  wire       [35:0]   _zz_1436;
  wire       [35:0]   _zz_1437;
  wire       [35:0]   _zz_1438;
  wire       [35:0]   _zz_1439;
  wire       [35:0]   _zz_1440;
  wire       [35:0]   _zz_1441;
  wire       [35:0]   _zz_1442;
  wire       [35:0]   _zz_1443;
  wire       [35:0]   _zz_1444;
  wire       [35:0]   _zz_1445;
  wire       [35:0]   _zz_1446;
  wire       [35:0]   _zz_1447;
  wire       [35:0]   _zz_1448;
  wire       [35:0]   _zz_1449;
  wire       [35:0]   _zz_1450;
  wire       [35:0]   _zz_1451;
  wire       [35:0]   _zz_1452;
  wire       [35:0]   _zz_1453;
  wire       [35:0]   _zz_1454;
  wire       [35:0]   _zz_1455;
  wire       [35:0]   _zz_1456;
  wire       [35:0]   _zz_1457;
  wire       [35:0]   _zz_1458;
  wire       [35:0]   _zz_1459;
  wire       [35:0]   _zz_1460;
  wire       [35:0]   _zz_1461;
  wire       [35:0]   _zz_1462;
  wire       [35:0]   _zz_1463;
  wire       [35:0]   _zz_1464;
  wire       [35:0]   _zz_1465;
  wire       [35:0]   _zz_1466;
  wire       [35:0]   _zz_1467;
  wire       [35:0]   _zz_1468;
  wire       [35:0]   _zz_1469;
  wire       [35:0]   _zz_1470;
  wire       [35:0]   _zz_1471;
  wire       [35:0]   _zz_1472;
  wire       [35:0]   _zz_1473;
  wire       [35:0]   _zz_1474;
  wire       [35:0]   _zz_1475;
  wire       [35:0]   _zz_1476;
  wire       [35:0]   _zz_1477;
  wire       [35:0]   _zz_1478;
  wire       [35:0]   _zz_1479;
  wire       [35:0]   _zz_1480;
  wire       [35:0]   _zz_1481;
  wire       [35:0]   _zz_1482;
  wire       [35:0]   _zz_1483;
  wire       [35:0]   _zz_1484;
  wire       [35:0]   _zz_1485;
  wire       [35:0]   _zz_1486;
  wire       [35:0]   _zz_1487;
  wire       [35:0]   _zz_1488;
  wire       [35:0]   _zz_1489;
  wire       [35:0]   _zz_1490;
  wire       [35:0]   _zz_1491;
  wire       [35:0]   _zz_1492;
  wire       [35:0]   _zz_1493;
  wire       [35:0]   _zz_1494;
  wire       [35:0]   _zz_1495;
  wire       [35:0]   _zz_1496;
  wire       [35:0]   _zz_1497;
  wire       [35:0]   _zz_1498;
  wire       [35:0]   _zz_1499;
  wire       [35:0]   _zz_1500;
  wire       [35:0]   _zz_1501;
  wire       [35:0]   _zz_1502;
  wire       [35:0]   _zz_1503;
  wire       [35:0]   _zz_1504;
  wire       [35:0]   _zz_1505;
  wire       [35:0]   _zz_1506;
  wire       [35:0]   _zz_1507;
  wire       [35:0]   _zz_1508;
  wire       [35:0]   _zz_1509;
  wire       [35:0]   _zz_1510;
  wire       [35:0]   _zz_1511;
  wire       [35:0]   _zz_1512;
  wire       [35:0]   _zz_1513;
  wire       [35:0]   _zz_1514;
  wire       [35:0]   _zz_1515;
  wire       [35:0]   _zz_1516;
  wire       [35:0]   _zz_1517;
  wire       [35:0]   _zz_1518;
  wire       [35:0]   _zz_1519;
  wire       [35:0]   _zz_1520;
  wire       [35:0]   _zz_1521;
  wire       [35:0]   _zz_1522;
  wire       [35:0]   _zz_1523;
  wire       [35:0]   _zz_1524;
  wire       [35:0]   _zz_1525;
  wire       [35:0]   _zz_1526;
  wire       [35:0]   _zz_1527;
  wire       [35:0]   _zz_1528;
  wire       [35:0]   _zz_1529;
  wire       [35:0]   _zz_1530;
  wire       [35:0]   _zz_1531;
  wire       [35:0]   _zz_1532;
  wire       [35:0]   _zz_1533;
  wire       [35:0]   _zz_1534;
  wire       [35:0]   _zz_1535;
  wire       [35:0]   _zz_1536;
  wire       [35:0]   _zz_1537;
  wire       [35:0]   _zz_1538;
  wire       [35:0]   _zz_1539;
  wire       [35:0]   _zz_1540;
  wire       [35:0]   _zz_1541;
  wire       [35:0]   _zz_1542;
  wire       [35:0]   _zz_1543;
  wire       [35:0]   _zz_1544;
  wire       [35:0]   _zz_1545;
  wire       [35:0]   _zz_1546;
  wire       [35:0]   _zz_1547;
  wire       [35:0]   _zz_1548;
  wire       [35:0]   _zz_1549;
  wire       [35:0]   _zz_1550;
  wire       [35:0]   _zz_1551;
  wire       [35:0]   _zz_1552;
  wire       [35:0]   _zz_1553;
  wire       [35:0]   _zz_1554;
  wire       [35:0]   _zz_1555;
  wire       [35:0]   _zz_1556;
  wire       [35:0]   _zz_1557;
  wire       [35:0]   _zz_1558;
  wire       [35:0]   _zz_1559;
  wire       [35:0]   _zz_1560;
  wire       [35:0]   _zz_1561;
  wire       [35:0]   _zz_1562;
  wire       [35:0]   _zz_1563;
  wire       [35:0]   _zz_1564;
  wire       [35:0]   _zz_1565;
  wire       [35:0]   _zz_1566;
  wire       [35:0]   _zz_1567;
  wire       [35:0]   _zz_1568;
  wire       [35:0]   _zz_1569;
  wire       [35:0]   _zz_1570;
  wire       [35:0]   _zz_1571;
  wire       [35:0]   _zz_1572;
  wire       [35:0]   _zz_1573;
  wire       [35:0]   _zz_1574;
  wire       [35:0]   _zz_1575;
  wire       [35:0]   _zz_1576;
  wire       [35:0]   _zz_1577;
  wire       [35:0]   _zz_1578;
  wire       [35:0]   _zz_1579;
  wire       [35:0]   _zz_1580;
  wire       [35:0]   _zz_1581;
  wire       [35:0]   _zz_1582;
  wire       [35:0]   _zz_1583;
  wire       [35:0]   _zz_1584;
  wire       [35:0]   _zz_1585;
  wire       [35:0]   _zz_1586;
  wire       [35:0]   _zz_1587;
  wire       [35:0]   _zz_1588;
  wire       [35:0]   _zz_1589;
  wire       [35:0]   _zz_1590;
  wire       [35:0]   _zz_1591;
  wire       [35:0]   _zz_1592;
  wire       [35:0]   _zz_1593;
  wire       [35:0]   _zz_1594;
  wire       [35:0]   _zz_1595;
  wire       [35:0]   _zz_1596;
  wire       [35:0]   _zz_1597;
  wire       [35:0]   _zz_1598;
  wire       [35:0]   _zz_1599;
  wire       [35:0]   _zz_1600;
  wire       [35:0]   _zz_1601;
  wire       [35:0]   _zz_1602;
  wire       [35:0]   _zz_1603;
  wire       [35:0]   _zz_1604;
  wire       [35:0]   _zz_1605;
  wire       [35:0]   _zz_1606;
  wire       [35:0]   _zz_1607;
  wire       [35:0]   _zz_1608;
  wire       [35:0]   _zz_1609;
  wire       [35:0]   _zz_1610;
  wire       [35:0]   _zz_1611;
  wire       [35:0]   _zz_1612;
  wire       [35:0]   _zz_1613;
  wire       [35:0]   _zz_1614;
  wire       [35:0]   _zz_1615;
  wire       [35:0]   _zz_1616;
  wire       [35:0]   _zz_1617;
  wire       [35:0]   _zz_1618;
  wire       [35:0]   _zz_1619;
  wire       [35:0]   _zz_1620;
  wire       [35:0]   _zz_1621;
  wire       [35:0]   _zz_1622;
  wire       [35:0]   _zz_1623;
  wire       [35:0]   _zz_1624;
  wire       [35:0]   _zz_1625;
  wire       [35:0]   _zz_1626;
  wire       [35:0]   _zz_1627;
  wire       [35:0]   _zz_1628;
  wire       [35:0]   _zz_1629;
  wire       [35:0]   _zz_1630;
  wire       [35:0]   _zz_1631;
  wire       [35:0]   _zz_1632;
  wire       [35:0]   _zz_1633;
  wire       [35:0]   _zz_1634;
  wire       [35:0]   _zz_1635;
  wire       [35:0]   _zz_1636;
  wire       [35:0]   _zz_1637;
  wire       [35:0]   _zz_1638;
  wire       [35:0]   _zz_1639;
  wire       [35:0]   _zz_1640;
  wire       [35:0]   _zz_1641;
  wire       [35:0]   _zz_1642;
  wire       [35:0]   _zz_1643;
  wire       [35:0]   _zz_1644;
  wire       [35:0]   _zz_1645;
  wire       [35:0]   _zz_1646;
  wire       [35:0]   _zz_1647;
  wire       [35:0]   _zz_1648;
  wire       [35:0]   _zz_1649;
  wire       [35:0]   _zz_1650;
  wire       [35:0]   _zz_1651;
  wire       [35:0]   _zz_1652;
  wire       [35:0]   _zz_1653;
  wire       [35:0]   _zz_1654;
  wire       [35:0]   _zz_1655;
  wire       [35:0]   _zz_1656;
  wire       [35:0]   _zz_1657;
  wire       [35:0]   _zz_1658;
  wire       [35:0]   _zz_1659;
  wire       [35:0]   _zz_1660;
  wire       [35:0]   _zz_1661;
  wire       [35:0]   _zz_1662;
  wire       [35:0]   _zz_1663;
  wire       [35:0]   _zz_1664;
  wire       [35:0]   _zz_1665;
  wire       [35:0]   _zz_1666;
  wire       [35:0]   _zz_1667;
  wire       [35:0]   _zz_1668;
  wire       [35:0]   _zz_1669;
  wire       [35:0]   _zz_1670;
  wire       [35:0]   _zz_1671;
  wire       [35:0]   _zz_1672;
  wire       [35:0]   _zz_1673;
  wire       [35:0]   _zz_1674;
  wire       [35:0]   _zz_1675;
  wire       [35:0]   _zz_1676;
  wire       [35:0]   _zz_1677;
  wire       [35:0]   _zz_1678;
  wire       [35:0]   _zz_1679;
  wire       [35:0]   _zz_1680;
  wire       [35:0]   _zz_1681;
  wire       [35:0]   _zz_1682;
  wire       [35:0]   _zz_1683;
  wire       [35:0]   _zz_1684;
  wire       [35:0]   _zz_1685;
  wire       [35:0]   _zz_1686;
  wire       [35:0]   _zz_1687;
  wire       [35:0]   _zz_1688;
  wire       [35:0]   _zz_1689;
  wire       [35:0]   _zz_1690;
  wire       [35:0]   _zz_1691;
  wire       [35:0]   _zz_1692;
  wire       [35:0]   _zz_1693;
  wire       [35:0]   _zz_1694;
  wire       [35:0]   _zz_1695;
  wire       [35:0]   _zz_1696;
  wire       [35:0]   _zz_1697;
  wire       [35:0]   _zz_1698;
  wire       [35:0]   _zz_1699;
  wire       [35:0]   _zz_1700;
  wire       [35:0]   _zz_1701;
  wire       [35:0]   _zz_1702;
  wire       [35:0]   _zz_1703;
  wire       [35:0]   _zz_1704;
  wire       [35:0]   _zz_1705;
  wire       [35:0]   _zz_1706;
  wire       [35:0]   _zz_1707;
  wire       [35:0]   _zz_1708;
  wire       [35:0]   _zz_1709;
  wire       [35:0]   _zz_1710;
  wire       [35:0]   _zz_1711;
  wire       [35:0]   _zz_1712;
  wire       [35:0]   _zz_1713;
  wire       [35:0]   _zz_1714;
  wire       [35:0]   _zz_1715;
  wire       [35:0]   _zz_1716;
  wire       [35:0]   _zz_1717;
  wire       [35:0]   _zz_1718;
  wire       [35:0]   _zz_1719;
  wire       [35:0]   _zz_1720;
  wire       [35:0]   _zz_1721;
  wire       [35:0]   _zz_1722;
  wire       [35:0]   _zz_1723;
  wire       [35:0]   _zz_1724;
  wire       [35:0]   _zz_1725;
  wire       [35:0]   _zz_1726;
  wire       [35:0]   _zz_1727;
  wire       [35:0]   _zz_1728;
  wire       [35:0]   _zz_1729;
  wire       [35:0]   _zz_1730;
  wire       [35:0]   _zz_1731;
  wire       [35:0]   _zz_1732;
  wire       [35:0]   _zz_1733;
  wire       [35:0]   _zz_1734;
  wire       [35:0]   _zz_1735;
  wire       [35:0]   _zz_1736;
  wire       [35:0]   _zz_1737;
  wire       [35:0]   _zz_1738;
  wire       [35:0]   _zz_1739;
  wire       [35:0]   _zz_1740;
  wire       [35:0]   _zz_1741;
  wire       [35:0]   _zz_1742;
  wire       [35:0]   _zz_1743;
  wire       [35:0]   _zz_1744;
  wire       [35:0]   _zz_1745;
  wire       [35:0]   _zz_1746;
  wire       [35:0]   _zz_1747;
  wire       [35:0]   _zz_1748;
  wire       [35:0]   _zz_1749;
  wire       [35:0]   _zz_1750;
  wire       [35:0]   _zz_1751;
  wire       [35:0]   _zz_1752;
  wire       [35:0]   _zz_1753;
  wire       [35:0]   _zz_1754;
  wire       [35:0]   _zz_1755;
  wire       [35:0]   _zz_1756;
  wire       [35:0]   _zz_1757;
  wire       [35:0]   _zz_1758;
  wire       [35:0]   _zz_1759;
  wire       [35:0]   _zz_1760;
  wire       [35:0]   _zz_1761;
  wire       [35:0]   _zz_1762;
  wire       [35:0]   _zz_1763;
  wire       [35:0]   _zz_1764;
  wire       [35:0]   _zz_1765;
  wire       [35:0]   _zz_1766;
  wire       [35:0]   _zz_1767;
  wire       [35:0]   _zz_1768;
  wire       [35:0]   _zz_1769;
  wire       [35:0]   _zz_1770;
  wire       [35:0]   _zz_1771;
  wire       [35:0]   _zz_1772;
  wire       [35:0]   _zz_1773;
  wire       [35:0]   _zz_1774;
  wire       [35:0]   _zz_1775;
  wire       [35:0]   _zz_1776;
  wire       [35:0]   _zz_1777;
  wire       [35:0]   _zz_1778;
  wire       [35:0]   _zz_1779;
  wire       [35:0]   _zz_1780;
  wire       [35:0]   _zz_1781;
  wire       [35:0]   _zz_1782;
  wire       [35:0]   _zz_1783;
  wire       [35:0]   _zz_1784;
  wire       [35:0]   _zz_1785;
  wire       [35:0]   _zz_1786;
  wire       [35:0]   _zz_1787;
  wire       [35:0]   _zz_1788;
  wire       [35:0]   _zz_1789;
  wire       [35:0]   _zz_1790;
  wire       [35:0]   _zz_1791;
  wire       [35:0]   _zz_1792;
  wire       [35:0]   _zz_1793;
  wire       [35:0]   _zz_1794;
  wire       [35:0]   _zz_1795;
  wire       [35:0]   _zz_1796;
  wire       [35:0]   _zz_1797;
  wire       [35:0]   _zz_1798;
  wire       [35:0]   _zz_1799;
  wire       [35:0]   _zz_1800;
  wire       [35:0]   _zz_1801;
  wire       [35:0]   _zz_1802;
  wire       [35:0]   _zz_1803;
  wire       [35:0]   _zz_1804;
  wire       [35:0]   _zz_1805;
  wire       [35:0]   _zz_1806;
  wire       [35:0]   _zz_1807;
  wire       [35:0]   _zz_1808;
  wire       [35:0]   _zz_1809;
  wire       [35:0]   _zz_1810;
  wire       [35:0]   _zz_1811;
  wire       [35:0]   _zz_1812;
  wire       [35:0]   _zz_1813;
  wire       [35:0]   _zz_1814;
  wire       [35:0]   _zz_1815;
  wire       [35:0]   _zz_1816;
  wire       [35:0]   _zz_1817;
  wire       [35:0]   _zz_1818;
  wire       [35:0]   _zz_1819;
  wire       [35:0]   _zz_1820;
  wire       [35:0]   _zz_1821;
  wire       [35:0]   _zz_1822;
  wire       [35:0]   _zz_1823;
  wire       [35:0]   _zz_1824;
  wire       [35:0]   _zz_1825;
  wire       [35:0]   _zz_1826;
  wire       [35:0]   _zz_1827;
  wire       [35:0]   _zz_1828;
  wire       [35:0]   _zz_1829;
  wire       [35:0]   _zz_1830;
  wire       [35:0]   _zz_1831;
  wire       [35:0]   _zz_1832;
  wire       [35:0]   _zz_1833;
  wire       [35:0]   _zz_1834;
  wire       [35:0]   _zz_1835;
  wire       [35:0]   _zz_1836;
  wire       [35:0]   _zz_1837;
  wire       [35:0]   _zz_1838;
  wire       [35:0]   _zz_1839;
  wire       [35:0]   _zz_1840;
  wire       [35:0]   _zz_1841;
  wire       [35:0]   _zz_1842;
  wire       [35:0]   _zz_1843;
  wire       [35:0]   _zz_1844;
  wire       [35:0]   _zz_1845;
  wire       [35:0]   _zz_1846;
  wire       [35:0]   _zz_1847;
  wire       [35:0]   _zz_1848;
  wire       [35:0]   _zz_1849;
  wire       [35:0]   _zz_1850;
  wire       [35:0]   _zz_1851;
  wire       [35:0]   _zz_1852;
  wire       [35:0]   _zz_1853;
  wire       [35:0]   _zz_1854;
  wire       [35:0]   _zz_1855;
  wire       [35:0]   _zz_1856;
  wire       [35:0]   _zz_1857;
  wire       [35:0]   _zz_1858;
  wire       [35:0]   _zz_1859;
  wire       [35:0]   _zz_1860;
  wire       [35:0]   _zz_1861;
  wire       [35:0]   _zz_1862;
  wire       [35:0]   _zz_1863;
  wire       [35:0]   _zz_1864;
  wire       [35:0]   _zz_1865;
  wire       [35:0]   _zz_1866;
  wire       [35:0]   _zz_1867;
  wire       [35:0]   _zz_1868;
  wire       [35:0]   _zz_1869;
  wire       [35:0]   _zz_1870;
  wire       [35:0]   _zz_1871;
  wire       [35:0]   _zz_1872;
  wire       [35:0]   _zz_1873;
  wire       [35:0]   _zz_1874;
  wire       [35:0]   _zz_1875;
  wire       [35:0]   _zz_1876;
  wire       [35:0]   _zz_1877;
  wire       [35:0]   _zz_1878;
  wire       [35:0]   _zz_1879;
  wire       [35:0]   _zz_1880;
  wire       [35:0]   _zz_1881;
  wire       [35:0]   _zz_1882;
  wire       [35:0]   _zz_1883;
  wire       [35:0]   _zz_1884;
  wire       [35:0]   _zz_1885;
  wire       [35:0]   _zz_1886;
  wire       [35:0]   _zz_1887;
  wire       [35:0]   _zz_1888;
  wire       [35:0]   _zz_1889;
  wire       [35:0]   _zz_1890;
  wire       [35:0]   _zz_1891;
  wire       [35:0]   _zz_1892;
  wire       [35:0]   _zz_1893;
  wire       [35:0]   _zz_1894;
  wire       [35:0]   _zz_1895;
  wire       [35:0]   _zz_1896;
  wire       [35:0]   _zz_1897;
  wire       [35:0]   _zz_1898;
  wire       [35:0]   _zz_1899;
  wire       [35:0]   _zz_1900;
  wire       [35:0]   _zz_1901;
  wire       [35:0]   _zz_1902;
  wire       [35:0]   _zz_1903;
  wire       [35:0]   _zz_1904;
  wire       [35:0]   _zz_1905;
  wire       [35:0]   _zz_1906;
  wire       [35:0]   _zz_1907;
  wire       [35:0]   _zz_1908;
  wire       [35:0]   _zz_1909;
  wire       [35:0]   _zz_1910;
  wire       [35:0]   _zz_1911;
  wire       [35:0]   _zz_1912;
  wire       [35:0]   _zz_1913;
  wire       [35:0]   _zz_1914;
  wire       [35:0]   _zz_1915;
  wire       [35:0]   _zz_1916;
  wire       [35:0]   _zz_1917;
  wire       [35:0]   _zz_1918;
  wire       [35:0]   _zz_1919;
  wire       [35:0]   _zz_1920;
  wire       [35:0]   _zz_1921;
  wire       [35:0]   _zz_1922;
  wire       [35:0]   _zz_1923;
  wire       [35:0]   _zz_1924;
  wire       [35:0]   _zz_1925;
  wire       [35:0]   _zz_1926;
  wire       [35:0]   _zz_1927;
  wire       [35:0]   _zz_1928;
  wire       [35:0]   _zz_1929;
  wire       [35:0]   _zz_1930;
  wire       [35:0]   _zz_1931;
  wire       [35:0]   _zz_1932;
  wire       [35:0]   _zz_1933;
  wire       [35:0]   _zz_1934;
  wire       [35:0]   _zz_1935;
  wire       [35:0]   _zz_1936;
  wire       [35:0]   _zz_1937;
  wire       [35:0]   _zz_1938;
  wire       [35:0]   _zz_1939;
  wire       [35:0]   _zz_1940;
  wire       [35:0]   _zz_1941;
  wire       [35:0]   _zz_1942;
  wire       [35:0]   _zz_1943;
  wire       [35:0]   _zz_1944;
  wire       [35:0]   _zz_1945;
  wire       [35:0]   _zz_1946;
  wire       [35:0]   _zz_1947;
  wire       [35:0]   _zz_1948;
  wire       [35:0]   _zz_1949;
  wire       [35:0]   _zz_1950;
  wire       [35:0]   _zz_1951;
  wire       [35:0]   _zz_1952;
  wire       [35:0]   _zz_1953;
  wire       [35:0]   _zz_1954;
  wire       [35:0]   _zz_1955;
  wire       [35:0]   _zz_1956;
  wire       [35:0]   _zz_1957;
  wire       [35:0]   _zz_1958;
  wire       [35:0]   _zz_1959;
  wire       [35:0]   _zz_1960;
  wire       [35:0]   _zz_1961;
  wire       [35:0]   _zz_1962;
  wire       [35:0]   _zz_1963;
  wire       [35:0]   _zz_1964;
  wire       [35:0]   _zz_1965;
  wire       [35:0]   _zz_1966;
  wire       [35:0]   _zz_1967;
  wire       [35:0]   _zz_1968;
  wire       [35:0]   _zz_1969;
  wire       [35:0]   _zz_1970;
  wire       [35:0]   _zz_1971;
  wire       [35:0]   _zz_1972;
  wire       [35:0]   _zz_1973;
  wire       [35:0]   _zz_1974;
  wire       [35:0]   _zz_1975;
  wire       [35:0]   _zz_1976;
  wire       [35:0]   _zz_1977;
  wire       [35:0]   _zz_1978;
  wire       [35:0]   _zz_1979;
  wire       [35:0]   _zz_1980;
  wire       [35:0]   _zz_1981;
  wire       [35:0]   _zz_1982;
  wire       [35:0]   _zz_1983;
  wire       [35:0]   _zz_1984;
  wire       [35:0]   _zz_1985;
  wire       [35:0]   _zz_1986;
  wire       [35:0]   _zz_1987;
  wire       [35:0]   _zz_1988;
  wire       [35:0]   _zz_1989;
  wire       [35:0]   _zz_1990;
  wire       [35:0]   _zz_1991;
  wire       [35:0]   _zz_1992;
  wire       [35:0]   _zz_1993;
  wire       [35:0]   _zz_1994;
  wire       [35:0]   _zz_1995;
  wire       [35:0]   _zz_1996;
  wire       [35:0]   _zz_1997;
  wire       [35:0]   _zz_1998;
  wire       [35:0]   _zz_1999;
  wire       [35:0]   _zz_2000;
  wire       [35:0]   _zz_2001;
  wire       [35:0]   _zz_2002;
  wire       [35:0]   _zz_2003;
  wire       [35:0]   _zz_2004;
  wire       [35:0]   _zz_2005;
  wire       [35:0]   _zz_2006;
  wire       [35:0]   _zz_2007;
  wire       [35:0]   _zz_2008;
  wire       [35:0]   _zz_2009;
  wire       [35:0]   _zz_2010;
  wire       [35:0]   _zz_2011;
  wire       [35:0]   _zz_2012;
  wire       [35:0]   _zz_2013;
  wire       [35:0]   _zz_2014;
  wire       [35:0]   _zz_2015;
  wire       [35:0]   _zz_2016;
  wire       [35:0]   _zz_2017;
  wire       [35:0]   _zz_2018;
  wire       [35:0]   _zz_2019;
  wire       [35:0]   _zz_2020;
  wire       [35:0]   _zz_2021;
  wire       [35:0]   _zz_2022;
  wire       [35:0]   _zz_2023;
  wire       [35:0]   _zz_2024;
  wire       [35:0]   _zz_2025;
  wire       [35:0]   _zz_2026;
  wire       [35:0]   _zz_2027;
  wire       [35:0]   _zz_2028;
  wire       [35:0]   _zz_2029;
  wire       [35:0]   _zz_2030;
  wire       [35:0]   _zz_2031;
  wire       [35:0]   _zz_2032;
  wire       [35:0]   _zz_2033;
  wire       [35:0]   _zz_2034;
  wire       [35:0]   _zz_2035;
  wire       [35:0]   _zz_2036;
  wire       [35:0]   _zz_2037;
  wire       [35:0]   _zz_2038;
  wire       [35:0]   _zz_2039;
  wire       [35:0]   _zz_2040;
  wire       [35:0]   _zz_2041;
  wire       [35:0]   _zz_2042;
  wire       [35:0]   _zz_2043;
  wire       [35:0]   _zz_2044;
  wire       [35:0]   _zz_2045;
  wire       [35:0]   _zz_2046;
  wire       [35:0]   _zz_2047;
  wire       [35:0]   _zz_2048;
  wire       [35:0]   _zz_2049;
  wire       [35:0]   _zz_2050;
  wire       [35:0]   _zz_2051;
  wire       [35:0]   _zz_2052;
  wire       [35:0]   _zz_2053;
  wire       [35:0]   _zz_2054;
  wire       [35:0]   _zz_2055;
  wire       [35:0]   _zz_2056;
  wire       [35:0]   _zz_2057;
  wire       [35:0]   _zz_2058;
  wire       [35:0]   _zz_2059;
  wire       [35:0]   _zz_2060;
  wire       [35:0]   _zz_2061;
  wire       [35:0]   _zz_2062;
  wire       [35:0]   _zz_2063;
  wire       [35:0]   _zz_2064;
  wire       [35:0]   _zz_2065;
  wire       [35:0]   _zz_2066;
  wire       [35:0]   _zz_2067;
  wire       [35:0]   _zz_2068;
  wire       [35:0]   _zz_2069;
  wire       [35:0]   _zz_2070;
  wire       [35:0]   _zz_2071;
  wire       [35:0]   _zz_2072;
  wire       [35:0]   _zz_2073;
  wire       [35:0]   _zz_2074;
  wire       [35:0]   _zz_2075;
  wire       [35:0]   _zz_2076;
  wire       [35:0]   _zz_2077;
  wire       [35:0]   _zz_2078;
  wire       [35:0]   _zz_2079;
  wire       [35:0]   _zz_2080;
  wire       [35:0]   _zz_2081;
  wire       [35:0]   _zz_2082;
  wire       [35:0]   _zz_2083;
  wire       [35:0]   _zz_2084;
  wire       [35:0]   _zz_2085;
  wire       [35:0]   _zz_2086;
  wire       [35:0]   _zz_2087;
  wire       [35:0]   _zz_2088;
  wire       [35:0]   _zz_2089;
  wire       [35:0]   _zz_2090;
  wire       [35:0]   _zz_2091;
  wire       [35:0]   _zz_2092;
  wire       [35:0]   _zz_2093;
  wire       [35:0]   _zz_2094;
  wire       [35:0]   _zz_2095;
  wire       [35:0]   _zz_2096;
  wire       [35:0]   _zz_2097;
  wire       [35:0]   _zz_2098;
  wire       [35:0]   _zz_2099;
  wire       [35:0]   _zz_2100;
  wire       [35:0]   _zz_2101;
  wire       [35:0]   _zz_2102;
  wire       [35:0]   _zz_2103;
  wire       [35:0]   _zz_2104;
  wire       [35:0]   _zz_2105;
  wire       [35:0]   _zz_2106;
  wire       [35:0]   _zz_2107;
  wire       [35:0]   _zz_2108;
  wire       [35:0]   _zz_2109;
  wire       [35:0]   _zz_2110;
  wire       [35:0]   _zz_2111;
  wire       [35:0]   _zz_2112;
  wire       [35:0]   fixTo_dout;
  wire       [35:0]   fixTo_1_dout;
  wire       [17:0]   fixTo_2_dout;
  wire       [17:0]   fixTo_3_dout;
  wire       [17:0]   fixTo_4_dout;
  wire       [17:0]   fixTo_5_dout;
  wire       [35:0]   fixTo_6_dout;
  wire       [35:0]   fixTo_7_dout;
  wire       [17:0]   fixTo_8_dout;
  wire       [17:0]   fixTo_9_dout;
  wire       [17:0]   fixTo_10_dout;
  wire       [17:0]   fixTo_11_dout;
  wire       [35:0]   fixTo_12_dout;
  wire       [35:0]   fixTo_13_dout;
  wire       [17:0]   fixTo_14_dout;
  wire       [17:0]   fixTo_15_dout;
  wire       [17:0]   fixTo_16_dout;
  wire       [17:0]   fixTo_17_dout;
  wire       [35:0]   fixTo_18_dout;
  wire       [35:0]   fixTo_19_dout;
  wire       [17:0]   fixTo_20_dout;
  wire       [17:0]   fixTo_21_dout;
  wire       [17:0]   fixTo_22_dout;
  wire       [17:0]   fixTo_23_dout;
  wire       [35:0]   fixTo_24_dout;
  wire       [35:0]   fixTo_25_dout;
  wire       [17:0]   fixTo_26_dout;
  wire       [17:0]   fixTo_27_dout;
  wire       [17:0]   fixTo_28_dout;
  wire       [17:0]   fixTo_29_dout;
  wire       [35:0]   fixTo_30_dout;
  wire       [35:0]   fixTo_31_dout;
  wire       [17:0]   fixTo_32_dout;
  wire       [17:0]   fixTo_33_dout;
  wire       [17:0]   fixTo_34_dout;
  wire       [17:0]   fixTo_35_dout;
  wire       [35:0]   fixTo_36_dout;
  wire       [35:0]   fixTo_37_dout;
  wire       [17:0]   fixTo_38_dout;
  wire       [17:0]   fixTo_39_dout;
  wire       [17:0]   fixTo_40_dout;
  wire       [17:0]   fixTo_41_dout;
  wire       [35:0]   fixTo_42_dout;
  wire       [35:0]   fixTo_43_dout;
  wire       [17:0]   fixTo_44_dout;
  wire       [17:0]   fixTo_45_dout;
  wire       [17:0]   fixTo_46_dout;
  wire       [17:0]   fixTo_47_dout;
  wire       [35:0]   fixTo_48_dout;
  wire       [35:0]   fixTo_49_dout;
  wire       [17:0]   fixTo_50_dout;
  wire       [17:0]   fixTo_51_dout;
  wire       [17:0]   fixTo_52_dout;
  wire       [17:0]   fixTo_53_dout;
  wire       [35:0]   fixTo_54_dout;
  wire       [35:0]   fixTo_55_dout;
  wire       [17:0]   fixTo_56_dout;
  wire       [17:0]   fixTo_57_dout;
  wire       [17:0]   fixTo_58_dout;
  wire       [17:0]   fixTo_59_dout;
  wire       [35:0]   fixTo_60_dout;
  wire       [35:0]   fixTo_61_dout;
  wire       [17:0]   fixTo_62_dout;
  wire       [17:0]   fixTo_63_dout;
  wire       [17:0]   fixTo_64_dout;
  wire       [17:0]   fixTo_65_dout;
  wire       [35:0]   fixTo_66_dout;
  wire       [35:0]   fixTo_67_dout;
  wire       [17:0]   fixTo_68_dout;
  wire       [17:0]   fixTo_69_dout;
  wire       [17:0]   fixTo_70_dout;
  wire       [17:0]   fixTo_71_dout;
  wire       [35:0]   fixTo_72_dout;
  wire       [35:0]   fixTo_73_dout;
  wire       [17:0]   fixTo_74_dout;
  wire       [17:0]   fixTo_75_dout;
  wire       [17:0]   fixTo_76_dout;
  wire       [17:0]   fixTo_77_dout;
  wire       [35:0]   fixTo_78_dout;
  wire       [35:0]   fixTo_79_dout;
  wire       [17:0]   fixTo_80_dout;
  wire       [17:0]   fixTo_81_dout;
  wire       [17:0]   fixTo_82_dout;
  wire       [17:0]   fixTo_83_dout;
  wire       [35:0]   fixTo_84_dout;
  wire       [35:0]   fixTo_85_dout;
  wire       [17:0]   fixTo_86_dout;
  wire       [17:0]   fixTo_87_dout;
  wire       [17:0]   fixTo_88_dout;
  wire       [17:0]   fixTo_89_dout;
  wire       [35:0]   fixTo_90_dout;
  wire       [35:0]   fixTo_91_dout;
  wire       [17:0]   fixTo_92_dout;
  wire       [17:0]   fixTo_93_dout;
  wire       [17:0]   fixTo_94_dout;
  wire       [17:0]   fixTo_95_dout;
  wire       [35:0]   fixTo_96_dout;
  wire       [35:0]   fixTo_97_dout;
  wire       [17:0]   fixTo_98_dout;
  wire       [17:0]   fixTo_99_dout;
  wire       [17:0]   fixTo_100_dout;
  wire       [17:0]   fixTo_101_dout;
  wire       [35:0]   fixTo_102_dout;
  wire       [35:0]   fixTo_103_dout;
  wire       [17:0]   fixTo_104_dout;
  wire       [17:0]   fixTo_105_dout;
  wire       [17:0]   fixTo_106_dout;
  wire       [17:0]   fixTo_107_dout;
  wire       [35:0]   fixTo_108_dout;
  wire       [35:0]   fixTo_109_dout;
  wire       [17:0]   fixTo_110_dout;
  wire       [17:0]   fixTo_111_dout;
  wire       [17:0]   fixTo_112_dout;
  wire       [17:0]   fixTo_113_dout;
  wire       [35:0]   fixTo_114_dout;
  wire       [35:0]   fixTo_115_dout;
  wire       [17:0]   fixTo_116_dout;
  wire       [17:0]   fixTo_117_dout;
  wire       [17:0]   fixTo_118_dout;
  wire       [17:0]   fixTo_119_dout;
  wire       [35:0]   fixTo_120_dout;
  wire       [35:0]   fixTo_121_dout;
  wire       [17:0]   fixTo_122_dout;
  wire       [17:0]   fixTo_123_dout;
  wire       [17:0]   fixTo_124_dout;
  wire       [17:0]   fixTo_125_dout;
  wire       [35:0]   fixTo_126_dout;
  wire       [35:0]   fixTo_127_dout;
  wire       [17:0]   fixTo_128_dout;
  wire       [17:0]   fixTo_129_dout;
  wire       [17:0]   fixTo_130_dout;
  wire       [17:0]   fixTo_131_dout;
  wire       [35:0]   fixTo_132_dout;
  wire       [35:0]   fixTo_133_dout;
  wire       [17:0]   fixTo_134_dout;
  wire       [17:0]   fixTo_135_dout;
  wire       [17:0]   fixTo_136_dout;
  wire       [17:0]   fixTo_137_dout;
  wire       [35:0]   fixTo_138_dout;
  wire       [35:0]   fixTo_139_dout;
  wire       [17:0]   fixTo_140_dout;
  wire       [17:0]   fixTo_141_dout;
  wire       [17:0]   fixTo_142_dout;
  wire       [17:0]   fixTo_143_dout;
  wire       [35:0]   fixTo_144_dout;
  wire       [35:0]   fixTo_145_dout;
  wire       [17:0]   fixTo_146_dout;
  wire       [17:0]   fixTo_147_dout;
  wire       [17:0]   fixTo_148_dout;
  wire       [17:0]   fixTo_149_dout;
  wire       [35:0]   fixTo_150_dout;
  wire       [35:0]   fixTo_151_dout;
  wire       [17:0]   fixTo_152_dout;
  wire       [17:0]   fixTo_153_dout;
  wire       [17:0]   fixTo_154_dout;
  wire       [17:0]   fixTo_155_dout;
  wire       [35:0]   fixTo_156_dout;
  wire       [35:0]   fixTo_157_dout;
  wire       [17:0]   fixTo_158_dout;
  wire       [17:0]   fixTo_159_dout;
  wire       [17:0]   fixTo_160_dout;
  wire       [17:0]   fixTo_161_dout;
  wire       [35:0]   fixTo_162_dout;
  wire       [35:0]   fixTo_163_dout;
  wire       [17:0]   fixTo_164_dout;
  wire       [17:0]   fixTo_165_dout;
  wire       [17:0]   fixTo_166_dout;
  wire       [17:0]   fixTo_167_dout;
  wire       [35:0]   fixTo_168_dout;
  wire       [35:0]   fixTo_169_dout;
  wire       [17:0]   fixTo_170_dout;
  wire       [17:0]   fixTo_171_dout;
  wire       [17:0]   fixTo_172_dout;
  wire       [17:0]   fixTo_173_dout;
  wire       [35:0]   fixTo_174_dout;
  wire       [35:0]   fixTo_175_dout;
  wire       [17:0]   fixTo_176_dout;
  wire       [17:0]   fixTo_177_dout;
  wire       [17:0]   fixTo_178_dout;
  wire       [17:0]   fixTo_179_dout;
  wire       [35:0]   fixTo_180_dout;
  wire       [35:0]   fixTo_181_dout;
  wire       [17:0]   fixTo_182_dout;
  wire       [17:0]   fixTo_183_dout;
  wire       [17:0]   fixTo_184_dout;
  wire       [17:0]   fixTo_185_dout;
  wire       [35:0]   fixTo_186_dout;
  wire       [35:0]   fixTo_187_dout;
  wire       [17:0]   fixTo_188_dout;
  wire       [17:0]   fixTo_189_dout;
  wire       [17:0]   fixTo_190_dout;
  wire       [17:0]   fixTo_191_dout;
  wire       [35:0]   fixTo_192_dout;
  wire       [35:0]   fixTo_193_dout;
  wire       [17:0]   fixTo_194_dout;
  wire       [17:0]   fixTo_195_dout;
  wire       [17:0]   fixTo_196_dout;
  wire       [17:0]   fixTo_197_dout;
  wire       [35:0]   fixTo_198_dout;
  wire       [35:0]   fixTo_199_dout;
  wire       [17:0]   fixTo_200_dout;
  wire       [17:0]   fixTo_201_dout;
  wire       [17:0]   fixTo_202_dout;
  wire       [17:0]   fixTo_203_dout;
  wire       [35:0]   fixTo_204_dout;
  wire       [35:0]   fixTo_205_dout;
  wire       [17:0]   fixTo_206_dout;
  wire       [17:0]   fixTo_207_dout;
  wire       [17:0]   fixTo_208_dout;
  wire       [17:0]   fixTo_209_dout;
  wire       [35:0]   fixTo_210_dout;
  wire       [35:0]   fixTo_211_dout;
  wire       [17:0]   fixTo_212_dout;
  wire       [17:0]   fixTo_213_dout;
  wire       [17:0]   fixTo_214_dout;
  wire       [17:0]   fixTo_215_dout;
  wire       [35:0]   fixTo_216_dout;
  wire       [35:0]   fixTo_217_dout;
  wire       [17:0]   fixTo_218_dout;
  wire       [17:0]   fixTo_219_dout;
  wire       [17:0]   fixTo_220_dout;
  wire       [17:0]   fixTo_221_dout;
  wire       [35:0]   fixTo_222_dout;
  wire       [35:0]   fixTo_223_dout;
  wire       [17:0]   fixTo_224_dout;
  wire       [17:0]   fixTo_225_dout;
  wire       [17:0]   fixTo_226_dout;
  wire       [17:0]   fixTo_227_dout;
  wire       [35:0]   fixTo_228_dout;
  wire       [35:0]   fixTo_229_dout;
  wire       [17:0]   fixTo_230_dout;
  wire       [17:0]   fixTo_231_dout;
  wire       [17:0]   fixTo_232_dout;
  wire       [17:0]   fixTo_233_dout;
  wire       [35:0]   fixTo_234_dout;
  wire       [35:0]   fixTo_235_dout;
  wire       [17:0]   fixTo_236_dout;
  wire       [17:0]   fixTo_237_dout;
  wire       [17:0]   fixTo_238_dout;
  wire       [17:0]   fixTo_239_dout;
  wire       [35:0]   fixTo_240_dout;
  wire       [35:0]   fixTo_241_dout;
  wire       [17:0]   fixTo_242_dout;
  wire       [17:0]   fixTo_243_dout;
  wire       [17:0]   fixTo_244_dout;
  wire       [17:0]   fixTo_245_dout;
  wire       [35:0]   fixTo_246_dout;
  wire       [35:0]   fixTo_247_dout;
  wire       [17:0]   fixTo_248_dout;
  wire       [17:0]   fixTo_249_dout;
  wire       [17:0]   fixTo_250_dout;
  wire       [17:0]   fixTo_251_dout;
  wire       [35:0]   fixTo_252_dout;
  wire       [35:0]   fixTo_253_dout;
  wire       [17:0]   fixTo_254_dout;
  wire       [17:0]   fixTo_255_dout;
  wire       [17:0]   fixTo_256_dout;
  wire       [17:0]   fixTo_257_dout;
  wire       [35:0]   fixTo_258_dout;
  wire       [35:0]   fixTo_259_dout;
  wire       [17:0]   fixTo_260_dout;
  wire       [17:0]   fixTo_261_dout;
  wire       [17:0]   fixTo_262_dout;
  wire       [17:0]   fixTo_263_dout;
  wire       [35:0]   fixTo_264_dout;
  wire       [35:0]   fixTo_265_dout;
  wire       [17:0]   fixTo_266_dout;
  wire       [17:0]   fixTo_267_dout;
  wire       [17:0]   fixTo_268_dout;
  wire       [17:0]   fixTo_269_dout;
  wire       [35:0]   fixTo_270_dout;
  wire       [35:0]   fixTo_271_dout;
  wire       [17:0]   fixTo_272_dout;
  wire       [17:0]   fixTo_273_dout;
  wire       [17:0]   fixTo_274_dout;
  wire       [17:0]   fixTo_275_dout;
  wire       [35:0]   fixTo_276_dout;
  wire       [35:0]   fixTo_277_dout;
  wire       [17:0]   fixTo_278_dout;
  wire       [17:0]   fixTo_279_dout;
  wire       [17:0]   fixTo_280_dout;
  wire       [17:0]   fixTo_281_dout;
  wire       [35:0]   fixTo_282_dout;
  wire       [35:0]   fixTo_283_dout;
  wire       [17:0]   fixTo_284_dout;
  wire       [17:0]   fixTo_285_dout;
  wire       [17:0]   fixTo_286_dout;
  wire       [17:0]   fixTo_287_dout;
  wire       [35:0]   fixTo_288_dout;
  wire       [35:0]   fixTo_289_dout;
  wire       [17:0]   fixTo_290_dout;
  wire       [17:0]   fixTo_291_dout;
  wire       [17:0]   fixTo_292_dout;
  wire       [17:0]   fixTo_293_dout;
  wire       [35:0]   fixTo_294_dout;
  wire       [35:0]   fixTo_295_dout;
  wire       [17:0]   fixTo_296_dout;
  wire       [17:0]   fixTo_297_dout;
  wire       [17:0]   fixTo_298_dout;
  wire       [17:0]   fixTo_299_dout;
  wire       [35:0]   fixTo_300_dout;
  wire       [35:0]   fixTo_301_dout;
  wire       [17:0]   fixTo_302_dout;
  wire       [17:0]   fixTo_303_dout;
  wire       [17:0]   fixTo_304_dout;
  wire       [17:0]   fixTo_305_dout;
  wire       [35:0]   fixTo_306_dout;
  wire       [35:0]   fixTo_307_dout;
  wire       [17:0]   fixTo_308_dout;
  wire       [17:0]   fixTo_309_dout;
  wire       [17:0]   fixTo_310_dout;
  wire       [17:0]   fixTo_311_dout;
  wire       [35:0]   fixTo_312_dout;
  wire       [35:0]   fixTo_313_dout;
  wire       [17:0]   fixTo_314_dout;
  wire       [17:0]   fixTo_315_dout;
  wire       [17:0]   fixTo_316_dout;
  wire       [17:0]   fixTo_317_dout;
  wire       [35:0]   fixTo_318_dout;
  wire       [35:0]   fixTo_319_dout;
  wire       [17:0]   fixTo_320_dout;
  wire       [17:0]   fixTo_321_dout;
  wire       [17:0]   fixTo_322_dout;
  wire       [17:0]   fixTo_323_dout;
  wire       [35:0]   fixTo_324_dout;
  wire       [35:0]   fixTo_325_dout;
  wire       [17:0]   fixTo_326_dout;
  wire       [17:0]   fixTo_327_dout;
  wire       [17:0]   fixTo_328_dout;
  wire       [17:0]   fixTo_329_dout;
  wire       [35:0]   fixTo_330_dout;
  wire       [35:0]   fixTo_331_dout;
  wire       [17:0]   fixTo_332_dout;
  wire       [17:0]   fixTo_333_dout;
  wire       [17:0]   fixTo_334_dout;
  wire       [17:0]   fixTo_335_dout;
  wire       [35:0]   fixTo_336_dout;
  wire       [35:0]   fixTo_337_dout;
  wire       [17:0]   fixTo_338_dout;
  wire       [17:0]   fixTo_339_dout;
  wire       [17:0]   fixTo_340_dout;
  wire       [17:0]   fixTo_341_dout;
  wire       [35:0]   fixTo_342_dout;
  wire       [35:0]   fixTo_343_dout;
  wire       [17:0]   fixTo_344_dout;
  wire       [17:0]   fixTo_345_dout;
  wire       [17:0]   fixTo_346_dout;
  wire       [17:0]   fixTo_347_dout;
  wire       [35:0]   fixTo_348_dout;
  wire       [35:0]   fixTo_349_dout;
  wire       [17:0]   fixTo_350_dout;
  wire       [17:0]   fixTo_351_dout;
  wire       [17:0]   fixTo_352_dout;
  wire       [17:0]   fixTo_353_dout;
  wire       [35:0]   fixTo_354_dout;
  wire       [35:0]   fixTo_355_dout;
  wire       [17:0]   fixTo_356_dout;
  wire       [17:0]   fixTo_357_dout;
  wire       [17:0]   fixTo_358_dout;
  wire       [17:0]   fixTo_359_dout;
  wire       [35:0]   fixTo_360_dout;
  wire       [35:0]   fixTo_361_dout;
  wire       [17:0]   fixTo_362_dout;
  wire       [17:0]   fixTo_363_dout;
  wire       [17:0]   fixTo_364_dout;
  wire       [17:0]   fixTo_365_dout;
  wire       [35:0]   fixTo_366_dout;
  wire       [35:0]   fixTo_367_dout;
  wire       [17:0]   fixTo_368_dout;
  wire       [17:0]   fixTo_369_dout;
  wire       [17:0]   fixTo_370_dout;
  wire       [17:0]   fixTo_371_dout;
  wire       [35:0]   fixTo_372_dout;
  wire       [35:0]   fixTo_373_dout;
  wire       [17:0]   fixTo_374_dout;
  wire       [17:0]   fixTo_375_dout;
  wire       [17:0]   fixTo_376_dout;
  wire       [17:0]   fixTo_377_dout;
  wire       [35:0]   fixTo_378_dout;
  wire       [35:0]   fixTo_379_dout;
  wire       [17:0]   fixTo_380_dout;
  wire       [17:0]   fixTo_381_dout;
  wire       [17:0]   fixTo_382_dout;
  wire       [17:0]   fixTo_383_dout;
  wire       [35:0]   fixTo_384_dout;
  wire       [35:0]   fixTo_385_dout;
  wire       [17:0]   fixTo_386_dout;
  wire       [17:0]   fixTo_387_dout;
  wire       [17:0]   fixTo_388_dout;
  wire       [17:0]   fixTo_389_dout;
  wire       [35:0]   fixTo_390_dout;
  wire       [35:0]   fixTo_391_dout;
  wire       [17:0]   fixTo_392_dout;
  wire       [17:0]   fixTo_393_dout;
  wire       [17:0]   fixTo_394_dout;
  wire       [17:0]   fixTo_395_dout;
  wire       [35:0]   fixTo_396_dout;
  wire       [35:0]   fixTo_397_dout;
  wire       [17:0]   fixTo_398_dout;
  wire       [17:0]   fixTo_399_dout;
  wire       [17:0]   fixTo_400_dout;
  wire       [17:0]   fixTo_401_dout;
  wire       [35:0]   fixTo_402_dout;
  wire       [35:0]   fixTo_403_dout;
  wire       [17:0]   fixTo_404_dout;
  wire       [17:0]   fixTo_405_dout;
  wire       [17:0]   fixTo_406_dout;
  wire       [17:0]   fixTo_407_dout;
  wire       [35:0]   fixTo_408_dout;
  wire       [35:0]   fixTo_409_dout;
  wire       [17:0]   fixTo_410_dout;
  wire       [17:0]   fixTo_411_dout;
  wire       [17:0]   fixTo_412_dout;
  wire       [17:0]   fixTo_413_dout;
  wire       [35:0]   fixTo_414_dout;
  wire       [35:0]   fixTo_415_dout;
  wire       [17:0]   fixTo_416_dout;
  wire       [17:0]   fixTo_417_dout;
  wire       [17:0]   fixTo_418_dout;
  wire       [17:0]   fixTo_419_dout;
  wire       [35:0]   fixTo_420_dout;
  wire       [35:0]   fixTo_421_dout;
  wire       [17:0]   fixTo_422_dout;
  wire       [17:0]   fixTo_423_dout;
  wire       [17:0]   fixTo_424_dout;
  wire       [17:0]   fixTo_425_dout;
  wire       [35:0]   fixTo_426_dout;
  wire       [35:0]   fixTo_427_dout;
  wire       [17:0]   fixTo_428_dout;
  wire       [17:0]   fixTo_429_dout;
  wire       [17:0]   fixTo_430_dout;
  wire       [17:0]   fixTo_431_dout;
  wire       [35:0]   fixTo_432_dout;
  wire       [35:0]   fixTo_433_dout;
  wire       [17:0]   fixTo_434_dout;
  wire       [17:0]   fixTo_435_dout;
  wire       [17:0]   fixTo_436_dout;
  wire       [17:0]   fixTo_437_dout;
  wire       [35:0]   fixTo_438_dout;
  wire       [35:0]   fixTo_439_dout;
  wire       [17:0]   fixTo_440_dout;
  wire       [17:0]   fixTo_441_dout;
  wire       [17:0]   fixTo_442_dout;
  wire       [17:0]   fixTo_443_dout;
  wire       [35:0]   fixTo_444_dout;
  wire       [35:0]   fixTo_445_dout;
  wire       [17:0]   fixTo_446_dout;
  wire       [17:0]   fixTo_447_dout;
  wire       [17:0]   fixTo_448_dout;
  wire       [17:0]   fixTo_449_dout;
  wire       [35:0]   fixTo_450_dout;
  wire       [35:0]   fixTo_451_dout;
  wire       [17:0]   fixTo_452_dout;
  wire       [17:0]   fixTo_453_dout;
  wire       [17:0]   fixTo_454_dout;
  wire       [17:0]   fixTo_455_dout;
  wire       [35:0]   fixTo_456_dout;
  wire       [35:0]   fixTo_457_dout;
  wire       [17:0]   fixTo_458_dout;
  wire       [17:0]   fixTo_459_dout;
  wire       [17:0]   fixTo_460_dout;
  wire       [17:0]   fixTo_461_dout;
  wire       [35:0]   fixTo_462_dout;
  wire       [35:0]   fixTo_463_dout;
  wire       [17:0]   fixTo_464_dout;
  wire       [17:0]   fixTo_465_dout;
  wire       [17:0]   fixTo_466_dout;
  wire       [17:0]   fixTo_467_dout;
  wire       [35:0]   fixTo_468_dout;
  wire       [35:0]   fixTo_469_dout;
  wire       [17:0]   fixTo_470_dout;
  wire       [17:0]   fixTo_471_dout;
  wire       [17:0]   fixTo_472_dout;
  wire       [17:0]   fixTo_473_dout;
  wire       [35:0]   fixTo_474_dout;
  wire       [35:0]   fixTo_475_dout;
  wire       [17:0]   fixTo_476_dout;
  wire       [17:0]   fixTo_477_dout;
  wire       [17:0]   fixTo_478_dout;
  wire       [17:0]   fixTo_479_dout;
  wire       [35:0]   fixTo_480_dout;
  wire       [35:0]   fixTo_481_dout;
  wire       [17:0]   fixTo_482_dout;
  wire       [17:0]   fixTo_483_dout;
  wire       [17:0]   fixTo_484_dout;
  wire       [17:0]   fixTo_485_dout;
  wire       [35:0]   fixTo_486_dout;
  wire       [35:0]   fixTo_487_dout;
  wire       [17:0]   fixTo_488_dout;
  wire       [17:0]   fixTo_489_dout;
  wire       [17:0]   fixTo_490_dout;
  wire       [17:0]   fixTo_491_dout;
  wire       [35:0]   fixTo_492_dout;
  wire       [35:0]   fixTo_493_dout;
  wire       [17:0]   fixTo_494_dout;
  wire       [17:0]   fixTo_495_dout;
  wire       [17:0]   fixTo_496_dout;
  wire       [17:0]   fixTo_497_dout;
  wire       [35:0]   fixTo_498_dout;
  wire       [35:0]   fixTo_499_dout;
  wire       [17:0]   fixTo_500_dout;
  wire       [17:0]   fixTo_501_dout;
  wire       [17:0]   fixTo_502_dout;
  wire       [17:0]   fixTo_503_dout;
  wire       [35:0]   fixTo_504_dout;
  wire       [35:0]   fixTo_505_dout;
  wire       [17:0]   fixTo_506_dout;
  wire       [17:0]   fixTo_507_dout;
  wire       [17:0]   fixTo_508_dout;
  wire       [17:0]   fixTo_509_dout;
  wire       [35:0]   fixTo_510_dout;
  wire       [35:0]   fixTo_511_dout;
  wire       [17:0]   fixTo_512_dout;
  wire       [17:0]   fixTo_513_dout;
  wire       [17:0]   fixTo_514_dout;
  wire       [17:0]   fixTo_515_dout;
  wire       [35:0]   fixTo_516_dout;
  wire       [35:0]   fixTo_517_dout;
  wire       [17:0]   fixTo_518_dout;
  wire       [17:0]   fixTo_519_dout;
  wire       [17:0]   fixTo_520_dout;
  wire       [17:0]   fixTo_521_dout;
  wire       [35:0]   fixTo_522_dout;
  wire       [35:0]   fixTo_523_dout;
  wire       [17:0]   fixTo_524_dout;
  wire       [17:0]   fixTo_525_dout;
  wire       [17:0]   fixTo_526_dout;
  wire       [17:0]   fixTo_527_dout;
  wire       [35:0]   fixTo_528_dout;
  wire       [35:0]   fixTo_529_dout;
  wire       [17:0]   fixTo_530_dout;
  wire       [17:0]   fixTo_531_dout;
  wire       [17:0]   fixTo_532_dout;
  wire       [17:0]   fixTo_533_dout;
  wire       [35:0]   fixTo_534_dout;
  wire       [35:0]   fixTo_535_dout;
  wire       [17:0]   fixTo_536_dout;
  wire       [17:0]   fixTo_537_dout;
  wire       [17:0]   fixTo_538_dout;
  wire       [17:0]   fixTo_539_dout;
  wire       [35:0]   fixTo_540_dout;
  wire       [35:0]   fixTo_541_dout;
  wire       [17:0]   fixTo_542_dout;
  wire       [17:0]   fixTo_543_dout;
  wire       [17:0]   fixTo_544_dout;
  wire       [17:0]   fixTo_545_dout;
  wire       [35:0]   fixTo_546_dout;
  wire       [35:0]   fixTo_547_dout;
  wire       [17:0]   fixTo_548_dout;
  wire       [17:0]   fixTo_549_dout;
  wire       [17:0]   fixTo_550_dout;
  wire       [17:0]   fixTo_551_dout;
  wire       [35:0]   fixTo_552_dout;
  wire       [35:0]   fixTo_553_dout;
  wire       [17:0]   fixTo_554_dout;
  wire       [17:0]   fixTo_555_dout;
  wire       [17:0]   fixTo_556_dout;
  wire       [17:0]   fixTo_557_dout;
  wire       [35:0]   fixTo_558_dout;
  wire       [35:0]   fixTo_559_dout;
  wire       [17:0]   fixTo_560_dout;
  wire       [17:0]   fixTo_561_dout;
  wire       [17:0]   fixTo_562_dout;
  wire       [17:0]   fixTo_563_dout;
  wire       [35:0]   fixTo_564_dout;
  wire       [35:0]   fixTo_565_dout;
  wire       [17:0]   fixTo_566_dout;
  wire       [17:0]   fixTo_567_dout;
  wire       [17:0]   fixTo_568_dout;
  wire       [17:0]   fixTo_569_dout;
  wire       [35:0]   fixTo_570_dout;
  wire       [35:0]   fixTo_571_dout;
  wire       [17:0]   fixTo_572_dout;
  wire       [17:0]   fixTo_573_dout;
  wire       [17:0]   fixTo_574_dout;
  wire       [17:0]   fixTo_575_dout;
  wire       [35:0]   fixTo_576_dout;
  wire       [35:0]   fixTo_577_dout;
  wire       [17:0]   fixTo_578_dout;
  wire       [17:0]   fixTo_579_dout;
  wire       [17:0]   fixTo_580_dout;
  wire       [17:0]   fixTo_581_dout;
  wire       [35:0]   fixTo_582_dout;
  wire       [35:0]   fixTo_583_dout;
  wire       [17:0]   fixTo_584_dout;
  wire       [17:0]   fixTo_585_dout;
  wire       [17:0]   fixTo_586_dout;
  wire       [17:0]   fixTo_587_dout;
  wire       [35:0]   fixTo_588_dout;
  wire       [35:0]   fixTo_589_dout;
  wire       [17:0]   fixTo_590_dout;
  wire       [17:0]   fixTo_591_dout;
  wire       [17:0]   fixTo_592_dout;
  wire       [17:0]   fixTo_593_dout;
  wire       [35:0]   fixTo_594_dout;
  wire       [35:0]   fixTo_595_dout;
  wire       [17:0]   fixTo_596_dout;
  wire       [17:0]   fixTo_597_dout;
  wire       [17:0]   fixTo_598_dout;
  wire       [17:0]   fixTo_599_dout;
  wire       [35:0]   fixTo_600_dout;
  wire       [35:0]   fixTo_601_dout;
  wire       [17:0]   fixTo_602_dout;
  wire       [17:0]   fixTo_603_dout;
  wire       [17:0]   fixTo_604_dout;
  wire       [17:0]   fixTo_605_dout;
  wire       [35:0]   fixTo_606_dout;
  wire       [35:0]   fixTo_607_dout;
  wire       [17:0]   fixTo_608_dout;
  wire       [17:0]   fixTo_609_dout;
  wire       [17:0]   fixTo_610_dout;
  wire       [17:0]   fixTo_611_dout;
  wire       [35:0]   fixTo_612_dout;
  wire       [35:0]   fixTo_613_dout;
  wire       [17:0]   fixTo_614_dout;
  wire       [17:0]   fixTo_615_dout;
  wire       [17:0]   fixTo_616_dout;
  wire       [17:0]   fixTo_617_dout;
  wire       [35:0]   fixTo_618_dout;
  wire       [35:0]   fixTo_619_dout;
  wire       [17:0]   fixTo_620_dout;
  wire       [17:0]   fixTo_621_dout;
  wire       [17:0]   fixTo_622_dout;
  wire       [17:0]   fixTo_623_dout;
  wire       [35:0]   fixTo_624_dout;
  wire       [35:0]   fixTo_625_dout;
  wire       [17:0]   fixTo_626_dout;
  wire       [17:0]   fixTo_627_dout;
  wire       [17:0]   fixTo_628_dout;
  wire       [17:0]   fixTo_629_dout;
  wire       [35:0]   fixTo_630_dout;
  wire       [35:0]   fixTo_631_dout;
  wire       [17:0]   fixTo_632_dout;
  wire       [17:0]   fixTo_633_dout;
  wire       [17:0]   fixTo_634_dout;
  wire       [17:0]   fixTo_635_dout;
  wire       [35:0]   fixTo_636_dout;
  wire       [35:0]   fixTo_637_dout;
  wire       [17:0]   fixTo_638_dout;
  wire       [17:0]   fixTo_639_dout;
  wire       [17:0]   fixTo_640_dout;
  wire       [17:0]   fixTo_641_dout;
  wire       [35:0]   fixTo_642_dout;
  wire       [35:0]   fixTo_643_dout;
  wire       [17:0]   fixTo_644_dout;
  wire       [17:0]   fixTo_645_dout;
  wire       [17:0]   fixTo_646_dout;
  wire       [17:0]   fixTo_647_dout;
  wire       [35:0]   fixTo_648_dout;
  wire       [35:0]   fixTo_649_dout;
  wire       [17:0]   fixTo_650_dout;
  wire       [17:0]   fixTo_651_dout;
  wire       [17:0]   fixTo_652_dout;
  wire       [17:0]   fixTo_653_dout;
  wire       [35:0]   fixTo_654_dout;
  wire       [35:0]   fixTo_655_dout;
  wire       [17:0]   fixTo_656_dout;
  wire       [17:0]   fixTo_657_dout;
  wire       [17:0]   fixTo_658_dout;
  wire       [17:0]   fixTo_659_dout;
  wire       [35:0]   fixTo_660_dout;
  wire       [35:0]   fixTo_661_dout;
  wire       [17:0]   fixTo_662_dout;
  wire       [17:0]   fixTo_663_dout;
  wire       [17:0]   fixTo_664_dout;
  wire       [17:0]   fixTo_665_dout;
  wire       [35:0]   fixTo_666_dout;
  wire       [35:0]   fixTo_667_dout;
  wire       [17:0]   fixTo_668_dout;
  wire       [17:0]   fixTo_669_dout;
  wire       [17:0]   fixTo_670_dout;
  wire       [17:0]   fixTo_671_dout;
  wire       [35:0]   fixTo_672_dout;
  wire       [35:0]   fixTo_673_dout;
  wire       [17:0]   fixTo_674_dout;
  wire       [17:0]   fixTo_675_dout;
  wire       [17:0]   fixTo_676_dout;
  wire       [17:0]   fixTo_677_dout;
  wire       [35:0]   fixTo_678_dout;
  wire       [35:0]   fixTo_679_dout;
  wire       [17:0]   fixTo_680_dout;
  wire       [17:0]   fixTo_681_dout;
  wire       [17:0]   fixTo_682_dout;
  wire       [17:0]   fixTo_683_dout;
  wire       [35:0]   fixTo_684_dout;
  wire       [35:0]   fixTo_685_dout;
  wire       [17:0]   fixTo_686_dout;
  wire       [17:0]   fixTo_687_dout;
  wire       [17:0]   fixTo_688_dout;
  wire       [17:0]   fixTo_689_dout;
  wire       [35:0]   fixTo_690_dout;
  wire       [35:0]   fixTo_691_dout;
  wire       [17:0]   fixTo_692_dout;
  wire       [17:0]   fixTo_693_dout;
  wire       [17:0]   fixTo_694_dout;
  wire       [17:0]   fixTo_695_dout;
  wire       [35:0]   fixTo_696_dout;
  wire       [35:0]   fixTo_697_dout;
  wire       [17:0]   fixTo_698_dout;
  wire       [17:0]   fixTo_699_dout;
  wire       [17:0]   fixTo_700_dout;
  wire       [17:0]   fixTo_701_dout;
  wire       [35:0]   fixTo_702_dout;
  wire       [35:0]   fixTo_703_dout;
  wire       [17:0]   fixTo_704_dout;
  wire       [17:0]   fixTo_705_dout;
  wire       [17:0]   fixTo_706_dout;
  wire       [17:0]   fixTo_707_dout;
  wire       [35:0]   fixTo_708_dout;
  wire       [35:0]   fixTo_709_dout;
  wire       [17:0]   fixTo_710_dout;
  wire       [17:0]   fixTo_711_dout;
  wire       [17:0]   fixTo_712_dout;
  wire       [17:0]   fixTo_713_dout;
  wire       [35:0]   fixTo_714_dout;
  wire       [35:0]   fixTo_715_dout;
  wire       [17:0]   fixTo_716_dout;
  wire       [17:0]   fixTo_717_dout;
  wire       [17:0]   fixTo_718_dout;
  wire       [17:0]   fixTo_719_dout;
  wire       [35:0]   fixTo_720_dout;
  wire       [35:0]   fixTo_721_dout;
  wire       [17:0]   fixTo_722_dout;
  wire       [17:0]   fixTo_723_dout;
  wire       [17:0]   fixTo_724_dout;
  wire       [17:0]   fixTo_725_dout;
  wire       [35:0]   fixTo_726_dout;
  wire       [35:0]   fixTo_727_dout;
  wire       [17:0]   fixTo_728_dout;
  wire       [17:0]   fixTo_729_dout;
  wire       [17:0]   fixTo_730_dout;
  wire       [17:0]   fixTo_731_dout;
  wire       [35:0]   fixTo_732_dout;
  wire       [35:0]   fixTo_733_dout;
  wire       [17:0]   fixTo_734_dout;
  wire       [17:0]   fixTo_735_dout;
  wire       [17:0]   fixTo_736_dout;
  wire       [17:0]   fixTo_737_dout;
  wire       [35:0]   fixTo_738_dout;
  wire       [35:0]   fixTo_739_dout;
  wire       [17:0]   fixTo_740_dout;
  wire       [17:0]   fixTo_741_dout;
  wire       [17:0]   fixTo_742_dout;
  wire       [17:0]   fixTo_743_dout;
  wire       [35:0]   fixTo_744_dout;
  wire       [35:0]   fixTo_745_dout;
  wire       [17:0]   fixTo_746_dout;
  wire       [17:0]   fixTo_747_dout;
  wire       [17:0]   fixTo_748_dout;
  wire       [17:0]   fixTo_749_dout;
  wire       [35:0]   fixTo_750_dout;
  wire       [35:0]   fixTo_751_dout;
  wire       [17:0]   fixTo_752_dout;
  wire       [17:0]   fixTo_753_dout;
  wire       [17:0]   fixTo_754_dout;
  wire       [17:0]   fixTo_755_dout;
  wire       [35:0]   fixTo_756_dout;
  wire       [35:0]   fixTo_757_dout;
  wire       [17:0]   fixTo_758_dout;
  wire       [17:0]   fixTo_759_dout;
  wire       [17:0]   fixTo_760_dout;
  wire       [17:0]   fixTo_761_dout;
  wire       [35:0]   fixTo_762_dout;
  wire       [35:0]   fixTo_763_dout;
  wire       [17:0]   fixTo_764_dout;
  wire       [17:0]   fixTo_765_dout;
  wire       [17:0]   fixTo_766_dout;
  wire       [17:0]   fixTo_767_dout;
  wire       [35:0]   fixTo_768_dout;
  wire       [35:0]   fixTo_769_dout;
  wire       [17:0]   fixTo_770_dout;
  wire       [17:0]   fixTo_771_dout;
  wire       [17:0]   fixTo_772_dout;
  wire       [17:0]   fixTo_773_dout;
  wire       [35:0]   fixTo_774_dout;
  wire       [35:0]   fixTo_775_dout;
  wire       [17:0]   fixTo_776_dout;
  wire       [17:0]   fixTo_777_dout;
  wire       [17:0]   fixTo_778_dout;
  wire       [17:0]   fixTo_779_dout;
  wire       [35:0]   fixTo_780_dout;
  wire       [35:0]   fixTo_781_dout;
  wire       [17:0]   fixTo_782_dout;
  wire       [17:0]   fixTo_783_dout;
  wire       [17:0]   fixTo_784_dout;
  wire       [17:0]   fixTo_785_dout;
  wire       [35:0]   fixTo_786_dout;
  wire       [35:0]   fixTo_787_dout;
  wire       [17:0]   fixTo_788_dout;
  wire       [17:0]   fixTo_789_dout;
  wire       [17:0]   fixTo_790_dout;
  wire       [17:0]   fixTo_791_dout;
  wire       [35:0]   fixTo_792_dout;
  wire       [35:0]   fixTo_793_dout;
  wire       [17:0]   fixTo_794_dout;
  wire       [17:0]   fixTo_795_dout;
  wire       [17:0]   fixTo_796_dout;
  wire       [17:0]   fixTo_797_dout;
  wire       [35:0]   fixTo_798_dout;
  wire       [35:0]   fixTo_799_dout;
  wire       [17:0]   fixTo_800_dout;
  wire       [17:0]   fixTo_801_dout;
  wire       [17:0]   fixTo_802_dout;
  wire       [17:0]   fixTo_803_dout;
  wire       [35:0]   fixTo_804_dout;
  wire       [35:0]   fixTo_805_dout;
  wire       [17:0]   fixTo_806_dout;
  wire       [17:0]   fixTo_807_dout;
  wire       [17:0]   fixTo_808_dout;
  wire       [17:0]   fixTo_809_dout;
  wire       [35:0]   fixTo_810_dout;
  wire       [35:0]   fixTo_811_dout;
  wire       [17:0]   fixTo_812_dout;
  wire       [17:0]   fixTo_813_dout;
  wire       [17:0]   fixTo_814_dout;
  wire       [17:0]   fixTo_815_dout;
  wire       [35:0]   fixTo_816_dout;
  wire       [35:0]   fixTo_817_dout;
  wire       [17:0]   fixTo_818_dout;
  wire       [17:0]   fixTo_819_dout;
  wire       [17:0]   fixTo_820_dout;
  wire       [17:0]   fixTo_821_dout;
  wire       [35:0]   fixTo_822_dout;
  wire       [35:0]   fixTo_823_dout;
  wire       [17:0]   fixTo_824_dout;
  wire       [17:0]   fixTo_825_dout;
  wire       [17:0]   fixTo_826_dout;
  wire       [17:0]   fixTo_827_dout;
  wire       [35:0]   fixTo_828_dout;
  wire       [35:0]   fixTo_829_dout;
  wire       [17:0]   fixTo_830_dout;
  wire       [17:0]   fixTo_831_dout;
  wire       [17:0]   fixTo_832_dout;
  wire       [17:0]   fixTo_833_dout;
  wire       [35:0]   fixTo_834_dout;
  wire       [35:0]   fixTo_835_dout;
  wire       [17:0]   fixTo_836_dout;
  wire       [17:0]   fixTo_837_dout;
  wire       [17:0]   fixTo_838_dout;
  wire       [17:0]   fixTo_839_dout;
  wire       [35:0]   fixTo_840_dout;
  wire       [35:0]   fixTo_841_dout;
  wire       [17:0]   fixTo_842_dout;
  wire       [17:0]   fixTo_843_dout;
  wire       [17:0]   fixTo_844_dout;
  wire       [17:0]   fixTo_845_dout;
  wire       [35:0]   fixTo_846_dout;
  wire       [35:0]   fixTo_847_dout;
  wire       [17:0]   fixTo_848_dout;
  wire       [17:0]   fixTo_849_dout;
  wire       [17:0]   fixTo_850_dout;
  wire       [17:0]   fixTo_851_dout;
  wire       [35:0]   fixTo_852_dout;
  wire       [35:0]   fixTo_853_dout;
  wire       [17:0]   fixTo_854_dout;
  wire       [17:0]   fixTo_855_dout;
  wire       [17:0]   fixTo_856_dout;
  wire       [17:0]   fixTo_857_dout;
  wire       [35:0]   fixTo_858_dout;
  wire       [35:0]   fixTo_859_dout;
  wire       [17:0]   fixTo_860_dout;
  wire       [17:0]   fixTo_861_dout;
  wire       [17:0]   fixTo_862_dout;
  wire       [17:0]   fixTo_863_dout;
  wire       [35:0]   fixTo_864_dout;
  wire       [35:0]   fixTo_865_dout;
  wire       [17:0]   fixTo_866_dout;
  wire       [17:0]   fixTo_867_dout;
  wire       [17:0]   fixTo_868_dout;
  wire       [17:0]   fixTo_869_dout;
  wire       [35:0]   fixTo_870_dout;
  wire       [35:0]   fixTo_871_dout;
  wire       [17:0]   fixTo_872_dout;
  wire       [17:0]   fixTo_873_dout;
  wire       [17:0]   fixTo_874_dout;
  wire       [17:0]   fixTo_875_dout;
  wire       [35:0]   fixTo_876_dout;
  wire       [35:0]   fixTo_877_dout;
  wire       [17:0]   fixTo_878_dout;
  wire       [17:0]   fixTo_879_dout;
  wire       [17:0]   fixTo_880_dout;
  wire       [17:0]   fixTo_881_dout;
  wire       [35:0]   fixTo_882_dout;
  wire       [35:0]   fixTo_883_dout;
  wire       [17:0]   fixTo_884_dout;
  wire       [17:0]   fixTo_885_dout;
  wire       [17:0]   fixTo_886_dout;
  wire       [17:0]   fixTo_887_dout;
  wire       [35:0]   fixTo_888_dout;
  wire       [35:0]   fixTo_889_dout;
  wire       [17:0]   fixTo_890_dout;
  wire       [17:0]   fixTo_891_dout;
  wire       [17:0]   fixTo_892_dout;
  wire       [17:0]   fixTo_893_dout;
  wire       [35:0]   fixTo_894_dout;
  wire       [35:0]   fixTo_895_dout;
  wire       [17:0]   fixTo_896_dout;
  wire       [17:0]   fixTo_897_dout;
  wire       [17:0]   fixTo_898_dout;
  wire       [17:0]   fixTo_899_dout;
  wire       [35:0]   fixTo_900_dout;
  wire       [35:0]   fixTo_901_dout;
  wire       [17:0]   fixTo_902_dout;
  wire       [17:0]   fixTo_903_dout;
  wire       [17:0]   fixTo_904_dout;
  wire       [17:0]   fixTo_905_dout;
  wire       [35:0]   fixTo_906_dout;
  wire       [35:0]   fixTo_907_dout;
  wire       [17:0]   fixTo_908_dout;
  wire       [17:0]   fixTo_909_dout;
  wire       [17:0]   fixTo_910_dout;
  wire       [17:0]   fixTo_911_dout;
  wire       [35:0]   fixTo_912_dout;
  wire       [35:0]   fixTo_913_dout;
  wire       [17:0]   fixTo_914_dout;
  wire       [17:0]   fixTo_915_dout;
  wire       [17:0]   fixTo_916_dout;
  wire       [17:0]   fixTo_917_dout;
  wire       [35:0]   fixTo_918_dout;
  wire       [35:0]   fixTo_919_dout;
  wire       [17:0]   fixTo_920_dout;
  wire       [17:0]   fixTo_921_dout;
  wire       [17:0]   fixTo_922_dout;
  wire       [17:0]   fixTo_923_dout;
  wire       [35:0]   fixTo_924_dout;
  wire       [35:0]   fixTo_925_dout;
  wire       [17:0]   fixTo_926_dout;
  wire       [17:0]   fixTo_927_dout;
  wire       [17:0]   fixTo_928_dout;
  wire       [17:0]   fixTo_929_dout;
  wire       [35:0]   fixTo_930_dout;
  wire       [35:0]   fixTo_931_dout;
  wire       [17:0]   fixTo_932_dout;
  wire       [17:0]   fixTo_933_dout;
  wire       [17:0]   fixTo_934_dout;
  wire       [17:0]   fixTo_935_dout;
  wire       [35:0]   fixTo_936_dout;
  wire       [35:0]   fixTo_937_dout;
  wire       [17:0]   fixTo_938_dout;
  wire       [17:0]   fixTo_939_dout;
  wire       [17:0]   fixTo_940_dout;
  wire       [17:0]   fixTo_941_dout;
  wire       [35:0]   fixTo_942_dout;
  wire       [35:0]   fixTo_943_dout;
  wire       [17:0]   fixTo_944_dout;
  wire       [17:0]   fixTo_945_dout;
  wire       [17:0]   fixTo_946_dout;
  wire       [17:0]   fixTo_947_dout;
  wire       [35:0]   fixTo_948_dout;
  wire       [35:0]   fixTo_949_dout;
  wire       [17:0]   fixTo_950_dout;
  wire       [17:0]   fixTo_951_dout;
  wire       [17:0]   fixTo_952_dout;
  wire       [17:0]   fixTo_953_dout;
  wire       [35:0]   fixTo_954_dout;
  wire       [35:0]   fixTo_955_dout;
  wire       [17:0]   fixTo_956_dout;
  wire       [17:0]   fixTo_957_dout;
  wire       [17:0]   fixTo_958_dout;
  wire       [17:0]   fixTo_959_dout;
  wire       [35:0]   fixTo_960_dout;
  wire       [35:0]   fixTo_961_dout;
  wire       [17:0]   fixTo_962_dout;
  wire       [17:0]   fixTo_963_dout;
  wire       [17:0]   fixTo_964_dout;
  wire       [17:0]   fixTo_965_dout;
  wire       [35:0]   fixTo_966_dout;
  wire       [35:0]   fixTo_967_dout;
  wire       [17:0]   fixTo_968_dout;
  wire       [17:0]   fixTo_969_dout;
  wire       [17:0]   fixTo_970_dout;
  wire       [17:0]   fixTo_971_dout;
  wire       [35:0]   fixTo_972_dout;
  wire       [35:0]   fixTo_973_dout;
  wire       [17:0]   fixTo_974_dout;
  wire       [17:0]   fixTo_975_dout;
  wire       [17:0]   fixTo_976_dout;
  wire       [17:0]   fixTo_977_dout;
  wire       [35:0]   fixTo_978_dout;
  wire       [35:0]   fixTo_979_dout;
  wire       [17:0]   fixTo_980_dout;
  wire       [17:0]   fixTo_981_dout;
  wire       [17:0]   fixTo_982_dout;
  wire       [17:0]   fixTo_983_dout;
  wire       [35:0]   fixTo_984_dout;
  wire       [35:0]   fixTo_985_dout;
  wire       [17:0]   fixTo_986_dout;
  wire       [17:0]   fixTo_987_dout;
  wire       [17:0]   fixTo_988_dout;
  wire       [17:0]   fixTo_989_dout;
  wire       [35:0]   fixTo_990_dout;
  wire       [35:0]   fixTo_991_dout;
  wire       [17:0]   fixTo_992_dout;
  wire       [17:0]   fixTo_993_dout;
  wire       [17:0]   fixTo_994_dout;
  wire       [17:0]   fixTo_995_dout;
  wire       [35:0]   fixTo_996_dout;
  wire       [35:0]   fixTo_997_dout;
  wire       [17:0]   fixTo_998_dout;
  wire       [17:0]   fixTo_999_dout;
  wire       [17:0]   fixTo_1000_dout;
  wire       [17:0]   fixTo_1001_dout;
  wire       [35:0]   fixTo_1002_dout;
  wire       [35:0]   fixTo_1003_dout;
  wire       [17:0]   fixTo_1004_dout;
  wire       [17:0]   fixTo_1005_dout;
  wire       [17:0]   fixTo_1006_dout;
  wire       [17:0]   fixTo_1007_dout;
  wire       [35:0]   fixTo_1008_dout;
  wire       [35:0]   fixTo_1009_dout;
  wire       [17:0]   fixTo_1010_dout;
  wire       [17:0]   fixTo_1011_dout;
  wire       [17:0]   fixTo_1012_dout;
  wire       [17:0]   fixTo_1013_dout;
  wire       [35:0]   fixTo_1014_dout;
  wire       [35:0]   fixTo_1015_dout;
  wire       [17:0]   fixTo_1016_dout;
  wire       [17:0]   fixTo_1017_dout;
  wire       [17:0]   fixTo_1018_dout;
  wire       [17:0]   fixTo_1019_dout;
  wire       [35:0]   fixTo_1020_dout;
  wire       [35:0]   fixTo_1021_dout;
  wire       [17:0]   fixTo_1022_dout;
  wire       [17:0]   fixTo_1023_dout;
  wire       [17:0]   fixTo_1024_dout;
  wire       [17:0]   fixTo_1025_dout;
  wire       [35:0]   fixTo_1026_dout;
  wire       [35:0]   fixTo_1027_dout;
  wire       [17:0]   fixTo_1028_dout;
  wire       [17:0]   fixTo_1029_dout;
  wire       [17:0]   fixTo_1030_dout;
  wire       [17:0]   fixTo_1031_dout;
  wire       [35:0]   fixTo_1032_dout;
  wire       [35:0]   fixTo_1033_dout;
  wire       [17:0]   fixTo_1034_dout;
  wire       [17:0]   fixTo_1035_dout;
  wire       [17:0]   fixTo_1036_dout;
  wire       [17:0]   fixTo_1037_dout;
  wire       [35:0]   fixTo_1038_dout;
  wire       [35:0]   fixTo_1039_dout;
  wire       [17:0]   fixTo_1040_dout;
  wire       [17:0]   fixTo_1041_dout;
  wire       [17:0]   fixTo_1042_dout;
  wire       [17:0]   fixTo_1043_dout;
  wire       [35:0]   fixTo_1044_dout;
  wire       [35:0]   fixTo_1045_dout;
  wire       [17:0]   fixTo_1046_dout;
  wire       [17:0]   fixTo_1047_dout;
  wire       [17:0]   fixTo_1048_dout;
  wire       [17:0]   fixTo_1049_dout;
  wire       [35:0]   fixTo_1050_dout;
  wire       [35:0]   fixTo_1051_dout;
  wire       [17:0]   fixTo_1052_dout;
  wire       [17:0]   fixTo_1053_dout;
  wire       [17:0]   fixTo_1054_dout;
  wire       [17:0]   fixTo_1055_dout;
  wire       [35:0]   fixTo_1056_dout;
  wire       [35:0]   fixTo_1057_dout;
  wire       [17:0]   fixTo_1058_dout;
  wire       [17:0]   fixTo_1059_dout;
  wire       [17:0]   fixTo_1060_dout;
  wire       [17:0]   fixTo_1061_dout;
  wire       [35:0]   fixTo_1062_dout;
  wire       [35:0]   fixTo_1063_dout;
  wire       [17:0]   fixTo_1064_dout;
  wire       [17:0]   fixTo_1065_dout;
  wire       [17:0]   fixTo_1066_dout;
  wire       [17:0]   fixTo_1067_dout;
  wire       [35:0]   fixTo_1068_dout;
  wire       [35:0]   fixTo_1069_dout;
  wire       [17:0]   fixTo_1070_dout;
  wire       [17:0]   fixTo_1071_dout;
  wire       [17:0]   fixTo_1072_dout;
  wire       [17:0]   fixTo_1073_dout;
  wire       [35:0]   fixTo_1074_dout;
  wire       [35:0]   fixTo_1075_dout;
  wire       [17:0]   fixTo_1076_dout;
  wire       [17:0]   fixTo_1077_dout;
  wire       [17:0]   fixTo_1078_dout;
  wire       [17:0]   fixTo_1079_dout;
  wire       [35:0]   fixTo_1080_dout;
  wire       [35:0]   fixTo_1081_dout;
  wire       [17:0]   fixTo_1082_dout;
  wire       [17:0]   fixTo_1083_dout;
  wire       [17:0]   fixTo_1084_dout;
  wire       [17:0]   fixTo_1085_dout;
  wire       [35:0]   fixTo_1086_dout;
  wire       [35:0]   fixTo_1087_dout;
  wire       [17:0]   fixTo_1088_dout;
  wire       [17:0]   fixTo_1089_dout;
  wire       [17:0]   fixTo_1090_dout;
  wire       [17:0]   fixTo_1091_dout;
  wire       [35:0]   fixTo_1092_dout;
  wire       [35:0]   fixTo_1093_dout;
  wire       [17:0]   fixTo_1094_dout;
  wire       [17:0]   fixTo_1095_dout;
  wire       [17:0]   fixTo_1096_dout;
  wire       [17:0]   fixTo_1097_dout;
  wire       [35:0]   fixTo_1098_dout;
  wire       [35:0]   fixTo_1099_dout;
  wire       [17:0]   fixTo_1100_dout;
  wire       [17:0]   fixTo_1101_dout;
  wire       [17:0]   fixTo_1102_dout;
  wire       [17:0]   fixTo_1103_dout;
  wire       [35:0]   fixTo_1104_dout;
  wire       [35:0]   fixTo_1105_dout;
  wire       [17:0]   fixTo_1106_dout;
  wire       [17:0]   fixTo_1107_dout;
  wire       [17:0]   fixTo_1108_dout;
  wire       [17:0]   fixTo_1109_dout;
  wire       [35:0]   fixTo_1110_dout;
  wire       [35:0]   fixTo_1111_dout;
  wire       [17:0]   fixTo_1112_dout;
  wire       [17:0]   fixTo_1113_dout;
  wire       [17:0]   fixTo_1114_dout;
  wire       [17:0]   fixTo_1115_dout;
  wire       [35:0]   fixTo_1116_dout;
  wire       [35:0]   fixTo_1117_dout;
  wire       [17:0]   fixTo_1118_dout;
  wire       [17:0]   fixTo_1119_dout;
  wire       [17:0]   fixTo_1120_dout;
  wire       [17:0]   fixTo_1121_dout;
  wire       [35:0]   fixTo_1122_dout;
  wire       [35:0]   fixTo_1123_dout;
  wire       [17:0]   fixTo_1124_dout;
  wire       [17:0]   fixTo_1125_dout;
  wire       [17:0]   fixTo_1126_dout;
  wire       [17:0]   fixTo_1127_dout;
  wire       [35:0]   fixTo_1128_dout;
  wire       [35:0]   fixTo_1129_dout;
  wire       [17:0]   fixTo_1130_dout;
  wire       [17:0]   fixTo_1131_dout;
  wire       [17:0]   fixTo_1132_dout;
  wire       [17:0]   fixTo_1133_dout;
  wire       [35:0]   fixTo_1134_dout;
  wire       [35:0]   fixTo_1135_dout;
  wire       [17:0]   fixTo_1136_dout;
  wire       [17:0]   fixTo_1137_dout;
  wire       [17:0]   fixTo_1138_dout;
  wire       [17:0]   fixTo_1139_dout;
  wire       [35:0]   fixTo_1140_dout;
  wire       [35:0]   fixTo_1141_dout;
  wire       [17:0]   fixTo_1142_dout;
  wire       [17:0]   fixTo_1143_dout;
  wire       [17:0]   fixTo_1144_dout;
  wire       [17:0]   fixTo_1145_dout;
  wire       [35:0]   fixTo_1146_dout;
  wire       [35:0]   fixTo_1147_dout;
  wire       [17:0]   fixTo_1148_dout;
  wire       [17:0]   fixTo_1149_dout;
  wire       [17:0]   fixTo_1150_dout;
  wire       [17:0]   fixTo_1151_dout;
  wire       [17:0]   _zz_2113;
  wire       [35:0]   _zz_2114;
  wire       [35:0]   _zz_2115;
  wire       [17:0]   _zz_2116;
  wire       [35:0]   _zz_2117;
  wire       [35:0]   _zz_2118;
  wire       [35:0]   _zz_2119;
  wire       [17:0]   _zz_2120;
  wire       [35:0]   _zz_2121;
  wire       [35:0]   _zz_2122;
  wire       [35:0]   _zz_2123;
  wire       [35:0]   _zz_2124;
  wire       [35:0]   _zz_2125;
  wire       [35:0]   _zz_2126;
  wire       [26:0]   _zz_2127;
  wire       [35:0]   _zz_2128;
  wire       [17:0]   _zz_2129;
  wire       [35:0]   _zz_2130;
  wire       [35:0]   _zz_2131;
  wire       [35:0]   _zz_2132;
  wire       [35:0]   _zz_2133;
  wire       [35:0]   _zz_2134;
  wire       [26:0]   _zz_2135;
  wire       [35:0]   _zz_2136;
  wire       [17:0]   _zz_2137;
  wire       [35:0]   _zz_2138;
  wire       [35:0]   _zz_2139;
  wire       [35:0]   _zz_2140;
  wire       [35:0]   _zz_2141;
  wire       [35:0]   _zz_2142;
  wire       [26:0]   _zz_2143;
  wire       [35:0]   _zz_2144;
  wire       [17:0]   _zz_2145;
  wire       [35:0]   _zz_2146;
  wire       [35:0]   _zz_2147;
  wire       [35:0]   _zz_2148;
  wire       [35:0]   _zz_2149;
  wire       [35:0]   _zz_2150;
  wire       [26:0]   _zz_2151;
  wire       [35:0]   _zz_2152;
  wire       [17:0]   _zz_2153;
  wire       [17:0]   _zz_2154;
  wire       [35:0]   _zz_2155;
  wire       [35:0]   _zz_2156;
  wire       [17:0]   _zz_2157;
  wire       [35:0]   _zz_2158;
  wire       [35:0]   _zz_2159;
  wire       [35:0]   _zz_2160;
  wire       [17:0]   _zz_2161;
  wire       [35:0]   _zz_2162;
  wire       [35:0]   _zz_2163;
  wire       [35:0]   _zz_2164;
  wire       [35:0]   _zz_2165;
  wire       [35:0]   _zz_2166;
  wire       [35:0]   _zz_2167;
  wire       [26:0]   _zz_2168;
  wire       [35:0]   _zz_2169;
  wire       [17:0]   _zz_2170;
  wire       [35:0]   _zz_2171;
  wire       [35:0]   _zz_2172;
  wire       [35:0]   _zz_2173;
  wire       [35:0]   _zz_2174;
  wire       [35:0]   _zz_2175;
  wire       [26:0]   _zz_2176;
  wire       [35:0]   _zz_2177;
  wire       [17:0]   _zz_2178;
  wire       [35:0]   _zz_2179;
  wire       [35:0]   _zz_2180;
  wire       [35:0]   _zz_2181;
  wire       [35:0]   _zz_2182;
  wire       [35:0]   _zz_2183;
  wire       [26:0]   _zz_2184;
  wire       [35:0]   _zz_2185;
  wire       [17:0]   _zz_2186;
  wire       [35:0]   _zz_2187;
  wire       [35:0]   _zz_2188;
  wire       [35:0]   _zz_2189;
  wire       [35:0]   _zz_2190;
  wire       [35:0]   _zz_2191;
  wire       [26:0]   _zz_2192;
  wire       [35:0]   _zz_2193;
  wire       [17:0]   _zz_2194;
  wire       [17:0]   _zz_2195;
  wire       [35:0]   _zz_2196;
  wire       [35:0]   _zz_2197;
  wire       [17:0]   _zz_2198;
  wire       [35:0]   _zz_2199;
  wire       [35:0]   _zz_2200;
  wire       [35:0]   _zz_2201;
  wire       [17:0]   _zz_2202;
  wire       [35:0]   _zz_2203;
  wire       [35:0]   _zz_2204;
  wire       [35:0]   _zz_2205;
  wire       [35:0]   _zz_2206;
  wire       [35:0]   _zz_2207;
  wire       [35:0]   _zz_2208;
  wire       [26:0]   _zz_2209;
  wire       [35:0]   _zz_2210;
  wire       [17:0]   _zz_2211;
  wire       [35:0]   _zz_2212;
  wire       [35:0]   _zz_2213;
  wire       [35:0]   _zz_2214;
  wire       [35:0]   _zz_2215;
  wire       [35:0]   _zz_2216;
  wire       [26:0]   _zz_2217;
  wire       [35:0]   _zz_2218;
  wire       [17:0]   _zz_2219;
  wire       [35:0]   _zz_2220;
  wire       [35:0]   _zz_2221;
  wire       [35:0]   _zz_2222;
  wire       [35:0]   _zz_2223;
  wire       [35:0]   _zz_2224;
  wire       [26:0]   _zz_2225;
  wire       [35:0]   _zz_2226;
  wire       [17:0]   _zz_2227;
  wire       [35:0]   _zz_2228;
  wire       [35:0]   _zz_2229;
  wire       [35:0]   _zz_2230;
  wire       [35:0]   _zz_2231;
  wire       [35:0]   _zz_2232;
  wire       [26:0]   _zz_2233;
  wire       [35:0]   _zz_2234;
  wire       [17:0]   _zz_2235;
  wire       [17:0]   _zz_2236;
  wire       [35:0]   _zz_2237;
  wire       [35:0]   _zz_2238;
  wire       [17:0]   _zz_2239;
  wire       [35:0]   _zz_2240;
  wire       [35:0]   _zz_2241;
  wire       [35:0]   _zz_2242;
  wire       [17:0]   _zz_2243;
  wire       [35:0]   _zz_2244;
  wire       [35:0]   _zz_2245;
  wire       [35:0]   _zz_2246;
  wire       [35:0]   _zz_2247;
  wire       [35:0]   _zz_2248;
  wire       [35:0]   _zz_2249;
  wire       [26:0]   _zz_2250;
  wire       [35:0]   _zz_2251;
  wire       [17:0]   _zz_2252;
  wire       [35:0]   _zz_2253;
  wire       [35:0]   _zz_2254;
  wire       [35:0]   _zz_2255;
  wire       [35:0]   _zz_2256;
  wire       [35:0]   _zz_2257;
  wire       [26:0]   _zz_2258;
  wire       [35:0]   _zz_2259;
  wire       [17:0]   _zz_2260;
  wire       [35:0]   _zz_2261;
  wire       [35:0]   _zz_2262;
  wire       [35:0]   _zz_2263;
  wire       [35:0]   _zz_2264;
  wire       [35:0]   _zz_2265;
  wire       [26:0]   _zz_2266;
  wire       [35:0]   _zz_2267;
  wire       [17:0]   _zz_2268;
  wire       [35:0]   _zz_2269;
  wire       [35:0]   _zz_2270;
  wire       [35:0]   _zz_2271;
  wire       [35:0]   _zz_2272;
  wire       [35:0]   _zz_2273;
  wire       [26:0]   _zz_2274;
  wire       [35:0]   _zz_2275;
  wire       [17:0]   _zz_2276;
  wire       [17:0]   _zz_2277;
  wire       [35:0]   _zz_2278;
  wire       [35:0]   _zz_2279;
  wire       [17:0]   _zz_2280;
  wire       [35:0]   _zz_2281;
  wire       [35:0]   _zz_2282;
  wire       [35:0]   _zz_2283;
  wire       [17:0]   _zz_2284;
  wire       [35:0]   _zz_2285;
  wire       [35:0]   _zz_2286;
  wire       [35:0]   _zz_2287;
  wire       [35:0]   _zz_2288;
  wire       [35:0]   _zz_2289;
  wire       [35:0]   _zz_2290;
  wire       [26:0]   _zz_2291;
  wire       [35:0]   _zz_2292;
  wire       [17:0]   _zz_2293;
  wire       [35:0]   _zz_2294;
  wire       [35:0]   _zz_2295;
  wire       [35:0]   _zz_2296;
  wire       [35:0]   _zz_2297;
  wire       [35:0]   _zz_2298;
  wire       [26:0]   _zz_2299;
  wire       [35:0]   _zz_2300;
  wire       [17:0]   _zz_2301;
  wire       [35:0]   _zz_2302;
  wire       [35:0]   _zz_2303;
  wire       [35:0]   _zz_2304;
  wire       [35:0]   _zz_2305;
  wire       [35:0]   _zz_2306;
  wire       [26:0]   _zz_2307;
  wire       [35:0]   _zz_2308;
  wire       [17:0]   _zz_2309;
  wire       [35:0]   _zz_2310;
  wire       [35:0]   _zz_2311;
  wire       [35:0]   _zz_2312;
  wire       [35:0]   _zz_2313;
  wire       [35:0]   _zz_2314;
  wire       [26:0]   _zz_2315;
  wire       [35:0]   _zz_2316;
  wire       [17:0]   _zz_2317;
  wire       [17:0]   _zz_2318;
  wire       [35:0]   _zz_2319;
  wire       [35:0]   _zz_2320;
  wire       [17:0]   _zz_2321;
  wire       [35:0]   _zz_2322;
  wire       [35:0]   _zz_2323;
  wire       [35:0]   _zz_2324;
  wire       [17:0]   _zz_2325;
  wire       [35:0]   _zz_2326;
  wire       [35:0]   _zz_2327;
  wire       [35:0]   _zz_2328;
  wire       [35:0]   _zz_2329;
  wire       [35:0]   _zz_2330;
  wire       [35:0]   _zz_2331;
  wire       [26:0]   _zz_2332;
  wire       [35:0]   _zz_2333;
  wire       [17:0]   _zz_2334;
  wire       [35:0]   _zz_2335;
  wire       [35:0]   _zz_2336;
  wire       [35:0]   _zz_2337;
  wire       [35:0]   _zz_2338;
  wire       [35:0]   _zz_2339;
  wire       [26:0]   _zz_2340;
  wire       [35:0]   _zz_2341;
  wire       [17:0]   _zz_2342;
  wire       [35:0]   _zz_2343;
  wire       [35:0]   _zz_2344;
  wire       [35:0]   _zz_2345;
  wire       [35:0]   _zz_2346;
  wire       [35:0]   _zz_2347;
  wire       [26:0]   _zz_2348;
  wire       [35:0]   _zz_2349;
  wire       [17:0]   _zz_2350;
  wire       [35:0]   _zz_2351;
  wire       [35:0]   _zz_2352;
  wire       [35:0]   _zz_2353;
  wire       [35:0]   _zz_2354;
  wire       [35:0]   _zz_2355;
  wire       [26:0]   _zz_2356;
  wire       [35:0]   _zz_2357;
  wire       [17:0]   _zz_2358;
  wire       [17:0]   _zz_2359;
  wire       [35:0]   _zz_2360;
  wire       [35:0]   _zz_2361;
  wire       [17:0]   _zz_2362;
  wire       [35:0]   _zz_2363;
  wire       [35:0]   _zz_2364;
  wire       [35:0]   _zz_2365;
  wire       [17:0]   _zz_2366;
  wire       [35:0]   _zz_2367;
  wire       [35:0]   _zz_2368;
  wire       [35:0]   _zz_2369;
  wire       [35:0]   _zz_2370;
  wire       [35:0]   _zz_2371;
  wire       [35:0]   _zz_2372;
  wire       [26:0]   _zz_2373;
  wire       [35:0]   _zz_2374;
  wire       [17:0]   _zz_2375;
  wire       [35:0]   _zz_2376;
  wire       [35:0]   _zz_2377;
  wire       [35:0]   _zz_2378;
  wire       [35:0]   _zz_2379;
  wire       [35:0]   _zz_2380;
  wire       [26:0]   _zz_2381;
  wire       [35:0]   _zz_2382;
  wire       [17:0]   _zz_2383;
  wire       [35:0]   _zz_2384;
  wire       [35:0]   _zz_2385;
  wire       [35:0]   _zz_2386;
  wire       [35:0]   _zz_2387;
  wire       [35:0]   _zz_2388;
  wire       [26:0]   _zz_2389;
  wire       [35:0]   _zz_2390;
  wire       [17:0]   _zz_2391;
  wire       [35:0]   _zz_2392;
  wire       [35:0]   _zz_2393;
  wire       [35:0]   _zz_2394;
  wire       [35:0]   _zz_2395;
  wire       [35:0]   _zz_2396;
  wire       [26:0]   _zz_2397;
  wire       [35:0]   _zz_2398;
  wire       [17:0]   _zz_2399;
  wire       [17:0]   _zz_2400;
  wire       [35:0]   _zz_2401;
  wire       [35:0]   _zz_2402;
  wire       [17:0]   _zz_2403;
  wire       [35:0]   _zz_2404;
  wire       [35:0]   _zz_2405;
  wire       [35:0]   _zz_2406;
  wire       [17:0]   _zz_2407;
  wire       [35:0]   _zz_2408;
  wire       [35:0]   _zz_2409;
  wire       [35:0]   _zz_2410;
  wire       [35:0]   _zz_2411;
  wire       [35:0]   _zz_2412;
  wire       [35:0]   _zz_2413;
  wire       [26:0]   _zz_2414;
  wire       [35:0]   _zz_2415;
  wire       [17:0]   _zz_2416;
  wire       [35:0]   _zz_2417;
  wire       [35:0]   _zz_2418;
  wire       [35:0]   _zz_2419;
  wire       [35:0]   _zz_2420;
  wire       [35:0]   _zz_2421;
  wire       [26:0]   _zz_2422;
  wire       [35:0]   _zz_2423;
  wire       [17:0]   _zz_2424;
  wire       [35:0]   _zz_2425;
  wire       [35:0]   _zz_2426;
  wire       [35:0]   _zz_2427;
  wire       [35:0]   _zz_2428;
  wire       [35:0]   _zz_2429;
  wire       [26:0]   _zz_2430;
  wire       [35:0]   _zz_2431;
  wire       [17:0]   _zz_2432;
  wire       [35:0]   _zz_2433;
  wire       [35:0]   _zz_2434;
  wire       [35:0]   _zz_2435;
  wire       [35:0]   _zz_2436;
  wire       [35:0]   _zz_2437;
  wire       [26:0]   _zz_2438;
  wire       [35:0]   _zz_2439;
  wire       [17:0]   _zz_2440;
  wire       [17:0]   _zz_2441;
  wire       [35:0]   _zz_2442;
  wire       [35:0]   _zz_2443;
  wire       [17:0]   _zz_2444;
  wire       [35:0]   _zz_2445;
  wire       [35:0]   _zz_2446;
  wire       [35:0]   _zz_2447;
  wire       [17:0]   _zz_2448;
  wire       [35:0]   _zz_2449;
  wire       [35:0]   _zz_2450;
  wire       [35:0]   _zz_2451;
  wire       [35:0]   _zz_2452;
  wire       [35:0]   _zz_2453;
  wire       [35:0]   _zz_2454;
  wire       [26:0]   _zz_2455;
  wire       [35:0]   _zz_2456;
  wire       [17:0]   _zz_2457;
  wire       [35:0]   _zz_2458;
  wire       [35:0]   _zz_2459;
  wire       [35:0]   _zz_2460;
  wire       [35:0]   _zz_2461;
  wire       [35:0]   _zz_2462;
  wire       [26:0]   _zz_2463;
  wire       [35:0]   _zz_2464;
  wire       [17:0]   _zz_2465;
  wire       [35:0]   _zz_2466;
  wire       [35:0]   _zz_2467;
  wire       [35:0]   _zz_2468;
  wire       [35:0]   _zz_2469;
  wire       [35:0]   _zz_2470;
  wire       [26:0]   _zz_2471;
  wire       [35:0]   _zz_2472;
  wire       [17:0]   _zz_2473;
  wire       [35:0]   _zz_2474;
  wire       [35:0]   _zz_2475;
  wire       [35:0]   _zz_2476;
  wire       [35:0]   _zz_2477;
  wire       [35:0]   _zz_2478;
  wire       [26:0]   _zz_2479;
  wire       [35:0]   _zz_2480;
  wire       [17:0]   _zz_2481;
  wire       [17:0]   _zz_2482;
  wire       [35:0]   _zz_2483;
  wire       [35:0]   _zz_2484;
  wire       [17:0]   _zz_2485;
  wire       [35:0]   _zz_2486;
  wire       [35:0]   _zz_2487;
  wire       [35:0]   _zz_2488;
  wire       [17:0]   _zz_2489;
  wire       [35:0]   _zz_2490;
  wire       [35:0]   _zz_2491;
  wire       [35:0]   _zz_2492;
  wire       [35:0]   _zz_2493;
  wire       [35:0]   _zz_2494;
  wire       [35:0]   _zz_2495;
  wire       [26:0]   _zz_2496;
  wire       [35:0]   _zz_2497;
  wire       [17:0]   _zz_2498;
  wire       [35:0]   _zz_2499;
  wire       [35:0]   _zz_2500;
  wire       [35:0]   _zz_2501;
  wire       [35:0]   _zz_2502;
  wire       [35:0]   _zz_2503;
  wire       [26:0]   _zz_2504;
  wire       [35:0]   _zz_2505;
  wire       [17:0]   _zz_2506;
  wire       [35:0]   _zz_2507;
  wire       [35:0]   _zz_2508;
  wire       [35:0]   _zz_2509;
  wire       [35:0]   _zz_2510;
  wire       [35:0]   _zz_2511;
  wire       [26:0]   _zz_2512;
  wire       [35:0]   _zz_2513;
  wire       [17:0]   _zz_2514;
  wire       [35:0]   _zz_2515;
  wire       [35:0]   _zz_2516;
  wire       [35:0]   _zz_2517;
  wire       [35:0]   _zz_2518;
  wire       [35:0]   _zz_2519;
  wire       [26:0]   _zz_2520;
  wire       [35:0]   _zz_2521;
  wire       [17:0]   _zz_2522;
  wire       [17:0]   _zz_2523;
  wire       [35:0]   _zz_2524;
  wire       [35:0]   _zz_2525;
  wire       [17:0]   _zz_2526;
  wire       [35:0]   _zz_2527;
  wire       [35:0]   _zz_2528;
  wire       [35:0]   _zz_2529;
  wire       [17:0]   _zz_2530;
  wire       [35:0]   _zz_2531;
  wire       [35:0]   _zz_2532;
  wire       [35:0]   _zz_2533;
  wire       [35:0]   _zz_2534;
  wire       [35:0]   _zz_2535;
  wire       [35:0]   _zz_2536;
  wire       [26:0]   _zz_2537;
  wire       [35:0]   _zz_2538;
  wire       [17:0]   _zz_2539;
  wire       [35:0]   _zz_2540;
  wire       [35:0]   _zz_2541;
  wire       [35:0]   _zz_2542;
  wire       [35:0]   _zz_2543;
  wire       [35:0]   _zz_2544;
  wire       [26:0]   _zz_2545;
  wire       [35:0]   _zz_2546;
  wire       [17:0]   _zz_2547;
  wire       [35:0]   _zz_2548;
  wire       [35:0]   _zz_2549;
  wire       [35:0]   _zz_2550;
  wire       [35:0]   _zz_2551;
  wire       [35:0]   _zz_2552;
  wire       [26:0]   _zz_2553;
  wire       [35:0]   _zz_2554;
  wire       [17:0]   _zz_2555;
  wire       [35:0]   _zz_2556;
  wire       [35:0]   _zz_2557;
  wire       [35:0]   _zz_2558;
  wire       [35:0]   _zz_2559;
  wire       [35:0]   _zz_2560;
  wire       [26:0]   _zz_2561;
  wire       [35:0]   _zz_2562;
  wire       [17:0]   _zz_2563;
  wire       [17:0]   _zz_2564;
  wire       [35:0]   _zz_2565;
  wire       [35:0]   _zz_2566;
  wire       [17:0]   _zz_2567;
  wire       [35:0]   _zz_2568;
  wire       [35:0]   _zz_2569;
  wire       [35:0]   _zz_2570;
  wire       [17:0]   _zz_2571;
  wire       [35:0]   _zz_2572;
  wire       [35:0]   _zz_2573;
  wire       [35:0]   _zz_2574;
  wire       [35:0]   _zz_2575;
  wire       [35:0]   _zz_2576;
  wire       [35:0]   _zz_2577;
  wire       [26:0]   _zz_2578;
  wire       [35:0]   _zz_2579;
  wire       [17:0]   _zz_2580;
  wire       [35:0]   _zz_2581;
  wire       [35:0]   _zz_2582;
  wire       [35:0]   _zz_2583;
  wire       [35:0]   _zz_2584;
  wire       [35:0]   _zz_2585;
  wire       [26:0]   _zz_2586;
  wire       [35:0]   _zz_2587;
  wire       [17:0]   _zz_2588;
  wire       [35:0]   _zz_2589;
  wire       [35:0]   _zz_2590;
  wire       [35:0]   _zz_2591;
  wire       [35:0]   _zz_2592;
  wire       [35:0]   _zz_2593;
  wire       [26:0]   _zz_2594;
  wire       [35:0]   _zz_2595;
  wire       [17:0]   _zz_2596;
  wire       [35:0]   _zz_2597;
  wire       [35:0]   _zz_2598;
  wire       [35:0]   _zz_2599;
  wire       [35:0]   _zz_2600;
  wire       [35:0]   _zz_2601;
  wire       [26:0]   _zz_2602;
  wire       [35:0]   _zz_2603;
  wire       [17:0]   _zz_2604;
  wire       [17:0]   _zz_2605;
  wire       [35:0]   _zz_2606;
  wire       [35:0]   _zz_2607;
  wire       [17:0]   _zz_2608;
  wire       [35:0]   _zz_2609;
  wire       [35:0]   _zz_2610;
  wire       [35:0]   _zz_2611;
  wire       [17:0]   _zz_2612;
  wire       [35:0]   _zz_2613;
  wire       [35:0]   _zz_2614;
  wire       [35:0]   _zz_2615;
  wire       [35:0]   _zz_2616;
  wire       [35:0]   _zz_2617;
  wire       [35:0]   _zz_2618;
  wire       [26:0]   _zz_2619;
  wire       [35:0]   _zz_2620;
  wire       [17:0]   _zz_2621;
  wire       [35:0]   _zz_2622;
  wire       [35:0]   _zz_2623;
  wire       [35:0]   _zz_2624;
  wire       [35:0]   _zz_2625;
  wire       [35:0]   _zz_2626;
  wire       [26:0]   _zz_2627;
  wire       [35:0]   _zz_2628;
  wire       [17:0]   _zz_2629;
  wire       [35:0]   _zz_2630;
  wire       [35:0]   _zz_2631;
  wire       [35:0]   _zz_2632;
  wire       [35:0]   _zz_2633;
  wire       [35:0]   _zz_2634;
  wire       [26:0]   _zz_2635;
  wire       [35:0]   _zz_2636;
  wire       [17:0]   _zz_2637;
  wire       [35:0]   _zz_2638;
  wire       [35:0]   _zz_2639;
  wire       [35:0]   _zz_2640;
  wire       [35:0]   _zz_2641;
  wire       [35:0]   _zz_2642;
  wire       [26:0]   _zz_2643;
  wire       [35:0]   _zz_2644;
  wire       [17:0]   _zz_2645;
  wire       [17:0]   _zz_2646;
  wire       [35:0]   _zz_2647;
  wire       [35:0]   _zz_2648;
  wire       [17:0]   _zz_2649;
  wire       [35:0]   _zz_2650;
  wire       [35:0]   _zz_2651;
  wire       [35:0]   _zz_2652;
  wire       [17:0]   _zz_2653;
  wire       [35:0]   _zz_2654;
  wire       [35:0]   _zz_2655;
  wire       [35:0]   _zz_2656;
  wire       [35:0]   _zz_2657;
  wire       [35:0]   _zz_2658;
  wire       [35:0]   _zz_2659;
  wire       [26:0]   _zz_2660;
  wire       [35:0]   _zz_2661;
  wire       [17:0]   _zz_2662;
  wire       [35:0]   _zz_2663;
  wire       [35:0]   _zz_2664;
  wire       [35:0]   _zz_2665;
  wire       [35:0]   _zz_2666;
  wire       [35:0]   _zz_2667;
  wire       [26:0]   _zz_2668;
  wire       [35:0]   _zz_2669;
  wire       [17:0]   _zz_2670;
  wire       [35:0]   _zz_2671;
  wire       [35:0]   _zz_2672;
  wire       [35:0]   _zz_2673;
  wire       [35:0]   _zz_2674;
  wire       [35:0]   _zz_2675;
  wire       [26:0]   _zz_2676;
  wire       [35:0]   _zz_2677;
  wire       [17:0]   _zz_2678;
  wire       [35:0]   _zz_2679;
  wire       [35:0]   _zz_2680;
  wire       [35:0]   _zz_2681;
  wire       [35:0]   _zz_2682;
  wire       [35:0]   _zz_2683;
  wire       [26:0]   _zz_2684;
  wire       [35:0]   _zz_2685;
  wire       [17:0]   _zz_2686;
  wire       [17:0]   _zz_2687;
  wire       [35:0]   _zz_2688;
  wire       [35:0]   _zz_2689;
  wire       [17:0]   _zz_2690;
  wire       [35:0]   _zz_2691;
  wire       [35:0]   _zz_2692;
  wire       [35:0]   _zz_2693;
  wire       [17:0]   _zz_2694;
  wire       [35:0]   _zz_2695;
  wire       [35:0]   _zz_2696;
  wire       [35:0]   _zz_2697;
  wire       [35:0]   _zz_2698;
  wire       [35:0]   _zz_2699;
  wire       [35:0]   _zz_2700;
  wire       [26:0]   _zz_2701;
  wire       [35:0]   _zz_2702;
  wire       [17:0]   _zz_2703;
  wire       [35:0]   _zz_2704;
  wire       [35:0]   _zz_2705;
  wire       [35:0]   _zz_2706;
  wire       [35:0]   _zz_2707;
  wire       [35:0]   _zz_2708;
  wire       [26:0]   _zz_2709;
  wire       [35:0]   _zz_2710;
  wire       [17:0]   _zz_2711;
  wire       [35:0]   _zz_2712;
  wire       [35:0]   _zz_2713;
  wire       [35:0]   _zz_2714;
  wire       [35:0]   _zz_2715;
  wire       [35:0]   _zz_2716;
  wire       [26:0]   _zz_2717;
  wire       [35:0]   _zz_2718;
  wire       [17:0]   _zz_2719;
  wire       [35:0]   _zz_2720;
  wire       [35:0]   _zz_2721;
  wire       [35:0]   _zz_2722;
  wire       [35:0]   _zz_2723;
  wire       [35:0]   _zz_2724;
  wire       [26:0]   _zz_2725;
  wire       [35:0]   _zz_2726;
  wire       [17:0]   _zz_2727;
  wire       [17:0]   _zz_2728;
  wire       [35:0]   _zz_2729;
  wire       [35:0]   _zz_2730;
  wire       [17:0]   _zz_2731;
  wire       [35:0]   _zz_2732;
  wire       [35:0]   _zz_2733;
  wire       [35:0]   _zz_2734;
  wire       [17:0]   _zz_2735;
  wire       [35:0]   _zz_2736;
  wire       [35:0]   _zz_2737;
  wire       [35:0]   _zz_2738;
  wire       [35:0]   _zz_2739;
  wire       [35:0]   _zz_2740;
  wire       [35:0]   _zz_2741;
  wire       [26:0]   _zz_2742;
  wire       [35:0]   _zz_2743;
  wire       [17:0]   _zz_2744;
  wire       [35:0]   _zz_2745;
  wire       [35:0]   _zz_2746;
  wire       [35:0]   _zz_2747;
  wire       [35:0]   _zz_2748;
  wire       [35:0]   _zz_2749;
  wire       [26:0]   _zz_2750;
  wire       [35:0]   _zz_2751;
  wire       [17:0]   _zz_2752;
  wire       [35:0]   _zz_2753;
  wire       [35:0]   _zz_2754;
  wire       [35:0]   _zz_2755;
  wire       [35:0]   _zz_2756;
  wire       [35:0]   _zz_2757;
  wire       [26:0]   _zz_2758;
  wire       [35:0]   _zz_2759;
  wire       [17:0]   _zz_2760;
  wire       [35:0]   _zz_2761;
  wire       [35:0]   _zz_2762;
  wire       [35:0]   _zz_2763;
  wire       [35:0]   _zz_2764;
  wire       [35:0]   _zz_2765;
  wire       [26:0]   _zz_2766;
  wire       [35:0]   _zz_2767;
  wire       [17:0]   _zz_2768;
  wire       [17:0]   _zz_2769;
  wire       [35:0]   _zz_2770;
  wire       [35:0]   _zz_2771;
  wire       [17:0]   _zz_2772;
  wire       [35:0]   _zz_2773;
  wire       [35:0]   _zz_2774;
  wire       [35:0]   _zz_2775;
  wire       [17:0]   _zz_2776;
  wire       [35:0]   _zz_2777;
  wire       [35:0]   _zz_2778;
  wire       [35:0]   _zz_2779;
  wire       [35:0]   _zz_2780;
  wire       [35:0]   _zz_2781;
  wire       [35:0]   _zz_2782;
  wire       [26:0]   _zz_2783;
  wire       [35:0]   _zz_2784;
  wire       [17:0]   _zz_2785;
  wire       [35:0]   _zz_2786;
  wire       [35:0]   _zz_2787;
  wire       [35:0]   _zz_2788;
  wire       [35:0]   _zz_2789;
  wire       [35:0]   _zz_2790;
  wire       [26:0]   _zz_2791;
  wire       [35:0]   _zz_2792;
  wire       [17:0]   _zz_2793;
  wire       [35:0]   _zz_2794;
  wire       [35:0]   _zz_2795;
  wire       [35:0]   _zz_2796;
  wire       [35:0]   _zz_2797;
  wire       [35:0]   _zz_2798;
  wire       [26:0]   _zz_2799;
  wire       [35:0]   _zz_2800;
  wire       [17:0]   _zz_2801;
  wire       [35:0]   _zz_2802;
  wire       [35:0]   _zz_2803;
  wire       [35:0]   _zz_2804;
  wire       [35:0]   _zz_2805;
  wire       [35:0]   _zz_2806;
  wire       [26:0]   _zz_2807;
  wire       [35:0]   _zz_2808;
  wire       [17:0]   _zz_2809;
  wire       [17:0]   _zz_2810;
  wire       [35:0]   _zz_2811;
  wire       [35:0]   _zz_2812;
  wire       [17:0]   _zz_2813;
  wire       [35:0]   _zz_2814;
  wire       [35:0]   _zz_2815;
  wire       [35:0]   _zz_2816;
  wire       [17:0]   _zz_2817;
  wire       [35:0]   _zz_2818;
  wire       [35:0]   _zz_2819;
  wire       [35:0]   _zz_2820;
  wire       [35:0]   _zz_2821;
  wire       [35:0]   _zz_2822;
  wire       [35:0]   _zz_2823;
  wire       [26:0]   _zz_2824;
  wire       [35:0]   _zz_2825;
  wire       [17:0]   _zz_2826;
  wire       [35:0]   _zz_2827;
  wire       [35:0]   _zz_2828;
  wire       [35:0]   _zz_2829;
  wire       [35:0]   _zz_2830;
  wire       [35:0]   _zz_2831;
  wire       [26:0]   _zz_2832;
  wire       [35:0]   _zz_2833;
  wire       [17:0]   _zz_2834;
  wire       [35:0]   _zz_2835;
  wire       [35:0]   _zz_2836;
  wire       [35:0]   _zz_2837;
  wire       [35:0]   _zz_2838;
  wire       [35:0]   _zz_2839;
  wire       [26:0]   _zz_2840;
  wire       [35:0]   _zz_2841;
  wire       [17:0]   _zz_2842;
  wire       [35:0]   _zz_2843;
  wire       [35:0]   _zz_2844;
  wire       [35:0]   _zz_2845;
  wire       [35:0]   _zz_2846;
  wire       [35:0]   _zz_2847;
  wire       [26:0]   _zz_2848;
  wire       [35:0]   _zz_2849;
  wire       [17:0]   _zz_2850;
  wire       [17:0]   _zz_2851;
  wire       [35:0]   _zz_2852;
  wire       [35:0]   _zz_2853;
  wire       [17:0]   _zz_2854;
  wire       [35:0]   _zz_2855;
  wire       [35:0]   _zz_2856;
  wire       [35:0]   _zz_2857;
  wire       [17:0]   _zz_2858;
  wire       [35:0]   _zz_2859;
  wire       [35:0]   _zz_2860;
  wire       [35:0]   _zz_2861;
  wire       [35:0]   _zz_2862;
  wire       [35:0]   _zz_2863;
  wire       [35:0]   _zz_2864;
  wire       [26:0]   _zz_2865;
  wire       [35:0]   _zz_2866;
  wire       [17:0]   _zz_2867;
  wire       [35:0]   _zz_2868;
  wire       [35:0]   _zz_2869;
  wire       [35:0]   _zz_2870;
  wire       [35:0]   _zz_2871;
  wire       [35:0]   _zz_2872;
  wire       [26:0]   _zz_2873;
  wire       [35:0]   _zz_2874;
  wire       [17:0]   _zz_2875;
  wire       [35:0]   _zz_2876;
  wire       [35:0]   _zz_2877;
  wire       [35:0]   _zz_2878;
  wire       [35:0]   _zz_2879;
  wire       [35:0]   _zz_2880;
  wire       [26:0]   _zz_2881;
  wire       [35:0]   _zz_2882;
  wire       [17:0]   _zz_2883;
  wire       [35:0]   _zz_2884;
  wire       [35:0]   _zz_2885;
  wire       [35:0]   _zz_2886;
  wire       [35:0]   _zz_2887;
  wire       [35:0]   _zz_2888;
  wire       [26:0]   _zz_2889;
  wire       [35:0]   _zz_2890;
  wire       [17:0]   _zz_2891;
  wire       [17:0]   _zz_2892;
  wire       [35:0]   _zz_2893;
  wire       [35:0]   _zz_2894;
  wire       [17:0]   _zz_2895;
  wire       [35:0]   _zz_2896;
  wire       [35:0]   _zz_2897;
  wire       [35:0]   _zz_2898;
  wire       [17:0]   _zz_2899;
  wire       [35:0]   _zz_2900;
  wire       [35:0]   _zz_2901;
  wire       [35:0]   _zz_2902;
  wire       [35:0]   _zz_2903;
  wire       [35:0]   _zz_2904;
  wire       [35:0]   _zz_2905;
  wire       [26:0]   _zz_2906;
  wire       [35:0]   _zz_2907;
  wire       [17:0]   _zz_2908;
  wire       [35:0]   _zz_2909;
  wire       [35:0]   _zz_2910;
  wire       [35:0]   _zz_2911;
  wire       [35:0]   _zz_2912;
  wire       [35:0]   _zz_2913;
  wire       [26:0]   _zz_2914;
  wire       [35:0]   _zz_2915;
  wire       [17:0]   _zz_2916;
  wire       [35:0]   _zz_2917;
  wire       [35:0]   _zz_2918;
  wire       [35:0]   _zz_2919;
  wire       [35:0]   _zz_2920;
  wire       [35:0]   _zz_2921;
  wire       [26:0]   _zz_2922;
  wire       [35:0]   _zz_2923;
  wire       [17:0]   _zz_2924;
  wire       [35:0]   _zz_2925;
  wire       [35:0]   _zz_2926;
  wire       [35:0]   _zz_2927;
  wire       [35:0]   _zz_2928;
  wire       [35:0]   _zz_2929;
  wire       [26:0]   _zz_2930;
  wire       [35:0]   _zz_2931;
  wire       [17:0]   _zz_2932;
  wire       [17:0]   _zz_2933;
  wire       [35:0]   _zz_2934;
  wire       [35:0]   _zz_2935;
  wire       [17:0]   _zz_2936;
  wire       [35:0]   _zz_2937;
  wire       [35:0]   _zz_2938;
  wire       [35:0]   _zz_2939;
  wire       [17:0]   _zz_2940;
  wire       [35:0]   _zz_2941;
  wire       [35:0]   _zz_2942;
  wire       [35:0]   _zz_2943;
  wire       [35:0]   _zz_2944;
  wire       [35:0]   _zz_2945;
  wire       [35:0]   _zz_2946;
  wire       [26:0]   _zz_2947;
  wire       [35:0]   _zz_2948;
  wire       [17:0]   _zz_2949;
  wire       [35:0]   _zz_2950;
  wire       [35:0]   _zz_2951;
  wire       [35:0]   _zz_2952;
  wire       [35:0]   _zz_2953;
  wire       [35:0]   _zz_2954;
  wire       [26:0]   _zz_2955;
  wire       [35:0]   _zz_2956;
  wire       [17:0]   _zz_2957;
  wire       [35:0]   _zz_2958;
  wire       [35:0]   _zz_2959;
  wire       [35:0]   _zz_2960;
  wire       [35:0]   _zz_2961;
  wire       [35:0]   _zz_2962;
  wire       [26:0]   _zz_2963;
  wire       [35:0]   _zz_2964;
  wire       [17:0]   _zz_2965;
  wire       [35:0]   _zz_2966;
  wire       [35:0]   _zz_2967;
  wire       [35:0]   _zz_2968;
  wire       [35:0]   _zz_2969;
  wire       [35:0]   _zz_2970;
  wire       [26:0]   _zz_2971;
  wire       [35:0]   _zz_2972;
  wire       [17:0]   _zz_2973;
  wire       [17:0]   _zz_2974;
  wire       [35:0]   _zz_2975;
  wire       [35:0]   _zz_2976;
  wire       [17:0]   _zz_2977;
  wire       [35:0]   _zz_2978;
  wire       [35:0]   _zz_2979;
  wire       [35:0]   _zz_2980;
  wire       [17:0]   _zz_2981;
  wire       [35:0]   _zz_2982;
  wire       [35:0]   _zz_2983;
  wire       [35:0]   _zz_2984;
  wire       [35:0]   _zz_2985;
  wire       [35:0]   _zz_2986;
  wire       [35:0]   _zz_2987;
  wire       [26:0]   _zz_2988;
  wire       [35:0]   _zz_2989;
  wire       [17:0]   _zz_2990;
  wire       [35:0]   _zz_2991;
  wire       [35:0]   _zz_2992;
  wire       [35:0]   _zz_2993;
  wire       [35:0]   _zz_2994;
  wire       [35:0]   _zz_2995;
  wire       [26:0]   _zz_2996;
  wire       [35:0]   _zz_2997;
  wire       [17:0]   _zz_2998;
  wire       [35:0]   _zz_2999;
  wire       [35:0]   _zz_3000;
  wire       [35:0]   _zz_3001;
  wire       [35:0]   _zz_3002;
  wire       [35:0]   _zz_3003;
  wire       [26:0]   _zz_3004;
  wire       [35:0]   _zz_3005;
  wire       [17:0]   _zz_3006;
  wire       [35:0]   _zz_3007;
  wire       [35:0]   _zz_3008;
  wire       [35:0]   _zz_3009;
  wire       [35:0]   _zz_3010;
  wire       [35:0]   _zz_3011;
  wire       [26:0]   _zz_3012;
  wire       [35:0]   _zz_3013;
  wire       [17:0]   _zz_3014;
  wire       [17:0]   _zz_3015;
  wire       [35:0]   _zz_3016;
  wire       [35:0]   _zz_3017;
  wire       [17:0]   _zz_3018;
  wire       [35:0]   _zz_3019;
  wire       [35:0]   _zz_3020;
  wire       [35:0]   _zz_3021;
  wire       [17:0]   _zz_3022;
  wire       [35:0]   _zz_3023;
  wire       [35:0]   _zz_3024;
  wire       [35:0]   _zz_3025;
  wire       [35:0]   _zz_3026;
  wire       [35:0]   _zz_3027;
  wire       [35:0]   _zz_3028;
  wire       [26:0]   _zz_3029;
  wire       [35:0]   _zz_3030;
  wire       [17:0]   _zz_3031;
  wire       [35:0]   _zz_3032;
  wire       [35:0]   _zz_3033;
  wire       [35:0]   _zz_3034;
  wire       [35:0]   _zz_3035;
  wire       [35:0]   _zz_3036;
  wire       [26:0]   _zz_3037;
  wire       [35:0]   _zz_3038;
  wire       [17:0]   _zz_3039;
  wire       [35:0]   _zz_3040;
  wire       [35:0]   _zz_3041;
  wire       [35:0]   _zz_3042;
  wire       [35:0]   _zz_3043;
  wire       [35:0]   _zz_3044;
  wire       [26:0]   _zz_3045;
  wire       [35:0]   _zz_3046;
  wire       [17:0]   _zz_3047;
  wire       [35:0]   _zz_3048;
  wire       [35:0]   _zz_3049;
  wire       [35:0]   _zz_3050;
  wire       [35:0]   _zz_3051;
  wire       [35:0]   _zz_3052;
  wire       [26:0]   _zz_3053;
  wire       [35:0]   _zz_3054;
  wire       [17:0]   _zz_3055;
  wire       [17:0]   _zz_3056;
  wire       [35:0]   _zz_3057;
  wire       [35:0]   _zz_3058;
  wire       [17:0]   _zz_3059;
  wire       [35:0]   _zz_3060;
  wire       [35:0]   _zz_3061;
  wire       [35:0]   _zz_3062;
  wire       [17:0]   _zz_3063;
  wire       [35:0]   _zz_3064;
  wire       [35:0]   _zz_3065;
  wire       [35:0]   _zz_3066;
  wire       [35:0]   _zz_3067;
  wire       [35:0]   _zz_3068;
  wire       [35:0]   _zz_3069;
  wire       [26:0]   _zz_3070;
  wire       [35:0]   _zz_3071;
  wire       [17:0]   _zz_3072;
  wire       [35:0]   _zz_3073;
  wire       [35:0]   _zz_3074;
  wire       [35:0]   _zz_3075;
  wire       [35:0]   _zz_3076;
  wire       [35:0]   _zz_3077;
  wire       [26:0]   _zz_3078;
  wire       [35:0]   _zz_3079;
  wire       [17:0]   _zz_3080;
  wire       [35:0]   _zz_3081;
  wire       [35:0]   _zz_3082;
  wire       [35:0]   _zz_3083;
  wire       [35:0]   _zz_3084;
  wire       [35:0]   _zz_3085;
  wire       [26:0]   _zz_3086;
  wire       [35:0]   _zz_3087;
  wire       [17:0]   _zz_3088;
  wire       [35:0]   _zz_3089;
  wire       [35:0]   _zz_3090;
  wire       [35:0]   _zz_3091;
  wire       [35:0]   _zz_3092;
  wire       [35:0]   _zz_3093;
  wire       [26:0]   _zz_3094;
  wire       [35:0]   _zz_3095;
  wire       [17:0]   _zz_3096;
  wire       [17:0]   _zz_3097;
  wire       [35:0]   _zz_3098;
  wire       [35:0]   _zz_3099;
  wire       [17:0]   _zz_3100;
  wire       [35:0]   _zz_3101;
  wire       [35:0]   _zz_3102;
  wire       [35:0]   _zz_3103;
  wire       [17:0]   _zz_3104;
  wire       [35:0]   _zz_3105;
  wire       [35:0]   _zz_3106;
  wire       [35:0]   _zz_3107;
  wire       [35:0]   _zz_3108;
  wire       [35:0]   _zz_3109;
  wire       [35:0]   _zz_3110;
  wire       [26:0]   _zz_3111;
  wire       [35:0]   _zz_3112;
  wire       [17:0]   _zz_3113;
  wire       [35:0]   _zz_3114;
  wire       [35:0]   _zz_3115;
  wire       [35:0]   _zz_3116;
  wire       [35:0]   _zz_3117;
  wire       [35:0]   _zz_3118;
  wire       [26:0]   _zz_3119;
  wire       [35:0]   _zz_3120;
  wire       [17:0]   _zz_3121;
  wire       [35:0]   _zz_3122;
  wire       [35:0]   _zz_3123;
  wire       [35:0]   _zz_3124;
  wire       [35:0]   _zz_3125;
  wire       [35:0]   _zz_3126;
  wire       [26:0]   _zz_3127;
  wire       [35:0]   _zz_3128;
  wire       [17:0]   _zz_3129;
  wire       [35:0]   _zz_3130;
  wire       [35:0]   _zz_3131;
  wire       [35:0]   _zz_3132;
  wire       [35:0]   _zz_3133;
  wire       [35:0]   _zz_3134;
  wire       [26:0]   _zz_3135;
  wire       [35:0]   _zz_3136;
  wire       [17:0]   _zz_3137;
  wire       [17:0]   _zz_3138;
  wire       [35:0]   _zz_3139;
  wire       [35:0]   _zz_3140;
  wire       [17:0]   _zz_3141;
  wire       [35:0]   _zz_3142;
  wire       [35:0]   _zz_3143;
  wire       [35:0]   _zz_3144;
  wire       [17:0]   _zz_3145;
  wire       [35:0]   _zz_3146;
  wire       [35:0]   _zz_3147;
  wire       [35:0]   _zz_3148;
  wire       [35:0]   _zz_3149;
  wire       [35:0]   _zz_3150;
  wire       [35:0]   _zz_3151;
  wire       [26:0]   _zz_3152;
  wire       [35:0]   _zz_3153;
  wire       [17:0]   _zz_3154;
  wire       [35:0]   _zz_3155;
  wire       [35:0]   _zz_3156;
  wire       [35:0]   _zz_3157;
  wire       [35:0]   _zz_3158;
  wire       [35:0]   _zz_3159;
  wire       [26:0]   _zz_3160;
  wire       [35:0]   _zz_3161;
  wire       [17:0]   _zz_3162;
  wire       [35:0]   _zz_3163;
  wire       [35:0]   _zz_3164;
  wire       [35:0]   _zz_3165;
  wire       [35:0]   _zz_3166;
  wire       [35:0]   _zz_3167;
  wire       [26:0]   _zz_3168;
  wire       [35:0]   _zz_3169;
  wire       [17:0]   _zz_3170;
  wire       [35:0]   _zz_3171;
  wire       [35:0]   _zz_3172;
  wire       [35:0]   _zz_3173;
  wire       [35:0]   _zz_3174;
  wire       [35:0]   _zz_3175;
  wire       [26:0]   _zz_3176;
  wire       [35:0]   _zz_3177;
  wire       [17:0]   _zz_3178;
  wire       [17:0]   _zz_3179;
  wire       [35:0]   _zz_3180;
  wire       [35:0]   _zz_3181;
  wire       [17:0]   _zz_3182;
  wire       [35:0]   _zz_3183;
  wire       [35:0]   _zz_3184;
  wire       [35:0]   _zz_3185;
  wire       [17:0]   _zz_3186;
  wire       [35:0]   _zz_3187;
  wire       [35:0]   _zz_3188;
  wire       [35:0]   _zz_3189;
  wire       [35:0]   _zz_3190;
  wire       [35:0]   _zz_3191;
  wire       [35:0]   _zz_3192;
  wire       [26:0]   _zz_3193;
  wire       [35:0]   _zz_3194;
  wire       [17:0]   _zz_3195;
  wire       [35:0]   _zz_3196;
  wire       [35:0]   _zz_3197;
  wire       [35:0]   _zz_3198;
  wire       [35:0]   _zz_3199;
  wire       [35:0]   _zz_3200;
  wire       [26:0]   _zz_3201;
  wire       [35:0]   _zz_3202;
  wire       [17:0]   _zz_3203;
  wire       [35:0]   _zz_3204;
  wire       [35:0]   _zz_3205;
  wire       [35:0]   _zz_3206;
  wire       [35:0]   _zz_3207;
  wire       [35:0]   _zz_3208;
  wire       [26:0]   _zz_3209;
  wire       [35:0]   _zz_3210;
  wire       [17:0]   _zz_3211;
  wire       [35:0]   _zz_3212;
  wire       [35:0]   _zz_3213;
  wire       [35:0]   _zz_3214;
  wire       [35:0]   _zz_3215;
  wire       [35:0]   _zz_3216;
  wire       [26:0]   _zz_3217;
  wire       [35:0]   _zz_3218;
  wire       [17:0]   _zz_3219;
  wire       [17:0]   _zz_3220;
  wire       [35:0]   _zz_3221;
  wire       [35:0]   _zz_3222;
  wire       [17:0]   _zz_3223;
  wire       [35:0]   _zz_3224;
  wire       [35:0]   _zz_3225;
  wire       [35:0]   _zz_3226;
  wire       [17:0]   _zz_3227;
  wire       [35:0]   _zz_3228;
  wire       [35:0]   _zz_3229;
  wire       [35:0]   _zz_3230;
  wire       [35:0]   _zz_3231;
  wire       [35:0]   _zz_3232;
  wire       [35:0]   _zz_3233;
  wire       [26:0]   _zz_3234;
  wire       [35:0]   _zz_3235;
  wire       [17:0]   _zz_3236;
  wire       [35:0]   _zz_3237;
  wire       [35:0]   _zz_3238;
  wire       [35:0]   _zz_3239;
  wire       [35:0]   _zz_3240;
  wire       [35:0]   _zz_3241;
  wire       [26:0]   _zz_3242;
  wire       [35:0]   _zz_3243;
  wire       [17:0]   _zz_3244;
  wire       [35:0]   _zz_3245;
  wire       [35:0]   _zz_3246;
  wire       [35:0]   _zz_3247;
  wire       [35:0]   _zz_3248;
  wire       [35:0]   _zz_3249;
  wire       [26:0]   _zz_3250;
  wire       [35:0]   _zz_3251;
  wire       [17:0]   _zz_3252;
  wire       [35:0]   _zz_3253;
  wire       [35:0]   _zz_3254;
  wire       [35:0]   _zz_3255;
  wire       [35:0]   _zz_3256;
  wire       [35:0]   _zz_3257;
  wire       [26:0]   _zz_3258;
  wire       [35:0]   _zz_3259;
  wire       [17:0]   _zz_3260;
  wire       [17:0]   _zz_3261;
  wire       [35:0]   _zz_3262;
  wire       [35:0]   _zz_3263;
  wire       [17:0]   _zz_3264;
  wire       [35:0]   _zz_3265;
  wire       [35:0]   _zz_3266;
  wire       [35:0]   _zz_3267;
  wire       [17:0]   _zz_3268;
  wire       [35:0]   _zz_3269;
  wire       [35:0]   _zz_3270;
  wire       [35:0]   _zz_3271;
  wire       [35:0]   _zz_3272;
  wire       [35:0]   _zz_3273;
  wire       [35:0]   _zz_3274;
  wire       [26:0]   _zz_3275;
  wire       [35:0]   _zz_3276;
  wire       [17:0]   _zz_3277;
  wire       [35:0]   _zz_3278;
  wire       [35:0]   _zz_3279;
  wire       [35:0]   _zz_3280;
  wire       [35:0]   _zz_3281;
  wire       [35:0]   _zz_3282;
  wire       [26:0]   _zz_3283;
  wire       [35:0]   _zz_3284;
  wire       [17:0]   _zz_3285;
  wire       [35:0]   _zz_3286;
  wire       [35:0]   _zz_3287;
  wire       [35:0]   _zz_3288;
  wire       [35:0]   _zz_3289;
  wire       [35:0]   _zz_3290;
  wire       [26:0]   _zz_3291;
  wire       [35:0]   _zz_3292;
  wire       [17:0]   _zz_3293;
  wire       [35:0]   _zz_3294;
  wire       [35:0]   _zz_3295;
  wire       [35:0]   _zz_3296;
  wire       [35:0]   _zz_3297;
  wire       [35:0]   _zz_3298;
  wire       [26:0]   _zz_3299;
  wire       [35:0]   _zz_3300;
  wire       [17:0]   _zz_3301;
  wire       [17:0]   _zz_3302;
  wire       [35:0]   _zz_3303;
  wire       [35:0]   _zz_3304;
  wire       [17:0]   _zz_3305;
  wire       [35:0]   _zz_3306;
  wire       [35:0]   _zz_3307;
  wire       [35:0]   _zz_3308;
  wire       [17:0]   _zz_3309;
  wire       [35:0]   _zz_3310;
  wire       [35:0]   _zz_3311;
  wire       [35:0]   _zz_3312;
  wire       [35:0]   _zz_3313;
  wire       [35:0]   _zz_3314;
  wire       [35:0]   _zz_3315;
  wire       [26:0]   _zz_3316;
  wire       [35:0]   _zz_3317;
  wire       [17:0]   _zz_3318;
  wire       [35:0]   _zz_3319;
  wire       [35:0]   _zz_3320;
  wire       [35:0]   _zz_3321;
  wire       [35:0]   _zz_3322;
  wire       [35:0]   _zz_3323;
  wire       [26:0]   _zz_3324;
  wire       [35:0]   _zz_3325;
  wire       [17:0]   _zz_3326;
  wire       [35:0]   _zz_3327;
  wire       [35:0]   _zz_3328;
  wire       [35:0]   _zz_3329;
  wire       [35:0]   _zz_3330;
  wire       [35:0]   _zz_3331;
  wire       [26:0]   _zz_3332;
  wire       [35:0]   _zz_3333;
  wire       [17:0]   _zz_3334;
  wire       [35:0]   _zz_3335;
  wire       [35:0]   _zz_3336;
  wire       [35:0]   _zz_3337;
  wire       [35:0]   _zz_3338;
  wire       [35:0]   _zz_3339;
  wire       [26:0]   _zz_3340;
  wire       [35:0]   _zz_3341;
  wire       [17:0]   _zz_3342;
  wire       [17:0]   _zz_3343;
  wire       [35:0]   _zz_3344;
  wire       [35:0]   _zz_3345;
  wire       [17:0]   _zz_3346;
  wire       [35:0]   _zz_3347;
  wire       [35:0]   _zz_3348;
  wire       [35:0]   _zz_3349;
  wire       [17:0]   _zz_3350;
  wire       [35:0]   _zz_3351;
  wire       [35:0]   _zz_3352;
  wire       [35:0]   _zz_3353;
  wire       [35:0]   _zz_3354;
  wire       [35:0]   _zz_3355;
  wire       [35:0]   _zz_3356;
  wire       [26:0]   _zz_3357;
  wire       [35:0]   _zz_3358;
  wire       [17:0]   _zz_3359;
  wire       [35:0]   _zz_3360;
  wire       [35:0]   _zz_3361;
  wire       [35:0]   _zz_3362;
  wire       [35:0]   _zz_3363;
  wire       [35:0]   _zz_3364;
  wire       [26:0]   _zz_3365;
  wire       [35:0]   _zz_3366;
  wire       [17:0]   _zz_3367;
  wire       [35:0]   _zz_3368;
  wire       [35:0]   _zz_3369;
  wire       [35:0]   _zz_3370;
  wire       [35:0]   _zz_3371;
  wire       [35:0]   _zz_3372;
  wire       [26:0]   _zz_3373;
  wire       [35:0]   _zz_3374;
  wire       [17:0]   _zz_3375;
  wire       [35:0]   _zz_3376;
  wire       [35:0]   _zz_3377;
  wire       [35:0]   _zz_3378;
  wire       [35:0]   _zz_3379;
  wire       [35:0]   _zz_3380;
  wire       [26:0]   _zz_3381;
  wire       [35:0]   _zz_3382;
  wire       [17:0]   _zz_3383;
  wire       [17:0]   _zz_3384;
  wire       [35:0]   _zz_3385;
  wire       [35:0]   _zz_3386;
  wire       [17:0]   _zz_3387;
  wire       [35:0]   _zz_3388;
  wire       [35:0]   _zz_3389;
  wire       [35:0]   _zz_3390;
  wire       [17:0]   _zz_3391;
  wire       [35:0]   _zz_3392;
  wire       [35:0]   _zz_3393;
  wire       [35:0]   _zz_3394;
  wire       [35:0]   _zz_3395;
  wire       [35:0]   _zz_3396;
  wire       [35:0]   _zz_3397;
  wire       [26:0]   _zz_3398;
  wire       [35:0]   _zz_3399;
  wire       [17:0]   _zz_3400;
  wire       [35:0]   _zz_3401;
  wire       [35:0]   _zz_3402;
  wire       [35:0]   _zz_3403;
  wire       [35:0]   _zz_3404;
  wire       [35:0]   _zz_3405;
  wire       [26:0]   _zz_3406;
  wire       [35:0]   _zz_3407;
  wire       [17:0]   _zz_3408;
  wire       [35:0]   _zz_3409;
  wire       [35:0]   _zz_3410;
  wire       [35:0]   _zz_3411;
  wire       [35:0]   _zz_3412;
  wire       [35:0]   _zz_3413;
  wire       [26:0]   _zz_3414;
  wire       [35:0]   _zz_3415;
  wire       [17:0]   _zz_3416;
  wire       [35:0]   _zz_3417;
  wire       [35:0]   _zz_3418;
  wire       [35:0]   _zz_3419;
  wire       [35:0]   _zz_3420;
  wire       [35:0]   _zz_3421;
  wire       [26:0]   _zz_3422;
  wire       [35:0]   _zz_3423;
  wire       [17:0]   _zz_3424;
  wire       [17:0]   _zz_3425;
  wire       [35:0]   _zz_3426;
  wire       [35:0]   _zz_3427;
  wire       [17:0]   _zz_3428;
  wire       [35:0]   _zz_3429;
  wire       [35:0]   _zz_3430;
  wire       [35:0]   _zz_3431;
  wire       [17:0]   _zz_3432;
  wire       [35:0]   _zz_3433;
  wire       [35:0]   _zz_3434;
  wire       [35:0]   _zz_3435;
  wire       [35:0]   _zz_3436;
  wire       [35:0]   _zz_3437;
  wire       [35:0]   _zz_3438;
  wire       [26:0]   _zz_3439;
  wire       [35:0]   _zz_3440;
  wire       [17:0]   _zz_3441;
  wire       [35:0]   _zz_3442;
  wire       [35:0]   _zz_3443;
  wire       [35:0]   _zz_3444;
  wire       [35:0]   _zz_3445;
  wire       [35:0]   _zz_3446;
  wire       [26:0]   _zz_3447;
  wire       [35:0]   _zz_3448;
  wire       [17:0]   _zz_3449;
  wire       [35:0]   _zz_3450;
  wire       [35:0]   _zz_3451;
  wire       [35:0]   _zz_3452;
  wire       [35:0]   _zz_3453;
  wire       [35:0]   _zz_3454;
  wire       [26:0]   _zz_3455;
  wire       [35:0]   _zz_3456;
  wire       [17:0]   _zz_3457;
  wire       [35:0]   _zz_3458;
  wire       [35:0]   _zz_3459;
  wire       [35:0]   _zz_3460;
  wire       [35:0]   _zz_3461;
  wire       [35:0]   _zz_3462;
  wire       [26:0]   _zz_3463;
  wire       [35:0]   _zz_3464;
  wire       [17:0]   _zz_3465;
  wire       [17:0]   _zz_3466;
  wire       [35:0]   _zz_3467;
  wire       [35:0]   _zz_3468;
  wire       [17:0]   _zz_3469;
  wire       [35:0]   _zz_3470;
  wire       [35:0]   _zz_3471;
  wire       [35:0]   _zz_3472;
  wire       [17:0]   _zz_3473;
  wire       [35:0]   _zz_3474;
  wire       [35:0]   _zz_3475;
  wire       [35:0]   _zz_3476;
  wire       [35:0]   _zz_3477;
  wire       [35:0]   _zz_3478;
  wire       [35:0]   _zz_3479;
  wire       [26:0]   _zz_3480;
  wire       [35:0]   _zz_3481;
  wire       [17:0]   _zz_3482;
  wire       [35:0]   _zz_3483;
  wire       [35:0]   _zz_3484;
  wire       [35:0]   _zz_3485;
  wire       [35:0]   _zz_3486;
  wire       [35:0]   _zz_3487;
  wire       [26:0]   _zz_3488;
  wire       [35:0]   _zz_3489;
  wire       [17:0]   _zz_3490;
  wire       [35:0]   _zz_3491;
  wire       [35:0]   _zz_3492;
  wire       [35:0]   _zz_3493;
  wire       [35:0]   _zz_3494;
  wire       [35:0]   _zz_3495;
  wire       [26:0]   _zz_3496;
  wire       [35:0]   _zz_3497;
  wire       [17:0]   _zz_3498;
  wire       [35:0]   _zz_3499;
  wire       [35:0]   _zz_3500;
  wire       [35:0]   _zz_3501;
  wire       [35:0]   _zz_3502;
  wire       [35:0]   _zz_3503;
  wire       [26:0]   _zz_3504;
  wire       [35:0]   _zz_3505;
  wire       [17:0]   _zz_3506;
  wire       [17:0]   _zz_3507;
  wire       [35:0]   _zz_3508;
  wire       [35:0]   _zz_3509;
  wire       [17:0]   _zz_3510;
  wire       [35:0]   _zz_3511;
  wire       [35:0]   _zz_3512;
  wire       [35:0]   _zz_3513;
  wire       [17:0]   _zz_3514;
  wire       [35:0]   _zz_3515;
  wire       [35:0]   _zz_3516;
  wire       [35:0]   _zz_3517;
  wire       [35:0]   _zz_3518;
  wire       [35:0]   _zz_3519;
  wire       [35:0]   _zz_3520;
  wire       [26:0]   _zz_3521;
  wire       [35:0]   _zz_3522;
  wire       [17:0]   _zz_3523;
  wire       [35:0]   _zz_3524;
  wire       [35:0]   _zz_3525;
  wire       [35:0]   _zz_3526;
  wire       [35:0]   _zz_3527;
  wire       [35:0]   _zz_3528;
  wire       [26:0]   _zz_3529;
  wire       [35:0]   _zz_3530;
  wire       [17:0]   _zz_3531;
  wire       [35:0]   _zz_3532;
  wire       [35:0]   _zz_3533;
  wire       [35:0]   _zz_3534;
  wire       [35:0]   _zz_3535;
  wire       [35:0]   _zz_3536;
  wire       [26:0]   _zz_3537;
  wire       [35:0]   _zz_3538;
  wire       [17:0]   _zz_3539;
  wire       [35:0]   _zz_3540;
  wire       [35:0]   _zz_3541;
  wire       [35:0]   _zz_3542;
  wire       [35:0]   _zz_3543;
  wire       [35:0]   _zz_3544;
  wire       [26:0]   _zz_3545;
  wire       [35:0]   _zz_3546;
  wire       [17:0]   _zz_3547;
  wire       [17:0]   _zz_3548;
  wire       [35:0]   _zz_3549;
  wire       [35:0]   _zz_3550;
  wire       [17:0]   _zz_3551;
  wire       [35:0]   _zz_3552;
  wire       [35:0]   _zz_3553;
  wire       [35:0]   _zz_3554;
  wire       [17:0]   _zz_3555;
  wire       [35:0]   _zz_3556;
  wire       [35:0]   _zz_3557;
  wire       [35:0]   _zz_3558;
  wire       [35:0]   _zz_3559;
  wire       [35:0]   _zz_3560;
  wire       [35:0]   _zz_3561;
  wire       [26:0]   _zz_3562;
  wire       [35:0]   _zz_3563;
  wire       [17:0]   _zz_3564;
  wire       [35:0]   _zz_3565;
  wire       [35:0]   _zz_3566;
  wire       [35:0]   _zz_3567;
  wire       [35:0]   _zz_3568;
  wire       [35:0]   _zz_3569;
  wire       [26:0]   _zz_3570;
  wire       [35:0]   _zz_3571;
  wire       [17:0]   _zz_3572;
  wire       [35:0]   _zz_3573;
  wire       [35:0]   _zz_3574;
  wire       [35:0]   _zz_3575;
  wire       [35:0]   _zz_3576;
  wire       [35:0]   _zz_3577;
  wire       [26:0]   _zz_3578;
  wire       [35:0]   _zz_3579;
  wire       [17:0]   _zz_3580;
  wire       [35:0]   _zz_3581;
  wire       [35:0]   _zz_3582;
  wire       [35:0]   _zz_3583;
  wire       [35:0]   _zz_3584;
  wire       [35:0]   _zz_3585;
  wire       [26:0]   _zz_3586;
  wire       [35:0]   _zz_3587;
  wire       [17:0]   _zz_3588;
  wire       [17:0]   _zz_3589;
  wire       [35:0]   _zz_3590;
  wire       [35:0]   _zz_3591;
  wire       [17:0]   _zz_3592;
  wire       [35:0]   _zz_3593;
  wire       [35:0]   _zz_3594;
  wire       [35:0]   _zz_3595;
  wire       [17:0]   _zz_3596;
  wire       [35:0]   _zz_3597;
  wire       [35:0]   _zz_3598;
  wire       [35:0]   _zz_3599;
  wire       [35:0]   _zz_3600;
  wire       [35:0]   _zz_3601;
  wire       [35:0]   _zz_3602;
  wire       [26:0]   _zz_3603;
  wire       [35:0]   _zz_3604;
  wire       [17:0]   _zz_3605;
  wire       [35:0]   _zz_3606;
  wire       [35:0]   _zz_3607;
  wire       [35:0]   _zz_3608;
  wire       [35:0]   _zz_3609;
  wire       [35:0]   _zz_3610;
  wire       [26:0]   _zz_3611;
  wire       [35:0]   _zz_3612;
  wire       [17:0]   _zz_3613;
  wire       [35:0]   _zz_3614;
  wire       [35:0]   _zz_3615;
  wire       [35:0]   _zz_3616;
  wire       [35:0]   _zz_3617;
  wire       [35:0]   _zz_3618;
  wire       [26:0]   _zz_3619;
  wire       [35:0]   _zz_3620;
  wire       [17:0]   _zz_3621;
  wire       [35:0]   _zz_3622;
  wire       [35:0]   _zz_3623;
  wire       [35:0]   _zz_3624;
  wire       [35:0]   _zz_3625;
  wire       [35:0]   _zz_3626;
  wire       [26:0]   _zz_3627;
  wire       [35:0]   _zz_3628;
  wire       [17:0]   _zz_3629;
  wire       [17:0]   _zz_3630;
  wire       [35:0]   _zz_3631;
  wire       [35:0]   _zz_3632;
  wire       [17:0]   _zz_3633;
  wire       [35:0]   _zz_3634;
  wire       [35:0]   _zz_3635;
  wire       [35:0]   _zz_3636;
  wire       [17:0]   _zz_3637;
  wire       [35:0]   _zz_3638;
  wire       [35:0]   _zz_3639;
  wire       [35:0]   _zz_3640;
  wire       [35:0]   _zz_3641;
  wire       [35:0]   _zz_3642;
  wire       [35:0]   _zz_3643;
  wire       [26:0]   _zz_3644;
  wire       [35:0]   _zz_3645;
  wire       [17:0]   _zz_3646;
  wire       [35:0]   _zz_3647;
  wire       [35:0]   _zz_3648;
  wire       [35:0]   _zz_3649;
  wire       [35:0]   _zz_3650;
  wire       [35:0]   _zz_3651;
  wire       [26:0]   _zz_3652;
  wire       [35:0]   _zz_3653;
  wire       [17:0]   _zz_3654;
  wire       [35:0]   _zz_3655;
  wire       [35:0]   _zz_3656;
  wire       [35:0]   _zz_3657;
  wire       [35:0]   _zz_3658;
  wire       [35:0]   _zz_3659;
  wire       [26:0]   _zz_3660;
  wire       [35:0]   _zz_3661;
  wire       [17:0]   _zz_3662;
  wire       [35:0]   _zz_3663;
  wire       [35:0]   _zz_3664;
  wire       [35:0]   _zz_3665;
  wire       [35:0]   _zz_3666;
  wire       [35:0]   _zz_3667;
  wire       [26:0]   _zz_3668;
  wire       [35:0]   _zz_3669;
  wire       [17:0]   _zz_3670;
  wire       [17:0]   _zz_3671;
  wire       [35:0]   _zz_3672;
  wire       [35:0]   _zz_3673;
  wire       [17:0]   _zz_3674;
  wire       [35:0]   _zz_3675;
  wire       [35:0]   _zz_3676;
  wire       [35:0]   _zz_3677;
  wire       [17:0]   _zz_3678;
  wire       [35:0]   _zz_3679;
  wire       [35:0]   _zz_3680;
  wire       [35:0]   _zz_3681;
  wire       [35:0]   _zz_3682;
  wire       [35:0]   _zz_3683;
  wire       [35:0]   _zz_3684;
  wire       [26:0]   _zz_3685;
  wire       [35:0]   _zz_3686;
  wire       [17:0]   _zz_3687;
  wire       [35:0]   _zz_3688;
  wire       [35:0]   _zz_3689;
  wire       [35:0]   _zz_3690;
  wire       [35:0]   _zz_3691;
  wire       [35:0]   _zz_3692;
  wire       [26:0]   _zz_3693;
  wire       [35:0]   _zz_3694;
  wire       [17:0]   _zz_3695;
  wire       [35:0]   _zz_3696;
  wire       [35:0]   _zz_3697;
  wire       [35:0]   _zz_3698;
  wire       [35:0]   _zz_3699;
  wire       [35:0]   _zz_3700;
  wire       [26:0]   _zz_3701;
  wire       [35:0]   _zz_3702;
  wire       [17:0]   _zz_3703;
  wire       [35:0]   _zz_3704;
  wire       [35:0]   _zz_3705;
  wire       [35:0]   _zz_3706;
  wire       [35:0]   _zz_3707;
  wire       [35:0]   _zz_3708;
  wire       [26:0]   _zz_3709;
  wire       [35:0]   _zz_3710;
  wire       [17:0]   _zz_3711;
  wire       [17:0]   _zz_3712;
  wire       [35:0]   _zz_3713;
  wire       [35:0]   _zz_3714;
  wire       [17:0]   _zz_3715;
  wire       [35:0]   _zz_3716;
  wire       [35:0]   _zz_3717;
  wire       [35:0]   _zz_3718;
  wire       [17:0]   _zz_3719;
  wire       [35:0]   _zz_3720;
  wire       [35:0]   _zz_3721;
  wire       [35:0]   _zz_3722;
  wire       [35:0]   _zz_3723;
  wire       [35:0]   _zz_3724;
  wire       [35:0]   _zz_3725;
  wire       [26:0]   _zz_3726;
  wire       [35:0]   _zz_3727;
  wire       [17:0]   _zz_3728;
  wire       [35:0]   _zz_3729;
  wire       [35:0]   _zz_3730;
  wire       [35:0]   _zz_3731;
  wire       [35:0]   _zz_3732;
  wire       [35:0]   _zz_3733;
  wire       [26:0]   _zz_3734;
  wire       [35:0]   _zz_3735;
  wire       [17:0]   _zz_3736;
  wire       [35:0]   _zz_3737;
  wire       [35:0]   _zz_3738;
  wire       [35:0]   _zz_3739;
  wire       [35:0]   _zz_3740;
  wire       [35:0]   _zz_3741;
  wire       [26:0]   _zz_3742;
  wire       [35:0]   _zz_3743;
  wire       [17:0]   _zz_3744;
  wire       [35:0]   _zz_3745;
  wire       [35:0]   _zz_3746;
  wire       [35:0]   _zz_3747;
  wire       [35:0]   _zz_3748;
  wire       [35:0]   _zz_3749;
  wire       [26:0]   _zz_3750;
  wire       [35:0]   _zz_3751;
  wire       [17:0]   _zz_3752;
  wire       [17:0]   _zz_3753;
  wire       [35:0]   _zz_3754;
  wire       [35:0]   _zz_3755;
  wire       [17:0]   _zz_3756;
  wire       [35:0]   _zz_3757;
  wire       [35:0]   _zz_3758;
  wire       [35:0]   _zz_3759;
  wire       [17:0]   _zz_3760;
  wire       [35:0]   _zz_3761;
  wire       [35:0]   _zz_3762;
  wire       [35:0]   _zz_3763;
  wire       [35:0]   _zz_3764;
  wire       [35:0]   _zz_3765;
  wire       [35:0]   _zz_3766;
  wire       [26:0]   _zz_3767;
  wire       [35:0]   _zz_3768;
  wire       [17:0]   _zz_3769;
  wire       [35:0]   _zz_3770;
  wire       [35:0]   _zz_3771;
  wire       [35:0]   _zz_3772;
  wire       [35:0]   _zz_3773;
  wire       [35:0]   _zz_3774;
  wire       [26:0]   _zz_3775;
  wire       [35:0]   _zz_3776;
  wire       [17:0]   _zz_3777;
  wire       [35:0]   _zz_3778;
  wire       [35:0]   _zz_3779;
  wire       [35:0]   _zz_3780;
  wire       [35:0]   _zz_3781;
  wire       [35:0]   _zz_3782;
  wire       [26:0]   _zz_3783;
  wire       [35:0]   _zz_3784;
  wire       [17:0]   _zz_3785;
  wire       [35:0]   _zz_3786;
  wire       [35:0]   _zz_3787;
  wire       [35:0]   _zz_3788;
  wire       [35:0]   _zz_3789;
  wire       [35:0]   _zz_3790;
  wire       [26:0]   _zz_3791;
  wire       [35:0]   _zz_3792;
  wire       [17:0]   _zz_3793;
  wire       [17:0]   _zz_3794;
  wire       [35:0]   _zz_3795;
  wire       [35:0]   _zz_3796;
  wire       [17:0]   _zz_3797;
  wire       [35:0]   _zz_3798;
  wire       [35:0]   _zz_3799;
  wire       [35:0]   _zz_3800;
  wire       [17:0]   _zz_3801;
  wire       [35:0]   _zz_3802;
  wire       [35:0]   _zz_3803;
  wire       [35:0]   _zz_3804;
  wire       [35:0]   _zz_3805;
  wire       [35:0]   _zz_3806;
  wire       [35:0]   _zz_3807;
  wire       [26:0]   _zz_3808;
  wire       [35:0]   _zz_3809;
  wire       [17:0]   _zz_3810;
  wire       [35:0]   _zz_3811;
  wire       [35:0]   _zz_3812;
  wire       [35:0]   _zz_3813;
  wire       [35:0]   _zz_3814;
  wire       [35:0]   _zz_3815;
  wire       [26:0]   _zz_3816;
  wire       [35:0]   _zz_3817;
  wire       [17:0]   _zz_3818;
  wire       [35:0]   _zz_3819;
  wire       [35:0]   _zz_3820;
  wire       [35:0]   _zz_3821;
  wire       [35:0]   _zz_3822;
  wire       [35:0]   _zz_3823;
  wire       [26:0]   _zz_3824;
  wire       [35:0]   _zz_3825;
  wire       [17:0]   _zz_3826;
  wire       [35:0]   _zz_3827;
  wire       [35:0]   _zz_3828;
  wire       [35:0]   _zz_3829;
  wire       [35:0]   _zz_3830;
  wire       [35:0]   _zz_3831;
  wire       [26:0]   _zz_3832;
  wire       [35:0]   _zz_3833;
  wire       [17:0]   _zz_3834;
  wire       [17:0]   _zz_3835;
  wire       [35:0]   _zz_3836;
  wire       [35:0]   _zz_3837;
  wire       [17:0]   _zz_3838;
  wire       [35:0]   _zz_3839;
  wire       [35:0]   _zz_3840;
  wire       [35:0]   _zz_3841;
  wire       [17:0]   _zz_3842;
  wire       [35:0]   _zz_3843;
  wire       [35:0]   _zz_3844;
  wire       [35:0]   _zz_3845;
  wire       [35:0]   _zz_3846;
  wire       [35:0]   _zz_3847;
  wire       [35:0]   _zz_3848;
  wire       [26:0]   _zz_3849;
  wire       [35:0]   _zz_3850;
  wire       [17:0]   _zz_3851;
  wire       [35:0]   _zz_3852;
  wire       [35:0]   _zz_3853;
  wire       [35:0]   _zz_3854;
  wire       [35:0]   _zz_3855;
  wire       [35:0]   _zz_3856;
  wire       [26:0]   _zz_3857;
  wire       [35:0]   _zz_3858;
  wire       [17:0]   _zz_3859;
  wire       [35:0]   _zz_3860;
  wire       [35:0]   _zz_3861;
  wire       [35:0]   _zz_3862;
  wire       [35:0]   _zz_3863;
  wire       [35:0]   _zz_3864;
  wire       [26:0]   _zz_3865;
  wire       [35:0]   _zz_3866;
  wire       [17:0]   _zz_3867;
  wire       [35:0]   _zz_3868;
  wire       [35:0]   _zz_3869;
  wire       [35:0]   _zz_3870;
  wire       [35:0]   _zz_3871;
  wire       [35:0]   _zz_3872;
  wire       [26:0]   _zz_3873;
  wire       [35:0]   _zz_3874;
  wire       [17:0]   _zz_3875;
  wire       [17:0]   _zz_3876;
  wire       [35:0]   _zz_3877;
  wire       [35:0]   _zz_3878;
  wire       [17:0]   _zz_3879;
  wire       [35:0]   _zz_3880;
  wire       [35:0]   _zz_3881;
  wire       [35:0]   _zz_3882;
  wire       [17:0]   _zz_3883;
  wire       [35:0]   _zz_3884;
  wire       [35:0]   _zz_3885;
  wire       [35:0]   _zz_3886;
  wire       [35:0]   _zz_3887;
  wire       [35:0]   _zz_3888;
  wire       [35:0]   _zz_3889;
  wire       [26:0]   _zz_3890;
  wire       [35:0]   _zz_3891;
  wire       [17:0]   _zz_3892;
  wire       [35:0]   _zz_3893;
  wire       [35:0]   _zz_3894;
  wire       [35:0]   _zz_3895;
  wire       [35:0]   _zz_3896;
  wire       [35:0]   _zz_3897;
  wire       [26:0]   _zz_3898;
  wire       [35:0]   _zz_3899;
  wire       [17:0]   _zz_3900;
  wire       [35:0]   _zz_3901;
  wire       [35:0]   _zz_3902;
  wire       [35:0]   _zz_3903;
  wire       [35:0]   _zz_3904;
  wire       [35:0]   _zz_3905;
  wire       [26:0]   _zz_3906;
  wire       [35:0]   _zz_3907;
  wire       [17:0]   _zz_3908;
  wire       [35:0]   _zz_3909;
  wire       [35:0]   _zz_3910;
  wire       [35:0]   _zz_3911;
  wire       [35:0]   _zz_3912;
  wire       [35:0]   _zz_3913;
  wire       [26:0]   _zz_3914;
  wire       [35:0]   _zz_3915;
  wire       [17:0]   _zz_3916;
  wire       [17:0]   _zz_3917;
  wire       [35:0]   _zz_3918;
  wire       [35:0]   _zz_3919;
  wire       [17:0]   _zz_3920;
  wire       [35:0]   _zz_3921;
  wire       [35:0]   _zz_3922;
  wire       [35:0]   _zz_3923;
  wire       [17:0]   _zz_3924;
  wire       [35:0]   _zz_3925;
  wire       [35:0]   _zz_3926;
  wire       [35:0]   _zz_3927;
  wire       [35:0]   _zz_3928;
  wire       [35:0]   _zz_3929;
  wire       [35:0]   _zz_3930;
  wire       [26:0]   _zz_3931;
  wire       [35:0]   _zz_3932;
  wire       [17:0]   _zz_3933;
  wire       [35:0]   _zz_3934;
  wire       [35:0]   _zz_3935;
  wire       [35:0]   _zz_3936;
  wire       [35:0]   _zz_3937;
  wire       [35:0]   _zz_3938;
  wire       [26:0]   _zz_3939;
  wire       [35:0]   _zz_3940;
  wire       [17:0]   _zz_3941;
  wire       [35:0]   _zz_3942;
  wire       [35:0]   _zz_3943;
  wire       [35:0]   _zz_3944;
  wire       [35:0]   _zz_3945;
  wire       [35:0]   _zz_3946;
  wire       [26:0]   _zz_3947;
  wire       [35:0]   _zz_3948;
  wire       [17:0]   _zz_3949;
  wire       [35:0]   _zz_3950;
  wire       [35:0]   _zz_3951;
  wire       [35:0]   _zz_3952;
  wire       [35:0]   _zz_3953;
  wire       [35:0]   _zz_3954;
  wire       [26:0]   _zz_3955;
  wire       [35:0]   _zz_3956;
  wire       [17:0]   _zz_3957;
  wire       [17:0]   _zz_3958;
  wire       [35:0]   _zz_3959;
  wire       [35:0]   _zz_3960;
  wire       [17:0]   _zz_3961;
  wire       [35:0]   _zz_3962;
  wire       [35:0]   _zz_3963;
  wire       [35:0]   _zz_3964;
  wire       [17:0]   _zz_3965;
  wire       [35:0]   _zz_3966;
  wire       [35:0]   _zz_3967;
  wire       [35:0]   _zz_3968;
  wire       [35:0]   _zz_3969;
  wire       [35:0]   _zz_3970;
  wire       [35:0]   _zz_3971;
  wire       [26:0]   _zz_3972;
  wire       [35:0]   _zz_3973;
  wire       [17:0]   _zz_3974;
  wire       [35:0]   _zz_3975;
  wire       [35:0]   _zz_3976;
  wire       [35:0]   _zz_3977;
  wire       [35:0]   _zz_3978;
  wire       [35:0]   _zz_3979;
  wire       [26:0]   _zz_3980;
  wire       [35:0]   _zz_3981;
  wire       [17:0]   _zz_3982;
  wire       [35:0]   _zz_3983;
  wire       [35:0]   _zz_3984;
  wire       [35:0]   _zz_3985;
  wire       [35:0]   _zz_3986;
  wire       [35:0]   _zz_3987;
  wire       [26:0]   _zz_3988;
  wire       [35:0]   _zz_3989;
  wire       [17:0]   _zz_3990;
  wire       [35:0]   _zz_3991;
  wire       [35:0]   _zz_3992;
  wire       [35:0]   _zz_3993;
  wire       [35:0]   _zz_3994;
  wire       [35:0]   _zz_3995;
  wire       [26:0]   _zz_3996;
  wire       [35:0]   _zz_3997;
  wire       [17:0]   _zz_3998;
  wire       [17:0]   _zz_3999;
  wire       [35:0]   _zz_4000;
  wire       [35:0]   _zz_4001;
  wire       [17:0]   _zz_4002;
  wire       [35:0]   _zz_4003;
  wire       [35:0]   _zz_4004;
  wire       [35:0]   _zz_4005;
  wire       [17:0]   _zz_4006;
  wire       [35:0]   _zz_4007;
  wire       [35:0]   _zz_4008;
  wire       [35:0]   _zz_4009;
  wire       [35:0]   _zz_4010;
  wire       [35:0]   _zz_4011;
  wire       [35:0]   _zz_4012;
  wire       [26:0]   _zz_4013;
  wire       [35:0]   _zz_4014;
  wire       [17:0]   _zz_4015;
  wire       [35:0]   _zz_4016;
  wire       [35:0]   _zz_4017;
  wire       [35:0]   _zz_4018;
  wire       [35:0]   _zz_4019;
  wire       [35:0]   _zz_4020;
  wire       [26:0]   _zz_4021;
  wire       [35:0]   _zz_4022;
  wire       [17:0]   _zz_4023;
  wire       [35:0]   _zz_4024;
  wire       [35:0]   _zz_4025;
  wire       [35:0]   _zz_4026;
  wire       [35:0]   _zz_4027;
  wire       [35:0]   _zz_4028;
  wire       [26:0]   _zz_4029;
  wire       [35:0]   _zz_4030;
  wire       [17:0]   _zz_4031;
  wire       [35:0]   _zz_4032;
  wire       [35:0]   _zz_4033;
  wire       [35:0]   _zz_4034;
  wire       [35:0]   _zz_4035;
  wire       [35:0]   _zz_4036;
  wire       [26:0]   _zz_4037;
  wire       [35:0]   _zz_4038;
  wire       [17:0]   _zz_4039;
  wire       [17:0]   _zz_4040;
  wire       [35:0]   _zz_4041;
  wire       [35:0]   _zz_4042;
  wire       [17:0]   _zz_4043;
  wire       [35:0]   _zz_4044;
  wire       [35:0]   _zz_4045;
  wire       [35:0]   _zz_4046;
  wire       [17:0]   _zz_4047;
  wire       [35:0]   _zz_4048;
  wire       [35:0]   _zz_4049;
  wire       [35:0]   _zz_4050;
  wire       [35:0]   _zz_4051;
  wire       [35:0]   _zz_4052;
  wire       [35:0]   _zz_4053;
  wire       [26:0]   _zz_4054;
  wire       [35:0]   _zz_4055;
  wire       [17:0]   _zz_4056;
  wire       [35:0]   _zz_4057;
  wire       [35:0]   _zz_4058;
  wire       [35:0]   _zz_4059;
  wire       [35:0]   _zz_4060;
  wire       [35:0]   _zz_4061;
  wire       [26:0]   _zz_4062;
  wire       [35:0]   _zz_4063;
  wire       [17:0]   _zz_4064;
  wire       [35:0]   _zz_4065;
  wire       [35:0]   _zz_4066;
  wire       [35:0]   _zz_4067;
  wire       [35:0]   _zz_4068;
  wire       [35:0]   _zz_4069;
  wire       [26:0]   _zz_4070;
  wire       [35:0]   _zz_4071;
  wire       [17:0]   _zz_4072;
  wire       [35:0]   _zz_4073;
  wire       [35:0]   _zz_4074;
  wire       [35:0]   _zz_4075;
  wire       [35:0]   _zz_4076;
  wire       [35:0]   _zz_4077;
  wire       [26:0]   _zz_4078;
  wire       [35:0]   _zz_4079;
  wire       [17:0]   _zz_4080;
  wire       [17:0]   _zz_4081;
  wire       [35:0]   _zz_4082;
  wire       [35:0]   _zz_4083;
  wire       [17:0]   _zz_4084;
  wire       [35:0]   _zz_4085;
  wire       [35:0]   _zz_4086;
  wire       [35:0]   _zz_4087;
  wire       [17:0]   _zz_4088;
  wire       [35:0]   _zz_4089;
  wire       [35:0]   _zz_4090;
  wire       [35:0]   _zz_4091;
  wire       [35:0]   _zz_4092;
  wire       [35:0]   _zz_4093;
  wire       [35:0]   _zz_4094;
  wire       [26:0]   _zz_4095;
  wire       [35:0]   _zz_4096;
  wire       [17:0]   _zz_4097;
  wire       [35:0]   _zz_4098;
  wire       [35:0]   _zz_4099;
  wire       [35:0]   _zz_4100;
  wire       [35:0]   _zz_4101;
  wire       [35:0]   _zz_4102;
  wire       [26:0]   _zz_4103;
  wire       [35:0]   _zz_4104;
  wire       [17:0]   _zz_4105;
  wire       [35:0]   _zz_4106;
  wire       [35:0]   _zz_4107;
  wire       [35:0]   _zz_4108;
  wire       [35:0]   _zz_4109;
  wire       [35:0]   _zz_4110;
  wire       [26:0]   _zz_4111;
  wire       [35:0]   _zz_4112;
  wire       [17:0]   _zz_4113;
  wire       [35:0]   _zz_4114;
  wire       [35:0]   _zz_4115;
  wire       [35:0]   _zz_4116;
  wire       [35:0]   _zz_4117;
  wire       [35:0]   _zz_4118;
  wire       [26:0]   _zz_4119;
  wire       [35:0]   _zz_4120;
  wire       [17:0]   _zz_4121;
  wire       [17:0]   _zz_4122;
  wire       [35:0]   _zz_4123;
  wire       [35:0]   _zz_4124;
  wire       [17:0]   _zz_4125;
  wire       [35:0]   _zz_4126;
  wire       [35:0]   _zz_4127;
  wire       [35:0]   _zz_4128;
  wire       [17:0]   _zz_4129;
  wire       [35:0]   _zz_4130;
  wire       [35:0]   _zz_4131;
  wire       [35:0]   _zz_4132;
  wire       [35:0]   _zz_4133;
  wire       [35:0]   _zz_4134;
  wire       [35:0]   _zz_4135;
  wire       [26:0]   _zz_4136;
  wire       [35:0]   _zz_4137;
  wire       [17:0]   _zz_4138;
  wire       [35:0]   _zz_4139;
  wire       [35:0]   _zz_4140;
  wire       [35:0]   _zz_4141;
  wire       [35:0]   _zz_4142;
  wire       [35:0]   _zz_4143;
  wire       [26:0]   _zz_4144;
  wire       [35:0]   _zz_4145;
  wire       [17:0]   _zz_4146;
  wire       [35:0]   _zz_4147;
  wire       [35:0]   _zz_4148;
  wire       [35:0]   _zz_4149;
  wire       [35:0]   _zz_4150;
  wire       [35:0]   _zz_4151;
  wire       [26:0]   _zz_4152;
  wire       [35:0]   _zz_4153;
  wire       [17:0]   _zz_4154;
  wire       [35:0]   _zz_4155;
  wire       [35:0]   _zz_4156;
  wire       [35:0]   _zz_4157;
  wire       [35:0]   _zz_4158;
  wire       [35:0]   _zz_4159;
  wire       [26:0]   _zz_4160;
  wire       [35:0]   _zz_4161;
  wire       [17:0]   _zz_4162;
  wire       [17:0]   _zz_4163;
  wire       [35:0]   _zz_4164;
  wire       [35:0]   _zz_4165;
  wire       [17:0]   _zz_4166;
  wire       [35:0]   _zz_4167;
  wire       [35:0]   _zz_4168;
  wire       [35:0]   _zz_4169;
  wire       [17:0]   _zz_4170;
  wire       [35:0]   _zz_4171;
  wire       [35:0]   _zz_4172;
  wire       [35:0]   _zz_4173;
  wire       [35:0]   _zz_4174;
  wire       [35:0]   _zz_4175;
  wire       [35:0]   _zz_4176;
  wire       [26:0]   _zz_4177;
  wire       [35:0]   _zz_4178;
  wire       [17:0]   _zz_4179;
  wire       [35:0]   _zz_4180;
  wire       [35:0]   _zz_4181;
  wire       [35:0]   _zz_4182;
  wire       [35:0]   _zz_4183;
  wire       [35:0]   _zz_4184;
  wire       [26:0]   _zz_4185;
  wire       [35:0]   _zz_4186;
  wire       [17:0]   _zz_4187;
  wire       [35:0]   _zz_4188;
  wire       [35:0]   _zz_4189;
  wire       [35:0]   _zz_4190;
  wire       [35:0]   _zz_4191;
  wire       [35:0]   _zz_4192;
  wire       [26:0]   _zz_4193;
  wire       [35:0]   _zz_4194;
  wire       [17:0]   _zz_4195;
  wire       [35:0]   _zz_4196;
  wire       [35:0]   _zz_4197;
  wire       [35:0]   _zz_4198;
  wire       [35:0]   _zz_4199;
  wire       [35:0]   _zz_4200;
  wire       [26:0]   _zz_4201;
  wire       [35:0]   _zz_4202;
  wire       [17:0]   _zz_4203;
  wire       [17:0]   _zz_4204;
  wire       [35:0]   _zz_4205;
  wire       [35:0]   _zz_4206;
  wire       [17:0]   _zz_4207;
  wire       [35:0]   _zz_4208;
  wire       [35:0]   _zz_4209;
  wire       [35:0]   _zz_4210;
  wire       [17:0]   _zz_4211;
  wire       [35:0]   _zz_4212;
  wire       [35:0]   _zz_4213;
  wire       [35:0]   _zz_4214;
  wire       [35:0]   _zz_4215;
  wire       [35:0]   _zz_4216;
  wire       [35:0]   _zz_4217;
  wire       [26:0]   _zz_4218;
  wire       [35:0]   _zz_4219;
  wire       [17:0]   _zz_4220;
  wire       [35:0]   _zz_4221;
  wire       [35:0]   _zz_4222;
  wire       [35:0]   _zz_4223;
  wire       [35:0]   _zz_4224;
  wire       [35:0]   _zz_4225;
  wire       [26:0]   _zz_4226;
  wire       [35:0]   _zz_4227;
  wire       [17:0]   _zz_4228;
  wire       [35:0]   _zz_4229;
  wire       [35:0]   _zz_4230;
  wire       [35:0]   _zz_4231;
  wire       [35:0]   _zz_4232;
  wire       [35:0]   _zz_4233;
  wire       [26:0]   _zz_4234;
  wire       [35:0]   _zz_4235;
  wire       [17:0]   _zz_4236;
  wire       [35:0]   _zz_4237;
  wire       [35:0]   _zz_4238;
  wire       [35:0]   _zz_4239;
  wire       [35:0]   _zz_4240;
  wire       [35:0]   _zz_4241;
  wire       [26:0]   _zz_4242;
  wire       [35:0]   _zz_4243;
  wire       [17:0]   _zz_4244;
  wire       [17:0]   _zz_4245;
  wire       [35:0]   _zz_4246;
  wire       [35:0]   _zz_4247;
  wire       [17:0]   _zz_4248;
  wire       [35:0]   _zz_4249;
  wire       [35:0]   _zz_4250;
  wire       [35:0]   _zz_4251;
  wire       [17:0]   _zz_4252;
  wire       [35:0]   _zz_4253;
  wire       [35:0]   _zz_4254;
  wire       [35:0]   _zz_4255;
  wire       [35:0]   _zz_4256;
  wire       [35:0]   _zz_4257;
  wire       [35:0]   _zz_4258;
  wire       [26:0]   _zz_4259;
  wire       [35:0]   _zz_4260;
  wire       [17:0]   _zz_4261;
  wire       [35:0]   _zz_4262;
  wire       [35:0]   _zz_4263;
  wire       [35:0]   _zz_4264;
  wire       [35:0]   _zz_4265;
  wire       [35:0]   _zz_4266;
  wire       [26:0]   _zz_4267;
  wire       [35:0]   _zz_4268;
  wire       [17:0]   _zz_4269;
  wire       [35:0]   _zz_4270;
  wire       [35:0]   _zz_4271;
  wire       [35:0]   _zz_4272;
  wire       [35:0]   _zz_4273;
  wire       [35:0]   _zz_4274;
  wire       [26:0]   _zz_4275;
  wire       [35:0]   _zz_4276;
  wire       [17:0]   _zz_4277;
  wire       [35:0]   _zz_4278;
  wire       [35:0]   _zz_4279;
  wire       [35:0]   _zz_4280;
  wire       [35:0]   _zz_4281;
  wire       [35:0]   _zz_4282;
  wire       [26:0]   _zz_4283;
  wire       [35:0]   _zz_4284;
  wire       [17:0]   _zz_4285;
  wire       [17:0]   _zz_4286;
  wire       [35:0]   _zz_4287;
  wire       [35:0]   _zz_4288;
  wire       [17:0]   _zz_4289;
  wire       [35:0]   _zz_4290;
  wire       [35:0]   _zz_4291;
  wire       [35:0]   _zz_4292;
  wire       [17:0]   _zz_4293;
  wire       [35:0]   _zz_4294;
  wire       [35:0]   _zz_4295;
  wire       [35:0]   _zz_4296;
  wire       [35:0]   _zz_4297;
  wire       [35:0]   _zz_4298;
  wire       [35:0]   _zz_4299;
  wire       [26:0]   _zz_4300;
  wire       [35:0]   _zz_4301;
  wire       [17:0]   _zz_4302;
  wire       [35:0]   _zz_4303;
  wire       [35:0]   _zz_4304;
  wire       [35:0]   _zz_4305;
  wire       [35:0]   _zz_4306;
  wire       [35:0]   _zz_4307;
  wire       [26:0]   _zz_4308;
  wire       [35:0]   _zz_4309;
  wire       [17:0]   _zz_4310;
  wire       [35:0]   _zz_4311;
  wire       [35:0]   _zz_4312;
  wire       [35:0]   _zz_4313;
  wire       [35:0]   _zz_4314;
  wire       [35:0]   _zz_4315;
  wire       [26:0]   _zz_4316;
  wire       [35:0]   _zz_4317;
  wire       [17:0]   _zz_4318;
  wire       [35:0]   _zz_4319;
  wire       [35:0]   _zz_4320;
  wire       [35:0]   _zz_4321;
  wire       [35:0]   _zz_4322;
  wire       [35:0]   _zz_4323;
  wire       [26:0]   _zz_4324;
  wire       [35:0]   _zz_4325;
  wire       [17:0]   _zz_4326;
  wire       [17:0]   _zz_4327;
  wire       [35:0]   _zz_4328;
  wire       [35:0]   _zz_4329;
  wire       [17:0]   _zz_4330;
  wire       [35:0]   _zz_4331;
  wire       [35:0]   _zz_4332;
  wire       [35:0]   _zz_4333;
  wire       [17:0]   _zz_4334;
  wire       [35:0]   _zz_4335;
  wire       [35:0]   _zz_4336;
  wire       [35:0]   _zz_4337;
  wire       [35:0]   _zz_4338;
  wire       [35:0]   _zz_4339;
  wire       [35:0]   _zz_4340;
  wire       [26:0]   _zz_4341;
  wire       [35:0]   _zz_4342;
  wire       [17:0]   _zz_4343;
  wire       [35:0]   _zz_4344;
  wire       [35:0]   _zz_4345;
  wire       [35:0]   _zz_4346;
  wire       [35:0]   _zz_4347;
  wire       [35:0]   _zz_4348;
  wire       [26:0]   _zz_4349;
  wire       [35:0]   _zz_4350;
  wire       [17:0]   _zz_4351;
  wire       [35:0]   _zz_4352;
  wire       [35:0]   _zz_4353;
  wire       [35:0]   _zz_4354;
  wire       [35:0]   _zz_4355;
  wire       [35:0]   _zz_4356;
  wire       [26:0]   _zz_4357;
  wire       [35:0]   _zz_4358;
  wire       [17:0]   _zz_4359;
  wire       [35:0]   _zz_4360;
  wire       [35:0]   _zz_4361;
  wire       [35:0]   _zz_4362;
  wire       [35:0]   _zz_4363;
  wire       [35:0]   _zz_4364;
  wire       [26:0]   _zz_4365;
  wire       [35:0]   _zz_4366;
  wire       [17:0]   _zz_4367;
  wire       [17:0]   _zz_4368;
  wire       [35:0]   _zz_4369;
  wire       [35:0]   _zz_4370;
  wire       [17:0]   _zz_4371;
  wire       [35:0]   _zz_4372;
  wire       [35:0]   _zz_4373;
  wire       [35:0]   _zz_4374;
  wire       [17:0]   _zz_4375;
  wire       [35:0]   _zz_4376;
  wire       [35:0]   _zz_4377;
  wire       [35:0]   _zz_4378;
  wire       [35:0]   _zz_4379;
  wire       [35:0]   _zz_4380;
  wire       [35:0]   _zz_4381;
  wire       [26:0]   _zz_4382;
  wire       [35:0]   _zz_4383;
  wire       [17:0]   _zz_4384;
  wire       [35:0]   _zz_4385;
  wire       [35:0]   _zz_4386;
  wire       [35:0]   _zz_4387;
  wire       [35:0]   _zz_4388;
  wire       [35:0]   _zz_4389;
  wire       [26:0]   _zz_4390;
  wire       [35:0]   _zz_4391;
  wire       [17:0]   _zz_4392;
  wire       [35:0]   _zz_4393;
  wire       [35:0]   _zz_4394;
  wire       [35:0]   _zz_4395;
  wire       [35:0]   _zz_4396;
  wire       [35:0]   _zz_4397;
  wire       [26:0]   _zz_4398;
  wire       [35:0]   _zz_4399;
  wire       [17:0]   _zz_4400;
  wire       [35:0]   _zz_4401;
  wire       [35:0]   _zz_4402;
  wire       [35:0]   _zz_4403;
  wire       [35:0]   _zz_4404;
  wire       [35:0]   _zz_4405;
  wire       [26:0]   _zz_4406;
  wire       [35:0]   _zz_4407;
  wire       [17:0]   _zz_4408;
  wire       [17:0]   _zz_4409;
  wire       [35:0]   _zz_4410;
  wire       [35:0]   _zz_4411;
  wire       [17:0]   _zz_4412;
  wire       [35:0]   _zz_4413;
  wire       [35:0]   _zz_4414;
  wire       [35:0]   _zz_4415;
  wire       [17:0]   _zz_4416;
  wire       [35:0]   _zz_4417;
  wire       [35:0]   _zz_4418;
  wire       [35:0]   _zz_4419;
  wire       [35:0]   _zz_4420;
  wire       [35:0]   _zz_4421;
  wire       [35:0]   _zz_4422;
  wire       [26:0]   _zz_4423;
  wire       [35:0]   _zz_4424;
  wire       [17:0]   _zz_4425;
  wire       [35:0]   _zz_4426;
  wire       [35:0]   _zz_4427;
  wire       [35:0]   _zz_4428;
  wire       [35:0]   _zz_4429;
  wire       [35:0]   _zz_4430;
  wire       [26:0]   _zz_4431;
  wire       [35:0]   _zz_4432;
  wire       [17:0]   _zz_4433;
  wire       [35:0]   _zz_4434;
  wire       [35:0]   _zz_4435;
  wire       [35:0]   _zz_4436;
  wire       [35:0]   _zz_4437;
  wire       [35:0]   _zz_4438;
  wire       [26:0]   _zz_4439;
  wire       [35:0]   _zz_4440;
  wire       [17:0]   _zz_4441;
  wire       [35:0]   _zz_4442;
  wire       [35:0]   _zz_4443;
  wire       [35:0]   _zz_4444;
  wire       [35:0]   _zz_4445;
  wire       [35:0]   _zz_4446;
  wire       [26:0]   _zz_4447;
  wire       [35:0]   _zz_4448;
  wire       [17:0]   _zz_4449;
  wire       [17:0]   _zz_4450;
  wire       [35:0]   _zz_4451;
  wire       [35:0]   _zz_4452;
  wire       [17:0]   _zz_4453;
  wire       [35:0]   _zz_4454;
  wire       [35:0]   _zz_4455;
  wire       [35:0]   _zz_4456;
  wire       [17:0]   _zz_4457;
  wire       [35:0]   _zz_4458;
  wire       [35:0]   _zz_4459;
  wire       [35:0]   _zz_4460;
  wire       [35:0]   _zz_4461;
  wire       [35:0]   _zz_4462;
  wire       [35:0]   _zz_4463;
  wire       [26:0]   _zz_4464;
  wire       [35:0]   _zz_4465;
  wire       [17:0]   _zz_4466;
  wire       [35:0]   _zz_4467;
  wire       [35:0]   _zz_4468;
  wire       [35:0]   _zz_4469;
  wire       [35:0]   _zz_4470;
  wire       [35:0]   _zz_4471;
  wire       [26:0]   _zz_4472;
  wire       [35:0]   _zz_4473;
  wire       [17:0]   _zz_4474;
  wire       [35:0]   _zz_4475;
  wire       [35:0]   _zz_4476;
  wire       [35:0]   _zz_4477;
  wire       [35:0]   _zz_4478;
  wire       [35:0]   _zz_4479;
  wire       [26:0]   _zz_4480;
  wire       [35:0]   _zz_4481;
  wire       [17:0]   _zz_4482;
  wire       [35:0]   _zz_4483;
  wire       [35:0]   _zz_4484;
  wire       [35:0]   _zz_4485;
  wire       [35:0]   _zz_4486;
  wire       [35:0]   _zz_4487;
  wire       [26:0]   _zz_4488;
  wire       [35:0]   _zz_4489;
  wire       [17:0]   _zz_4490;
  wire       [17:0]   _zz_4491;
  wire       [35:0]   _zz_4492;
  wire       [35:0]   _zz_4493;
  wire       [17:0]   _zz_4494;
  wire       [35:0]   _zz_4495;
  wire       [35:0]   _zz_4496;
  wire       [35:0]   _zz_4497;
  wire       [17:0]   _zz_4498;
  wire       [35:0]   _zz_4499;
  wire       [35:0]   _zz_4500;
  wire       [35:0]   _zz_4501;
  wire       [35:0]   _zz_4502;
  wire       [35:0]   _zz_4503;
  wire       [35:0]   _zz_4504;
  wire       [26:0]   _zz_4505;
  wire       [35:0]   _zz_4506;
  wire       [17:0]   _zz_4507;
  wire       [35:0]   _zz_4508;
  wire       [35:0]   _zz_4509;
  wire       [35:0]   _zz_4510;
  wire       [35:0]   _zz_4511;
  wire       [35:0]   _zz_4512;
  wire       [26:0]   _zz_4513;
  wire       [35:0]   _zz_4514;
  wire       [17:0]   _zz_4515;
  wire       [35:0]   _zz_4516;
  wire       [35:0]   _zz_4517;
  wire       [35:0]   _zz_4518;
  wire       [35:0]   _zz_4519;
  wire       [35:0]   _zz_4520;
  wire       [26:0]   _zz_4521;
  wire       [35:0]   _zz_4522;
  wire       [17:0]   _zz_4523;
  wire       [35:0]   _zz_4524;
  wire       [35:0]   _zz_4525;
  wire       [35:0]   _zz_4526;
  wire       [35:0]   _zz_4527;
  wire       [35:0]   _zz_4528;
  wire       [26:0]   _zz_4529;
  wire       [35:0]   _zz_4530;
  wire       [17:0]   _zz_4531;
  wire       [17:0]   _zz_4532;
  wire       [35:0]   _zz_4533;
  wire       [35:0]   _zz_4534;
  wire       [17:0]   _zz_4535;
  wire       [35:0]   _zz_4536;
  wire       [35:0]   _zz_4537;
  wire       [35:0]   _zz_4538;
  wire       [17:0]   _zz_4539;
  wire       [35:0]   _zz_4540;
  wire       [35:0]   _zz_4541;
  wire       [35:0]   _zz_4542;
  wire       [35:0]   _zz_4543;
  wire       [35:0]   _zz_4544;
  wire       [35:0]   _zz_4545;
  wire       [26:0]   _zz_4546;
  wire       [35:0]   _zz_4547;
  wire       [17:0]   _zz_4548;
  wire       [35:0]   _zz_4549;
  wire       [35:0]   _zz_4550;
  wire       [35:0]   _zz_4551;
  wire       [35:0]   _zz_4552;
  wire       [35:0]   _zz_4553;
  wire       [26:0]   _zz_4554;
  wire       [35:0]   _zz_4555;
  wire       [17:0]   _zz_4556;
  wire       [35:0]   _zz_4557;
  wire       [35:0]   _zz_4558;
  wire       [35:0]   _zz_4559;
  wire       [35:0]   _zz_4560;
  wire       [35:0]   _zz_4561;
  wire       [26:0]   _zz_4562;
  wire       [35:0]   _zz_4563;
  wire       [17:0]   _zz_4564;
  wire       [35:0]   _zz_4565;
  wire       [35:0]   _zz_4566;
  wire       [35:0]   _zz_4567;
  wire       [35:0]   _zz_4568;
  wire       [35:0]   _zz_4569;
  wire       [26:0]   _zz_4570;
  wire       [35:0]   _zz_4571;
  wire       [17:0]   _zz_4572;
  wire       [17:0]   _zz_4573;
  wire       [35:0]   _zz_4574;
  wire       [35:0]   _zz_4575;
  wire       [17:0]   _zz_4576;
  wire       [35:0]   _zz_4577;
  wire       [35:0]   _zz_4578;
  wire       [35:0]   _zz_4579;
  wire       [17:0]   _zz_4580;
  wire       [35:0]   _zz_4581;
  wire       [35:0]   _zz_4582;
  wire       [35:0]   _zz_4583;
  wire       [35:0]   _zz_4584;
  wire       [35:0]   _zz_4585;
  wire       [35:0]   _zz_4586;
  wire       [26:0]   _zz_4587;
  wire       [35:0]   _zz_4588;
  wire       [17:0]   _zz_4589;
  wire       [35:0]   _zz_4590;
  wire       [35:0]   _zz_4591;
  wire       [35:0]   _zz_4592;
  wire       [35:0]   _zz_4593;
  wire       [35:0]   _zz_4594;
  wire       [26:0]   _zz_4595;
  wire       [35:0]   _zz_4596;
  wire       [17:0]   _zz_4597;
  wire       [35:0]   _zz_4598;
  wire       [35:0]   _zz_4599;
  wire       [35:0]   _zz_4600;
  wire       [35:0]   _zz_4601;
  wire       [35:0]   _zz_4602;
  wire       [26:0]   _zz_4603;
  wire       [35:0]   _zz_4604;
  wire       [17:0]   _zz_4605;
  wire       [35:0]   _zz_4606;
  wire       [35:0]   _zz_4607;
  wire       [35:0]   _zz_4608;
  wire       [35:0]   _zz_4609;
  wire       [35:0]   _zz_4610;
  wire       [26:0]   _zz_4611;
  wire       [35:0]   _zz_4612;
  wire       [17:0]   _zz_4613;
  wire       [17:0]   _zz_4614;
  wire       [35:0]   _zz_4615;
  wire       [35:0]   _zz_4616;
  wire       [17:0]   _zz_4617;
  wire       [35:0]   _zz_4618;
  wire       [35:0]   _zz_4619;
  wire       [35:0]   _zz_4620;
  wire       [17:0]   _zz_4621;
  wire       [35:0]   _zz_4622;
  wire       [35:0]   _zz_4623;
  wire       [35:0]   _zz_4624;
  wire       [35:0]   _zz_4625;
  wire       [35:0]   _zz_4626;
  wire       [35:0]   _zz_4627;
  wire       [26:0]   _zz_4628;
  wire       [35:0]   _zz_4629;
  wire       [17:0]   _zz_4630;
  wire       [35:0]   _zz_4631;
  wire       [35:0]   _zz_4632;
  wire       [35:0]   _zz_4633;
  wire       [35:0]   _zz_4634;
  wire       [35:0]   _zz_4635;
  wire       [26:0]   _zz_4636;
  wire       [35:0]   _zz_4637;
  wire       [17:0]   _zz_4638;
  wire       [35:0]   _zz_4639;
  wire       [35:0]   _zz_4640;
  wire       [35:0]   _zz_4641;
  wire       [35:0]   _zz_4642;
  wire       [35:0]   _zz_4643;
  wire       [26:0]   _zz_4644;
  wire       [35:0]   _zz_4645;
  wire       [17:0]   _zz_4646;
  wire       [35:0]   _zz_4647;
  wire       [35:0]   _zz_4648;
  wire       [35:0]   _zz_4649;
  wire       [35:0]   _zz_4650;
  wire       [35:0]   _zz_4651;
  wire       [26:0]   _zz_4652;
  wire       [35:0]   _zz_4653;
  wire       [17:0]   _zz_4654;
  wire       [17:0]   _zz_4655;
  wire       [35:0]   _zz_4656;
  wire       [35:0]   _zz_4657;
  wire       [17:0]   _zz_4658;
  wire       [35:0]   _zz_4659;
  wire       [35:0]   _zz_4660;
  wire       [35:0]   _zz_4661;
  wire       [17:0]   _zz_4662;
  wire       [35:0]   _zz_4663;
  wire       [35:0]   _zz_4664;
  wire       [35:0]   _zz_4665;
  wire       [35:0]   _zz_4666;
  wire       [35:0]   _zz_4667;
  wire       [35:0]   _zz_4668;
  wire       [26:0]   _zz_4669;
  wire       [35:0]   _zz_4670;
  wire       [17:0]   _zz_4671;
  wire       [35:0]   _zz_4672;
  wire       [35:0]   _zz_4673;
  wire       [35:0]   _zz_4674;
  wire       [35:0]   _zz_4675;
  wire       [35:0]   _zz_4676;
  wire       [26:0]   _zz_4677;
  wire       [35:0]   _zz_4678;
  wire       [17:0]   _zz_4679;
  wire       [35:0]   _zz_4680;
  wire       [35:0]   _zz_4681;
  wire       [35:0]   _zz_4682;
  wire       [35:0]   _zz_4683;
  wire       [35:0]   _zz_4684;
  wire       [26:0]   _zz_4685;
  wire       [35:0]   _zz_4686;
  wire       [17:0]   _zz_4687;
  wire       [35:0]   _zz_4688;
  wire       [35:0]   _zz_4689;
  wire       [35:0]   _zz_4690;
  wire       [35:0]   _zz_4691;
  wire       [35:0]   _zz_4692;
  wire       [26:0]   _zz_4693;
  wire       [35:0]   _zz_4694;
  wire       [17:0]   _zz_4695;
  wire       [17:0]   _zz_4696;
  wire       [35:0]   _zz_4697;
  wire       [35:0]   _zz_4698;
  wire       [17:0]   _zz_4699;
  wire       [35:0]   _zz_4700;
  wire       [35:0]   _zz_4701;
  wire       [35:0]   _zz_4702;
  wire       [17:0]   _zz_4703;
  wire       [35:0]   _zz_4704;
  wire       [35:0]   _zz_4705;
  wire       [35:0]   _zz_4706;
  wire       [35:0]   _zz_4707;
  wire       [35:0]   _zz_4708;
  wire       [35:0]   _zz_4709;
  wire       [26:0]   _zz_4710;
  wire       [35:0]   _zz_4711;
  wire       [17:0]   _zz_4712;
  wire       [35:0]   _zz_4713;
  wire       [35:0]   _zz_4714;
  wire       [35:0]   _zz_4715;
  wire       [35:0]   _zz_4716;
  wire       [35:0]   _zz_4717;
  wire       [26:0]   _zz_4718;
  wire       [35:0]   _zz_4719;
  wire       [17:0]   _zz_4720;
  wire       [35:0]   _zz_4721;
  wire       [35:0]   _zz_4722;
  wire       [35:0]   _zz_4723;
  wire       [35:0]   _zz_4724;
  wire       [35:0]   _zz_4725;
  wire       [26:0]   _zz_4726;
  wire       [35:0]   _zz_4727;
  wire       [17:0]   _zz_4728;
  wire       [35:0]   _zz_4729;
  wire       [35:0]   _zz_4730;
  wire       [35:0]   _zz_4731;
  wire       [35:0]   _zz_4732;
  wire       [35:0]   _zz_4733;
  wire       [26:0]   _zz_4734;
  wire       [35:0]   _zz_4735;
  wire       [17:0]   _zz_4736;
  wire       [17:0]   _zz_4737;
  wire       [35:0]   _zz_4738;
  wire       [35:0]   _zz_4739;
  wire       [17:0]   _zz_4740;
  wire       [35:0]   _zz_4741;
  wire       [35:0]   _zz_4742;
  wire       [35:0]   _zz_4743;
  wire       [17:0]   _zz_4744;
  wire       [35:0]   _zz_4745;
  wire       [35:0]   _zz_4746;
  wire       [35:0]   _zz_4747;
  wire       [35:0]   _zz_4748;
  wire       [35:0]   _zz_4749;
  wire       [35:0]   _zz_4750;
  wire       [26:0]   _zz_4751;
  wire       [35:0]   _zz_4752;
  wire       [17:0]   _zz_4753;
  wire       [35:0]   _zz_4754;
  wire       [35:0]   _zz_4755;
  wire       [35:0]   _zz_4756;
  wire       [35:0]   _zz_4757;
  wire       [35:0]   _zz_4758;
  wire       [26:0]   _zz_4759;
  wire       [35:0]   _zz_4760;
  wire       [17:0]   _zz_4761;
  wire       [35:0]   _zz_4762;
  wire       [35:0]   _zz_4763;
  wire       [35:0]   _zz_4764;
  wire       [35:0]   _zz_4765;
  wire       [35:0]   _zz_4766;
  wire       [26:0]   _zz_4767;
  wire       [35:0]   _zz_4768;
  wire       [17:0]   _zz_4769;
  wire       [35:0]   _zz_4770;
  wire       [35:0]   _zz_4771;
  wire       [35:0]   _zz_4772;
  wire       [35:0]   _zz_4773;
  wire       [35:0]   _zz_4774;
  wire       [26:0]   _zz_4775;
  wire       [35:0]   _zz_4776;
  wire       [17:0]   _zz_4777;
  wire       [17:0]   _zz_4778;
  wire       [35:0]   _zz_4779;
  wire       [35:0]   _zz_4780;
  wire       [17:0]   _zz_4781;
  wire       [35:0]   _zz_4782;
  wire       [35:0]   _zz_4783;
  wire       [35:0]   _zz_4784;
  wire       [17:0]   _zz_4785;
  wire       [35:0]   _zz_4786;
  wire       [35:0]   _zz_4787;
  wire       [35:0]   _zz_4788;
  wire       [35:0]   _zz_4789;
  wire       [35:0]   _zz_4790;
  wire       [35:0]   _zz_4791;
  wire       [26:0]   _zz_4792;
  wire       [35:0]   _zz_4793;
  wire       [17:0]   _zz_4794;
  wire       [35:0]   _zz_4795;
  wire       [35:0]   _zz_4796;
  wire       [35:0]   _zz_4797;
  wire       [35:0]   _zz_4798;
  wire       [35:0]   _zz_4799;
  wire       [26:0]   _zz_4800;
  wire       [35:0]   _zz_4801;
  wire       [17:0]   _zz_4802;
  wire       [35:0]   _zz_4803;
  wire       [35:0]   _zz_4804;
  wire       [35:0]   _zz_4805;
  wire       [35:0]   _zz_4806;
  wire       [35:0]   _zz_4807;
  wire       [26:0]   _zz_4808;
  wire       [35:0]   _zz_4809;
  wire       [17:0]   _zz_4810;
  wire       [35:0]   _zz_4811;
  wire       [35:0]   _zz_4812;
  wire       [35:0]   _zz_4813;
  wire       [35:0]   _zz_4814;
  wire       [35:0]   _zz_4815;
  wire       [26:0]   _zz_4816;
  wire       [35:0]   _zz_4817;
  wire       [17:0]   _zz_4818;
  wire       [17:0]   _zz_4819;
  wire       [35:0]   _zz_4820;
  wire       [35:0]   _zz_4821;
  wire       [17:0]   _zz_4822;
  wire       [35:0]   _zz_4823;
  wire       [35:0]   _zz_4824;
  wire       [35:0]   _zz_4825;
  wire       [17:0]   _zz_4826;
  wire       [35:0]   _zz_4827;
  wire       [35:0]   _zz_4828;
  wire       [35:0]   _zz_4829;
  wire       [35:0]   _zz_4830;
  wire       [35:0]   _zz_4831;
  wire       [35:0]   _zz_4832;
  wire       [26:0]   _zz_4833;
  wire       [35:0]   _zz_4834;
  wire       [17:0]   _zz_4835;
  wire       [35:0]   _zz_4836;
  wire       [35:0]   _zz_4837;
  wire       [35:0]   _zz_4838;
  wire       [35:0]   _zz_4839;
  wire       [35:0]   _zz_4840;
  wire       [26:0]   _zz_4841;
  wire       [35:0]   _zz_4842;
  wire       [17:0]   _zz_4843;
  wire       [35:0]   _zz_4844;
  wire       [35:0]   _zz_4845;
  wire       [35:0]   _zz_4846;
  wire       [35:0]   _zz_4847;
  wire       [35:0]   _zz_4848;
  wire       [26:0]   _zz_4849;
  wire       [35:0]   _zz_4850;
  wire       [17:0]   _zz_4851;
  wire       [35:0]   _zz_4852;
  wire       [35:0]   _zz_4853;
  wire       [35:0]   _zz_4854;
  wire       [35:0]   _zz_4855;
  wire       [35:0]   _zz_4856;
  wire       [26:0]   _zz_4857;
  wire       [35:0]   _zz_4858;
  wire       [17:0]   _zz_4859;
  wire       [17:0]   _zz_4860;
  wire       [35:0]   _zz_4861;
  wire       [35:0]   _zz_4862;
  wire       [17:0]   _zz_4863;
  wire       [35:0]   _zz_4864;
  wire       [35:0]   _zz_4865;
  wire       [35:0]   _zz_4866;
  wire       [17:0]   _zz_4867;
  wire       [35:0]   _zz_4868;
  wire       [35:0]   _zz_4869;
  wire       [35:0]   _zz_4870;
  wire       [35:0]   _zz_4871;
  wire       [35:0]   _zz_4872;
  wire       [35:0]   _zz_4873;
  wire       [26:0]   _zz_4874;
  wire       [35:0]   _zz_4875;
  wire       [17:0]   _zz_4876;
  wire       [35:0]   _zz_4877;
  wire       [35:0]   _zz_4878;
  wire       [35:0]   _zz_4879;
  wire       [35:0]   _zz_4880;
  wire       [35:0]   _zz_4881;
  wire       [26:0]   _zz_4882;
  wire       [35:0]   _zz_4883;
  wire       [17:0]   _zz_4884;
  wire       [35:0]   _zz_4885;
  wire       [35:0]   _zz_4886;
  wire       [35:0]   _zz_4887;
  wire       [35:0]   _zz_4888;
  wire       [35:0]   _zz_4889;
  wire       [26:0]   _zz_4890;
  wire       [35:0]   _zz_4891;
  wire       [17:0]   _zz_4892;
  wire       [35:0]   _zz_4893;
  wire       [35:0]   _zz_4894;
  wire       [35:0]   _zz_4895;
  wire       [35:0]   _zz_4896;
  wire       [35:0]   _zz_4897;
  wire       [26:0]   _zz_4898;
  wire       [35:0]   _zz_4899;
  wire       [17:0]   _zz_4900;
  wire       [17:0]   _zz_4901;
  wire       [35:0]   _zz_4902;
  wire       [35:0]   _zz_4903;
  wire       [17:0]   _zz_4904;
  wire       [35:0]   _zz_4905;
  wire       [35:0]   _zz_4906;
  wire       [35:0]   _zz_4907;
  wire       [17:0]   _zz_4908;
  wire       [35:0]   _zz_4909;
  wire       [35:0]   _zz_4910;
  wire       [35:0]   _zz_4911;
  wire       [35:0]   _zz_4912;
  wire       [35:0]   _zz_4913;
  wire       [35:0]   _zz_4914;
  wire       [26:0]   _zz_4915;
  wire       [35:0]   _zz_4916;
  wire       [17:0]   _zz_4917;
  wire       [35:0]   _zz_4918;
  wire       [35:0]   _zz_4919;
  wire       [35:0]   _zz_4920;
  wire       [35:0]   _zz_4921;
  wire       [35:0]   _zz_4922;
  wire       [26:0]   _zz_4923;
  wire       [35:0]   _zz_4924;
  wire       [17:0]   _zz_4925;
  wire       [35:0]   _zz_4926;
  wire       [35:0]   _zz_4927;
  wire       [35:0]   _zz_4928;
  wire       [35:0]   _zz_4929;
  wire       [35:0]   _zz_4930;
  wire       [26:0]   _zz_4931;
  wire       [35:0]   _zz_4932;
  wire       [17:0]   _zz_4933;
  wire       [35:0]   _zz_4934;
  wire       [35:0]   _zz_4935;
  wire       [35:0]   _zz_4936;
  wire       [35:0]   _zz_4937;
  wire       [35:0]   _zz_4938;
  wire       [26:0]   _zz_4939;
  wire       [35:0]   _zz_4940;
  wire       [17:0]   _zz_4941;
  wire       [17:0]   _zz_4942;
  wire       [35:0]   _zz_4943;
  wire       [35:0]   _zz_4944;
  wire       [17:0]   _zz_4945;
  wire       [35:0]   _zz_4946;
  wire       [35:0]   _zz_4947;
  wire       [35:0]   _zz_4948;
  wire       [17:0]   _zz_4949;
  wire       [35:0]   _zz_4950;
  wire       [35:0]   _zz_4951;
  wire       [35:0]   _zz_4952;
  wire       [35:0]   _zz_4953;
  wire       [35:0]   _zz_4954;
  wire       [35:0]   _zz_4955;
  wire       [26:0]   _zz_4956;
  wire       [35:0]   _zz_4957;
  wire       [17:0]   _zz_4958;
  wire       [35:0]   _zz_4959;
  wire       [35:0]   _zz_4960;
  wire       [35:0]   _zz_4961;
  wire       [35:0]   _zz_4962;
  wire       [35:0]   _zz_4963;
  wire       [26:0]   _zz_4964;
  wire       [35:0]   _zz_4965;
  wire       [17:0]   _zz_4966;
  wire       [35:0]   _zz_4967;
  wire       [35:0]   _zz_4968;
  wire       [35:0]   _zz_4969;
  wire       [35:0]   _zz_4970;
  wire       [35:0]   _zz_4971;
  wire       [26:0]   _zz_4972;
  wire       [35:0]   _zz_4973;
  wire       [17:0]   _zz_4974;
  wire       [35:0]   _zz_4975;
  wire       [35:0]   _zz_4976;
  wire       [35:0]   _zz_4977;
  wire       [35:0]   _zz_4978;
  wire       [35:0]   _zz_4979;
  wire       [26:0]   _zz_4980;
  wire       [35:0]   _zz_4981;
  wire       [17:0]   _zz_4982;
  wire       [17:0]   _zz_4983;
  wire       [35:0]   _zz_4984;
  wire       [35:0]   _zz_4985;
  wire       [17:0]   _zz_4986;
  wire       [35:0]   _zz_4987;
  wire       [35:0]   _zz_4988;
  wire       [35:0]   _zz_4989;
  wire       [17:0]   _zz_4990;
  wire       [35:0]   _zz_4991;
  wire       [35:0]   _zz_4992;
  wire       [35:0]   _zz_4993;
  wire       [35:0]   _zz_4994;
  wire       [35:0]   _zz_4995;
  wire       [35:0]   _zz_4996;
  wire       [26:0]   _zz_4997;
  wire       [35:0]   _zz_4998;
  wire       [17:0]   _zz_4999;
  wire       [35:0]   _zz_5000;
  wire       [35:0]   _zz_5001;
  wire       [35:0]   _zz_5002;
  wire       [35:0]   _zz_5003;
  wire       [35:0]   _zz_5004;
  wire       [26:0]   _zz_5005;
  wire       [35:0]   _zz_5006;
  wire       [17:0]   _zz_5007;
  wire       [35:0]   _zz_5008;
  wire       [35:0]   _zz_5009;
  wire       [35:0]   _zz_5010;
  wire       [35:0]   _zz_5011;
  wire       [35:0]   _zz_5012;
  wire       [26:0]   _zz_5013;
  wire       [35:0]   _zz_5014;
  wire       [17:0]   _zz_5015;
  wire       [35:0]   _zz_5016;
  wire       [35:0]   _zz_5017;
  wire       [35:0]   _zz_5018;
  wire       [35:0]   _zz_5019;
  wire       [35:0]   _zz_5020;
  wire       [26:0]   _zz_5021;
  wire       [35:0]   _zz_5022;
  wire       [17:0]   _zz_5023;
  wire       [17:0]   _zz_5024;
  wire       [35:0]   _zz_5025;
  wire       [35:0]   _zz_5026;
  wire       [17:0]   _zz_5027;
  wire       [35:0]   _zz_5028;
  wire       [35:0]   _zz_5029;
  wire       [35:0]   _zz_5030;
  wire       [17:0]   _zz_5031;
  wire       [35:0]   _zz_5032;
  wire       [35:0]   _zz_5033;
  wire       [35:0]   _zz_5034;
  wire       [35:0]   _zz_5035;
  wire       [35:0]   _zz_5036;
  wire       [35:0]   _zz_5037;
  wire       [26:0]   _zz_5038;
  wire       [35:0]   _zz_5039;
  wire       [17:0]   _zz_5040;
  wire       [35:0]   _zz_5041;
  wire       [35:0]   _zz_5042;
  wire       [35:0]   _zz_5043;
  wire       [35:0]   _zz_5044;
  wire       [35:0]   _zz_5045;
  wire       [26:0]   _zz_5046;
  wire       [35:0]   _zz_5047;
  wire       [17:0]   _zz_5048;
  wire       [35:0]   _zz_5049;
  wire       [35:0]   _zz_5050;
  wire       [35:0]   _zz_5051;
  wire       [35:0]   _zz_5052;
  wire       [35:0]   _zz_5053;
  wire       [26:0]   _zz_5054;
  wire       [35:0]   _zz_5055;
  wire       [17:0]   _zz_5056;
  wire       [35:0]   _zz_5057;
  wire       [35:0]   _zz_5058;
  wire       [35:0]   _zz_5059;
  wire       [35:0]   _zz_5060;
  wire       [35:0]   _zz_5061;
  wire       [26:0]   _zz_5062;
  wire       [35:0]   _zz_5063;
  wire       [17:0]   _zz_5064;
  wire       [17:0]   _zz_5065;
  wire       [35:0]   _zz_5066;
  wire       [35:0]   _zz_5067;
  wire       [17:0]   _zz_5068;
  wire       [35:0]   _zz_5069;
  wire       [35:0]   _zz_5070;
  wire       [35:0]   _zz_5071;
  wire       [17:0]   _zz_5072;
  wire       [35:0]   _zz_5073;
  wire       [35:0]   _zz_5074;
  wire       [35:0]   _zz_5075;
  wire       [35:0]   _zz_5076;
  wire       [35:0]   _zz_5077;
  wire       [35:0]   _zz_5078;
  wire       [26:0]   _zz_5079;
  wire       [35:0]   _zz_5080;
  wire       [17:0]   _zz_5081;
  wire       [35:0]   _zz_5082;
  wire       [35:0]   _zz_5083;
  wire       [35:0]   _zz_5084;
  wire       [35:0]   _zz_5085;
  wire       [35:0]   _zz_5086;
  wire       [26:0]   _zz_5087;
  wire       [35:0]   _zz_5088;
  wire       [17:0]   _zz_5089;
  wire       [35:0]   _zz_5090;
  wire       [35:0]   _zz_5091;
  wire       [35:0]   _zz_5092;
  wire       [35:0]   _zz_5093;
  wire       [35:0]   _zz_5094;
  wire       [26:0]   _zz_5095;
  wire       [35:0]   _zz_5096;
  wire       [17:0]   _zz_5097;
  wire       [35:0]   _zz_5098;
  wire       [35:0]   _zz_5099;
  wire       [35:0]   _zz_5100;
  wire       [35:0]   _zz_5101;
  wire       [35:0]   _zz_5102;
  wire       [26:0]   _zz_5103;
  wire       [35:0]   _zz_5104;
  wire       [17:0]   _zz_5105;
  wire       [17:0]   _zz_5106;
  wire       [35:0]   _zz_5107;
  wire       [35:0]   _zz_5108;
  wire       [17:0]   _zz_5109;
  wire       [35:0]   _zz_5110;
  wire       [35:0]   _zz_5111;
  wire       [35:0]   _zz_5112;
  wire       [17:0]   _zz_5113;
  wire       [35:0]   _zz_5114;
  wire       [35:0]   _zz_5115;
  wire       [35:0]   _zz_5116;
  wire       [35:0]   _zz_5117;
  wire       [35:0]   _zz_5118;
  wire       [35:0]   _zz_5119;
  wire       [26:0]   _zz_5120;
  wire       [35:0]   _zz_5121;
  wire       [17:0]   _zz_5122;
  wire       [35:0]   _zz_5123;
  wire       [35:0]   _zz_5124;
  wire       [35:0]   _zz_5125;
  wire       [35:0]   _zz_5126;
  wire       [35:0]   _zz_5127;
  wire       [26:0]   _zz_5128;
  wire       [35:0]   _zz_5129;
  wire       [17:0]   _zz_5130;
  wire       [35:0]   _zz_5131;
  wire       [35:0]   _zz_5132;
  wire       [35:0]   _zz_5133;
  wire       [35:0]   _zz_5134;
  wire       [35:0]   _zz_5135;
  wire       [26:0]   _zz_5136;
  wire       [35:0]   _zz_5137;
  wire       [17:0]   _zz_5138;
  wire       [35:0]   _zz_5139;
  wire       [35:0]   _zz_5140;
  wire       [35:0]   _zz_5141;
  wire       [35:0]   _zz_5142;
  wire       [35:0]   _zz_5143;
  wire       [26:0]   _zz_5144;
  wire       [35:0]   _zz_5145;
  wire       [17:0]   _zz_5146;
  wire       [17:0]   _zz_5147;
  wire       [35:0]   _zz_5148;
  wire       [35:0]   _zz_5149;
  wire       [17:0]   _zz_5150;
  wire       [35:0]   _zz_5151;
  wire       [35:0]   _zz_5152;
  wire       [35:0]   _zz_5153;
  wire       [17:0]   _zz_5154;
  wire       [35:0]   _zz_5155;
  wire       [35:0]   _zz_5156;
  wire       [35:0]   _zz_5157;
  wire       [35:0]   _zz_5158;
  wire       [35:0]   _zz_5159;
  wire       [35:0]   _zz_5160;
  wire       [26:0]   _zz_5161;
  wire       [35:0]   _zz_5162;
  wire       [17:0]   _zz_5163;
  wire       [35:0]   _zz_5164;
  wire       [35:0]   _zz_5165;
  wire       [35:0]   _zz_5166;
  wire       [35:0]   _zz_5167;
  wire       [35:0]   _zz_5168;
  wire       [26:0]   _zz_5169;
  wire       [35:0]   _zz_5170;
  wire       [17:0]   _zz_5171;
  wire       [35:0]   _zz_5172;
  wire       [35:0]   _zz_5173;
  wire       [35:0]   _zz_5174;
  wire       [35:0]   _zz_5175;
  wire       [35:0]   _zz_5176;
  wire       [26:0]   _zz_5177;
  wire       [35:0]   _zz_5178;
  wire       [17:0]   _zz_5179;
  wire       [35:0]   _zz_5180;
  wire       [35:0]   _zz_5181;
  wire       [35:0]   _zz_5182;
  wire       [35:0]   _zz_5183;
  wire       [35:0]   _zz_5184;
  wire       [26:0]   _zz_5185;
  wire       [35:0]   _zz_5186;
  wire       [17:0]   _zz_5187;
  wire       [17:0]   _zz_5188;
  wire       [35:0]   _zz_5189;
  wire       [35:0]   _zz_5190;
  wire       [17:0]   _zz_5191;
  wire       [35:0]   _zz_5192;
  wire       [35:0]   _zz_5193;
  wire       [35:0]   _zz_5194;
  wire       [17:0]   _zz_5195;
  wire       [35:0]   _zz_5196;
  wire       [35:0]   _zz_5197;
  wire       [35:0]   _zz_5198;
  wire       [35:0]   _zz_5199;
  wire       [35:0]   _zz_5200;
  wire       [35:0]   _zz_5201;
  wire       [26:0]   _zz_5202;
  wire       [35:0]   _zz_5203;
  wire       [17:0]   _zz_5204;
  wire       [35:0]   _zz_5205;
  wire       [35:0]   _zz_5206;
  wire       [35:0]   _zz_5207;
  wire       [35:0]   _zz_5208;
  wire       [35:0]   _zz_5209;
  wire       [26:0]   _zz_5210;
  wire       [35:0]   _zz_5211;
  wire       [17:0]   _zz_5212;
  wire       [35:0]   _zz_5213;
  wire       [35:0]   _zz_5214;
  wire       [35:0]   _zz_5215;
  wire       [35:0]   _zz_5216;
  wire       [35:0]   _zz_5217;
  wire       [26:0]   _zz_5218;
  wire       [35:0]   _zz_5219;
  wire       [17:0]   _zz_5220;
  wire       [35:0]   _zz_5221;
  wire       [35:0]   _zz_5222;
  wire       [35:0]   _zz_5223;
  wire       [35:0]   _zz_5224;
  wire       [35:0]   _zz_5225;
  wire       [26:0]   _zz_5226;
  wire       [35:0]   _zz_5227;
  wire       [17:0]   _zz_5228;
  wire       [17:0]   _zz_5229;
  wire       [35:0]   _zz_5230;
  wire       [35:0]   _zz_5231;
  wire       [17:0]   _zz_5232;
  wire       [35:0]   _zz_5233;
  wire       [35:0]   _zz_5234;
  wire       [35:0]   _zz_5235;
  wire       [17:0]   _zz_5236;
  wire       [35:0]   _zz_5237;
  wire       [35:0]   _zz_5238;
  wire       [35:0]   _zz_5239;
  wire       [35:0]   _zz_5240;
  wire       [35:0]   _zz_5241;
  wire       [35:0]   _zz_5242;
  wire       [26:0]   _zz_5243;
  wire       [35:0]   _zz_5244;
  wire       [17:0]   _zz_5245;
  wire       [35:0]   _zz_5246;
  wire       [35:0]   _zz_5247;
  wire       [35:0]   _zz_5248;
  wire       [35:0]   _zz_5249;
  wire       [35:0]   _zz_5250;
  wire       [26:0]   _zz_5251;
  wire       [35:0]   _zz_5252;
  wire       [17:0]   _zz_5253;
  wire       [35:0]   _zz_5254;
  wire       [35:0]   _zz_5255;
  wire       [35:0]   _zz_5256;
  wire       [35:0]   _zz_5257;
  wire       [35:0]   _zz_5258;
  wire       [26:0]   _zz_5259;
  wire       [35:0]   _zz_5260;
  wire       [17:0]   _zz_5261;
  wire       [35:0]   _zz_5262;
  wire       [35:0]   _zz_5263;
  wire       [35:0]   _zz_5264;
  wire       [35:0]   _zz_5265;
  wire       [35:0]   _zz_5266;
  wire       [26:0]   _zz_5267;
  wire       [35:0]   _zz_5268;
  wire       [17:0]   _zz_5269;
  wire       [17:0]   _zz_5270;
  wire       [35:0]   _zz_5271;
  wire       [35:0]   _zz_5272;
  wire       [17:0]   _zz_5273;
  wire       [35:0]   _zz_5274;
  wire       [35:0]   _zz_5275;
  wire       [35:0]   _zz_5276;
  wire       [17:0]   _zz_5277;
  wire       [35:0]   _zz_5278;
  wire       [35:0]   _zz_5279;
  wire       [35:0]   _zz_5280;
  wire       [35:0]   _zz_5281;
  wire       [35:0]   _zz_5282;
  wire       [35:0]   _zz_5283;
  wire       [26:0]   _zz_5284;
  wire       [35:0]   _zz_5285;
  wire       [17:0]   _zz_5286;
  wire       [35:0]   _zz_5287;
  wire       [35:0]   _zz_5288;
  wire       [35:0]   _zz_5289;
  wire       [35:0]   _zz_5290;
  wire       [35:0]   _zz_5291;
  wire       [26:0]   _zz_5292;
  wire       [35:0]   _zz_5293;
  wire       [17:0]   _zz_5294;
  wire       [35:0]   _zz_5295;
  wire       [35:0]   _zz_5296;
  wire       [35:0]   _zz_5297;
  wire       [35:0]   _zz_5298;
  wire       [35:0]   _zz_5299;
  wire       [26:0]   _zz_5300;
  wire       [35:0]   _zz_5301;
  wire       [17:0]   _zz_5302;
  wire       [35:0]   _zz_5303;
  wire       [35:0]   _zz_5304;
  wire       [35:0]   _zz_5305;
  wire       [35:0]   _zz_5306;
  wire       [35:0]   _zz_5307;
  wire       [26:0]   _zz_5308;
  wire       [35:0]   _zz_5309;
  wire       [17:0]   _zz_5310;
  wire       [17:0]   _zz_5311;
  wire       [35:0]   _zz_5312;
  wire       [35:0]   _zz_5313;
  wire       [17:0]   _zz_5314;
  wire       [35:0]   _zz_5315;
  wire       [35:0]   _zz_5316;
  wire       [35:0]   _zz_5317;
  wire       [17:0]   _zz_5318;
  wire       [35:0]   _zz_5319;
  wire       [35:0]   _zz_5320;
  wire       [35:0]   _zz_5321;
  wire       [35:0]   _zz_5322;
  wire       [35:0]   _zz_5323;
  wire       [35:0]   _zz_5324;
  wire       [26:0]   _zz_5325;
  wire       [35:0]   _zz_5326;
  wire       [17:0]   _zz_5327;
  wire       [35:0]   _zz_5328;
  wire       [35:0]   _zz_5329;
  wire       [35:0]   _zz_5330;
  wire       [35:0]   _zz_5331;
  wire       [35:0]   _zz_5332;
  wire       [26:0]   _zz_5333;
  wire       [35:0]   _zz_5334;
  wire       [17:0]   _zz_5335;
  wire       [35:0]   _zz_5336;
  wire       [35:0]   _zz_5337;
  wire       [35:0]   _zz_5338;
  wire       [35:0]   _zz_5339;
  wire       [35:0]   _zz_5340;
  wire       [26:0]   _zz_5341;
  wire       [35:0]   _zz_5342;
  wire       [17:0]   _zz_5343;
  wire       [35:0]   _zz_5344;
  wire       [35:0]   _zz_5345;
  wire       [35:0]   _zz_5346;
  wire       [35:0]   _zz_5347;
  wire       [35:0]   _zz_5348;
  wire       [26:0]   _zz_5349;
  wire       [35:0]   _zz_5350;
  wire       [17:0]   _zz_5351;
  wire       [17:0]   _zz_5352;
  wire       [35:0]   _zz_5353;
  wire       [35:0]   _zz_5354;
  wire       [17:0]   _zz_5355;
  wire       [35:0]   _zz_5356;
  wire       [35:0]   _zz_5357;
  wire       [35:0]   _zz_5358;
  wire       [17:0]   _zz_5359;
  wire       [35:0]   _zz_5360;
  wire       [35:0]   _zz_5361;
  wire       [35:0]   _zz_5362;
  wire       [35:0]   _zz_5363;
  wire       [35:0]   _zz_5364;
  wire       [35:0]   _zz_5365;
  wire       [26:0]   _zz_5366;
  wire       [35:0]   _zz_5367;
  wire       [17:0]   _zz_5368;
  wire       [35:0]   _zz_5369;
  wire       [35:0]   _zz_5370;
  wire       [35:0]   _zz_5371;
  wire       [35:0]   _zz_5372;
  wire       [35:0]   _zz_5373;
  wire       [26:0]   _zz_5374;
  wire       [35:0]   _zz_5375;
  wire       [17:0]   _zz_5376;
  wire       [35:0]   _zz_5377;
  wire       [35:0]   _zz_5378;
  wire       [35:0]   _zz_5379;
  wire       [35:0]   _zz_5380;
  wire       [35:0]   _zz_5381;
  wire       [26:0]   _zz_5382;
  wire       [35:0]   _zz_5383;
  wire       [17:0]   _zz_5384;
  wire       [35:0]   _zz_5385;
  wire       [35:0]   _zz_5386;
  wire       [35:0]   _zz_5387;
  wire       [35:0]   _zz_5388;
  wire       [35:0]   _zz_5389;
  wire       [26:0]   _zz_5390;
  wire       [35:0]   _zz_5391;
  wire       [17:0]   _zz_5392;
  wire       [17:0]   _zz_5393;
  wire       [35:0]   _zz_5394;
  wire       [35:0]   _zz_5395;
  wire       [17:0]   _zz_5396;
  wire       [35:0]   _zz_5397;
  wire       [35:0]   _zz_5398;
  wire       [35:0]   _zz_5399;
  wire       [17:0]   _zz_5400;
  wire       [35:0]   _zz_5401;
  wire       [35:0]   _zz_5402;
  wire       [35:0]   _zz_5403;
  wire       [35:0]   _zz_5404;
  wire       [35:0]   _zz_5405;
  wire       [35:0]   _zz_5406;
  wire       [26:0]   _zz_5407;
  wire       [35:0]   _zz_5408;
  wire       [17:0]   _zz_5409;
  wire       [35:0]   _zz_5410;
  wire       [35:0]   _zz_5411;
  wire       [35:0]   _zz_5412;
  wire       [35:0]   _zz_5413;
  wire       [35:0]   _zz_5414;
  wire       [26:0]   _zz_5415;
  wire       [35:0]   _zz_5416;
  wire       [17:0]   _zz_5417;
  wire       [35:0]   _zz_5418;
  wire       [35:0]   _zz_5419;
  wire       [35:0]   _zz_5420;
  wire       [35:0]   _zz_5421;
  wire       [35:0]   _zz_5422;
  wire       [26:0]   _zz_5423;
  wire       [35:0]   _zz_5424;
  wire       [17:0]   _zz_5425;
  wire       [35:0]   _zz_5426;
  wire       [35:0]   _zz_5427;
  wire       [35:0]   _zz_5428;
  wire       [35:0]   _zz_5429;
  wire       [35:0]   _zz_5430;
  wire       [26:0]   _zz_5431;
  wire       [35:0]   _zz_5432;
  wire       [17:0]   _zz_5433;
  wire       [17:0]   _zz_5434;
  wire       [35:0]   _zz_5435;
  wire       [35:0]   _zz_5436;
  wire       [17:0]   _zz_5437;
  wire       [35:0]   _zz_5438;
  wire       [35:0]   _zz_5439;
  wire       [35:0]   _zz_5440;
  wire       [17:0]   _zz_5441;
  wire       [35:0]   _zz_5442;
  wire       [35:0]   _zz_5443;
  wire       [35:0]   _zz_5444;
  wire       [35:0]   _zz_5445;
  wire       [35:0]   _zz_5446;
  wire       [35:0]   _zz_5447;
  wire       [26:0]   _zz_5448;
  wire       [35:0]   _zz_5449;
  wire       [17:0]   _zz_5450;
  wire       [35:0]   _zz_5451;
  wire       [35:0]   _zz_5452;
  wire       [35:0]   _zz_5453;
  wire       [35:0]   _zz_5454;
  wire       [35:0]   _zz_5455;
  wire       [26:0]   _zz_5456;
  wire       [35:0]   _zz_5457;
  wire       [17:0]   _zz_5458;
  wire       [35:0]   _zz_5459;
  wire       [35:0]   _zz_5460;
  wire       [35:0]   _zz_5461;
  wire       [35:0]   _zz_5462;
  wire       [35:0]   _zz_5463;
  wire       [26:0]   _zz_5464;
  wire       [35:0]   _zz_5465;
  wire       [17:0]   _zz_5466;
  wire       [35:0]   _zz_5467;
  wire       [35:0]   _zz_5468;
  wire       [35:0]   _zz_5469;
  wire       [35:0]   _zz_5470;
  wire       [35:0]   _zz_5471;
  wire       [26:0]   _zz_5472;
  wire       [35:0]   _zz_5473;
  wire       [17:0]   _zz_5474;
  wire       [17:0]   _zz_5475;
  wire       [35:0]   _zz_5476;
  wire       [35:0]   _zz_5477;
  wire       [17:0]   _zz_5478;
  wire       [35:0]   _zz_5479;
  wire       [35:0]   _zz_5480;
  wire       [35:0]   _zz_5481;
  wire       [17:0]   _zz_5482;
  wire       [35:0]   _zz_5483;
  wire       [35:0]   _zz_5484;
  wire       [35:0]   _zz_5485;
  wire       [35:0]   _zz_5486;
  wire       [35:0]   _zz_5487;
  wire       [35:0]   _zz_5488;
  wire       [26:0]   _zz_5489;
  wire       [35:0]   _zz_5490;
  wire       [17:0]   _zz_5491;
  wire       [35:0]   _zz_5492;
  wire       [35:0]   _zz_5493;
  wire       [35:0]   _zz_5494;
  wire       [35:0]   _zz_5495;
  wire       [35:0]   _zz_5496;
  wire       [26:0]   _zz_5497;
  wire       [35:0]   _zz_5498;
  wire       [17:0]   _zz_5499;
  wire       [35:0]   _zz_5500;
  wire       [35:0]   _zz_5501;
  wire       [35:0]   _zz_5502;
  wire       [35:0]   _zz_5503;
  wire       [35:0]   _zz_5504;
  wire       [26:0]   _zz_5505;
  wire       [35:0]   _zz_5506;
  wire       [17:0]   _zz_5507;
  wire       [35:0]   _zz_5508;
  wire       [35:0]   _zz_5509;
  wire       [35:0]   _zz_5510;
  wire       [35:0]   _zz_5511;
  wire       [35:0]   _zz_5512;
  wire       [26:0]   _zz_5513;
  wire       [35:0]   _zz_5514;
  wire       [17:0]   _zz_5515;
  wire       [17:0]   _zz_5516;
  wire       [35:0]   _zz_5517;
  wire       [35:0]   _zz_5518;
  wire       [17:0]   _zz_5519;
  wire       [35:0]   _zz_5520;
  wire       [35:0]   _zz_5521;
  wire       [35:0]   _zz_5522;
  wire       [17:0]   _zz_5523;
  wire       [35:0]   _zz_5524;
  wire       [35:0]   _zz_5525;
  wire       [35:0]   _zz_5526;
  wire       [35:0]   _zz_5527;
  wire       [35:0]   _zz_5528;
  wire       [35:0]   _zz_5529;
  wire       [26:0]   _zz_5530;
  wire       [35:0]   _zz_5531;
  wire       [17:0]   _zz_5532;
  wire       [35:0]   _zz_5533;
  wire       [35:0]   _zz_5534;
  wire       [35:0]   _zz_5535;
  wire       [35:0]   _zz_5536;
  wire       [35:0]   _zz_5537;
  wire       [26:0]   _zz_5538;
  wire       [35:0]   _zz_5539;
  wire       [17:0]   _zz_5540;
  wire       [35:0]   _zz_5541;
  wire       [35:0]   _zz_5542;
  wire       [35:0]   _zz_5543;
  wire       [35:0]   _zz_5544;
  wire       [35:0]   _zz_5545;
  wire       [26:0]   _zz_5546;
  wire       [35:0]   _zz_5547;
  wire       [17:0]   _zz_5548;
  wire       [35:0]   _zz_5549;
  wire       [35:0]   _zz_5550;
  wire       [35:0]   _zz_5551;
  wire       [35:0]   _zz_5552;
  wire       [35:0]   _zz_5553;
  wire       [26:0]   _zz_5554;
  wire       [35:0]   _zz_5555;
  wire       [17:0]   _zz_5556;
  wire       [17:0]   _zz_5557;
  wire       [35:0]   _zz_5558;
  wire       [35:0]   _zz_5559;
  wire       [17:0]   _zz_5560;
  wire       [35:0]   _zz_5561;
  wire       [35:0]   _zz_5562;
  wire       [35:0]   _zz_5563;
  wire       [17:0]   _zz_5564;
  wire       [35:0]   _zz_5565;
  wire       [35:0]   _zz_5566;
  wire       [35:0]   _zz_5567;
  wire       [35:0]   _zz_5568;
  wire       [35:0]   _zz_5569;
  wire       [35:0]   _zz_5570;
  wire       [26:0]   _zz_5571;
  wire       [35:0]   _zz_5572;
  wire       [17:0]   _zz_5573;
  wire       [35:0]   _zz_5574;
  wire       [35:0]   _zz_5575;
  wire       [35:0]   _zz_5576;
  wire       [35:0]   _zz_5577;
  wire       [35:0]   _zz_5578;
  wire       [26:0]   _zz_5579;
  wire       [35:0]   _zz_5580;
  wire       [17:0]   _zz_5581;
  wire       [35:0]   _zz_5582;
  wire       [35:0]   _zz_5583;
  wire       [35:0]   _zz_5584;
  wire       [35:0]   _zz_5585;
  wire       [35:0]   _zz_5586;
  wire       [26:0]   _zz_5587;
  wire       [35:0]   _zz_5588;
  wire       [17:0]   _zz_5589;
  wire       [35:0]   _zz_5590;
  wire       [35:0]   _zz_5591;
  wire       [35:0]   _zz_5592;
  wire       [35:0]   _zz_5593;
  wire       [35:0]   _zz_5594;
  wire       [26:0]   _zz_5595;
  wire       [35:0]   _zz_5596;
  wire       [17:0]   _zz_5597;
  wire       [17:0]   _zz_5598;
  wire       [35:0]   _zz_5599;
  wire       [35:0]   _zz_5600;
  wire       [17:0]   _zz_5601;
  wire       [35:0]   _zz_5602;
  wire       [35:0]   _zz_5603;
  wire       [35:0]   _zz_5604;
  wire       [17:0]   _zz_5605;
  wire       [35:0]   _zz_5606;
  wire       [35:0]   _zz_5607;
  wire       [35:0]   _zz_5608;
  wire       [35:0]   _zz_5609;
  wire       [35:0]   _zz_5610;
  wire       [35:0]   _zz_5611;
  wire       [26:0]   _zz_5612;
  wire       [35:0]   _zz_5613;
  wire       [17:0]   _zz_5614;
  wire       [35:0]   _zz_5615;
  wire       [35:0]   _zz_5616;
  wire       [35:0]   _zz_5617;
  wire       [35:0]   _zz_5618;
  wire       [35:0]   _zz_5619;
  wire       [26:0]   _zz_5620;
  wire       [35:0]   _zz_5621;
  wire       [17:0]   _zz_5622;
  wire       [35:0]   _zz_5623;
  wire       [35:0]   _zz_5624;
  wire       [35:0]   _zz_5625;
  wire       [35:0]   _zz_5626;
  wire       [35:0]   _zz_5627;
  wire       [26:0]   _zz_5628;
  wire       [35:0]   _zz_5629;
  wire       [17:0]   _zz_5630;
  wire       [35:0]   _zz_5631;
  wire       [35:0]   _zz_5632;
  wire       [35:0]   _zz_5633;
  wire       [35:0]   _zz_5634;
  wire       [35:0]   _zz_5635;
  wire       [26:0]   _zz_5636;
  wire       [35:0]   _zz_5637;
  wire       [17:0]   _zz_5638;
  wire       [17:0]   _zz_5639;
  wire       [35:0]   _zz_5640;
  wire       [35:0]   _zz_5641;
  wire       [17:0]   _zz_5642;
  wire       [35:0]   _zz_5643;
  wire       [35:0]   _zz_5644;
  wire       [35:0]   _zz_5645;
  wire       [17:0]   _zz_5646;
  wire       [35:0]   _zz_5647;
  wire       [35:0]   _zz_5648;
  wire       [35:0]   _zz_5649;
  wire       [35:0]   _zz_5650;
  wire       [35:0]   _zz_5651;
  wire       [35:0]   _zz_5652;
  wire       [26:0]   _zz_5653;
  wire       [35:0]   _zz_5654;
  wire       [17:0]   _zz_5655;
  wire       [35:0]   _zz_5656;
  wire       [35:0]   _zz_5657;
  wire       [35:0]   _zz_5658;
  wire       [35:0]   _zz_5659;
  wire       [35:0]   _zz_5660;
  wire       [26:0]   _zz_5661;
  wire       [35:0]   _zz_5662;
  wire       [17:0]   _zz_5663;
  wire       [35:0]   _zz_5664;
  wire       [35:0]   _zz_5665;
  wire       [35:0]   _zz_5666;
  wire       [35:0]   _zz_5667;
  wire       [35:0]   _zz_5668;
  wire       [26:0]   _zz_5669;
  wire       [35:0]   _zz_5670;
  wire       [17:0]   _zz_5671;
  wire       [35:0]   _zz_5672;
  wire       [35:0]   _zz_5673;
  wire       [35:0]   _zz_5674;
  wire       [35:0]   _zz_5675;
  wire       [35:0]   _zz_5676;
  wire       [26:0]   _zz_5677;
  wire       [35:0]   _zz_5678;
  wire       [17:0]   _zz_5679;
  wire       [17:0]   _zz_5680;
  wire       [35:0]   _zz_5681;
  wire       [35:0]   _zz_5682;
  wire       [17:0]   _zz_5683;
  wire       [35:0]   _zz_5684;
  wire       [35:0]   _zz_5685;
  wire       [35:0]   _zz_5686;
  wire       [17:0]   _zz_5687;
  wire       [35:0]   _zz_5688;
  wire       [35:0]   _zz_5689;
  wire       [35:0]   _zz_5690;
  wire       [35:0]   _zz_5691;
  wire       [35:0]   _zz_5692;
  wire       [35:0]   _zz_5693;
  wire       [26:0]   _zz_5694;
  wire       [35:0]   _zz_5695;
  wire       [17:0]   _zz_5696;
  wire       [35:0]   _zz_5697;
  wire       [35:0]   _zz_5698;
  wire       [35:0]   _zz_5699;
  wire       [35:0]   _zz_5700;
  wire       [35:0]   _zz_5701;
  wire       [26:0]   _zz_5702;
  wire       [35:0]   _zz_5703;
  wire       [17:0]   _zz_5704;
  wire       [35:0]   _zz_5705;
  wire       [35:0]   _zz_5706;
  wire       [35:0]   _zz_5707;
  wire       [35:0]   _zz_5708;
  wire       [35:0]   _zz_5709;
  wire       [26:0]   _zz_5710;
  wire       [35:0]   _zz_5711;
  wire       [17:0]   _zz_5712;
  wire       [35:0]   _zz_5713;
  wire       [35:0]   _zz_5714;
  wire       [35:0]   _zz_5715;
  wire       [35:0]   _zz_5716;
  wire       [35:0]   _zz_5717;
  wire       [26:0]   _zz_5718;
  wire       [35:0]   _zz_5719;
  wire       [17:0]   _zz_5720;
  wire       [17:0]   _zz_5721;
  wire       [35:0]   _zz_5722;
  wire       [35:0]   _zz_5723;
  wire       [17:0]   _zz_5724;
  wire       [35:0]   _zz_5725;
  wire       [35:0]   _zz_5726;
  wire       [35:0]   _zz_5727;
  wire       [17:0]   _zz_5728;
  wire       [35:0]   _zz_5729;
  wire       [35:0]   _zz_5730;
  wire       [35:0]   _zz_5731;
  wire       [35:0]   _zz_5732;
  wire       [35:0]   _zz_5733;
  wire       [35:0]   _zz_5734;
  wire       [26:0]   _zz_5735;
  wire       [35:0]   _zz_5736;
  wire       [17:0]   _zz_5737;
  wire       [35:0]   _zz_5738;
  wire       [35:0]   _zz_5739;
  wire       [35:0]   _zz_5740;
  wire       [35:0]   _zz_5741;
  wire       [35:0]   _zz_5742;
  wire       [26:0]   _zz_5743;
  wire       [35:0]   _zz_5744;
  wire       [17:0]   _zz_5745;
  wire       [35:0]   _zz_5746;
  wire       [35:0]   _zz_5747;
  wire       [35:0]   _zz_5748;
  wire       [35:0]   _zz_5749;
  wire       [35:0]   _zz_5750;
  wire       [26:0]   _zz_5751;
  wire       [35:0]   _zz_5752;
  wire       [17:0]   _zz_5753;
  wire       [35:0]   _zz_5754;
  wire       [35:0]   _zz_5755;
  wire       [35:0]   _zz_5756;
  wire       [35:0]   _zz_5757;
  wire       [35:0]   _zz_5758;
  wire       [26:0]   _zz_5759;
  wire       [35:0]   _zz_5760;
  wire       [17:0]   _zz_5761;
  wire       [17:0]   _zz_5762;
  wire       [35:0]   _zz_5763;
  wire       [35:0]   _zz_5764;
  wire       [17:0]   _zz_5765;
  wire       [35:0]   _zz_5766;
  wire       [35:0]   _zz_5767;
  wire       [35:0]   _zz_5768;
  wire       [17:0]   _zz_5769;
  wire       [35:0]   _zz_5770;
  wire       [35:0]   _zz_5771;
  wire       [35:0]   _zz_5772;
  wire       [35:0]   _zz_5773;
  wire       [35:0]   _zz_5774;
  wire       [35:0]   _zz_5775;
  wire       [26:0]   _zz_5776;
  wire       [35:0]   _zz_5777;
  wire       [17:0]   _zz_5778;
  wire       [35:0]   _zz_5779;
  wire       [35:0]   _zz_5780;
  wire       [35:0]   _zz_5781;
  wire       [35:0]   _zz_5782;
  wire       [35:0]   _zz_5783;
  wire       [26:0]   _zz_5784;
  wire       [35:0]   _zz_5785;
  wire       [17:0]   _zz_5786;
  wire       [35:0]   _zz_5787;
  wire       [35:0]   _zz_5788;
  wire       [35:0]   _zz_5789;
  wire       [35:0]   _zz_5790;
  wire       [35:0]   _zz_5791;
  wire       [26:0]   _zz_5792;
  wire       [35:0]   _zz_5793;
  wire       [17:0]   _zz_5794;
  wire       [35:0]   _zz_5795;
  wire       [35:0]   _zz_5796;
  wire       [35:0]   _zz_5797;
  wire       [35:0]   _zz_5798;
  wire       [35:0]   _zz_5799;
  wire       [26:0]   _zz_5800;
  wire       [35:0]   _zz_5801;
  wire       [17:0]   _zz_5802;
  wire       [17:0]   _zz_5803;
  wire       [35:0]   _zz_5804;
  wire       [35:0]   _zz_5805;
  wire       [17:0]   _zz_5806;
  wire       [35:0]   _zz_5807;
  wire       [35:0]   _zz_5808;
  wire       [35:0]   _zz_5809;
  wire       [17:0]   _zz_5810;
  wire       [35:0]   _zz_5811;
  wire       [35:0]   _zz_5812;
  wire       [35:0]   _zz_5813;
  wire       [35:0]   _zz_5814;
  wire       [35:0]   _zz_5815;
  wire       [35:0]   _zz_5816;
  wire       [26:0]   _zz_5817;
  wire       [35:0]   _zz_5818;
  wire       [17:0]   _zz_5819;
  wire       [35:0]   _zz_5820;
  wire       [35:0]   _zz_5821;
  wire       [35:0]   _zz_5822;
  wire       [35:0]   _zz_5823;
  wire       [35:0]   _zz_5824;
  wire       [26:0]   _zz_5825;
  wire       [35:0]   _zz_5826;
  wire       [17:0]   _zz_5827;
  wire       [35:0]   _zz_5828;
  wire       [35:0]   _zz_5829;
  wire       [35:0]   _zz_5830;
  wire       [35:0]   _zz_5831;
  wire       [35:0]   _zz_5832;
  wire       [26:0]   _zz_5833;
  wire       [35:0]   _zz_5834;
  wire       [17:0]   _zz_5835;
  wire       [35:0]   _zz_5836;
  wire       [35:0]   _zz_5837;
  wire       [35:0]   _zz_5838;
  wire       [35:0]   _zz_5839;
  wire       [35:0]   _zz_5840;
  wire       [26:0]   _zz_5841;
  wire       [35:0]   _zz_5842;
  wire       [17:0]   _zz_5843;
  wire       [17:0]   _zz_5844;
  wire       [35:0]   _zz_5845;
  wire       [35:0]   _zz_5846;
  wire       [17:0]   _zz_5847;
  wire       [35:0]   _zz_5848;
  wire       [35:0]   _zz_5849;
  wire       [35:0]   _zz_5850;
  wire       [17:0]   _zz_5851;
  wire       [35:0]   _zz_5852;
  wire       [35:0]   _zz_5853;
  wire       [35:0]   _zz_5854;
  wire       [35:0]   _zz_5855;
  wire       [35:0]   _zz_5856;
  wire       [35:0]   _zz_5857;
  wire       [26:0]   _zz_5858;
  wire       [35:0]   _zz_5859;
  wire       [17:0]   _zz_5860;
  wire       [35:0]   _zz_5861;
  wire       [35:0]   _zz_5862;
  wire       [35:0]   _zz_5863;
  wire       [35:0]   _zz_5864;
  wire       [35:0]   _zz_5865;
  wire       [26:0]   _zz_5866;
  wire       [35:0]   _zz_5867;
  wire       [17:0]   _zz_5868;
  wire       [35:0]   _zz_5869;
  wire       [35:0]   _zz_5870;
  wire       [35:0]   _zz_5871;
  wire       [35:0]   _zz_5872;
  wire       [35:0]   _zz_5873;
  wire       [26:0]   _zz_5874;
  wire       [35:0]   _zz_5875;
  wire       [17:0]   _zz_5876;
  wire       [35:0]   _zz_5877;
  wire       [35:0]   _zz_5878;
  wire       [35:0]   _zz_5879;
  wire       [35:0]   _zz_5880;
  wire       [35:0]   _zz_5881;
  wire       [26:0]   _zz_5882;
  wire       [35:0]   _zz_5883;
  wire       [17:0]   _zz_5884;
  wire       [17:0]   _zz_5885;
  wire       [35:0]   _zz_5886;
  wire       [35:0]   _zz_5887;
  wire       [17:0]   _zz_5888;
  wire       [35:0]   _zz_5889;
  wire       [35:0]   _zz_5890;
  wire       [35:0]   _zz_5891;
  wire       [17:0]   _zz_5892;
  wire       [35:0]   _zz_5893;
  wire       [35:0]   _zz_5894;
  wire       [35:0]   _zz_5895;
  wire       [35:0]   _zz_5896;
  wire       [35:0]   _zz_5897;
  wire       [35:0]   _zz_5898;
  wire       [26:0]   _zz_5899;
  wire       [35:0]   _zz_5900;
  wire       [17:0]   _zz_5901;
  wire       [35:0]   _zz_5902;
  wire       [35:0]   _zz_5903;
  wire       [35:0]   _zz_5904;
  wire       [35:0]   _zz_5905;
  wire       [35:0]   _zz_5906;
  wire       [26:0]   _zz_5907;
  wire       [35:0]   _zz_5908;
  wire       [17:0]   _zz_5909;
  wire       [35:0]   _zz_5910;
  wire       [35:0]   _zz_5911;
  wire       [35:0]   _zz_5912;
  wire       [35:0]   _zz_5913;
  wire       [35:0]   _zz_5914;
  wire       [26:0]   _zz_5915;
  wire       [35:0]   _zz_5916;
  wire       [17:0]   _zz_5917;
  wire       [35:0]   _zz_5918;
  wire       [35:0]   _zz_5919;
  wire       [35:0]   _zz_5920;
  wire       [35:0]   _zz_5921;
  wire       [35:0]   _zz_5922;
  wire       [26:0]   _zz_5923;
  wire       [35:0]   _zz_5924;
  wire       [17:0]   _zz_5925;
  wire       [17:0]   _zz_5926;
  wire       [35:0]   _zz_5927;
  wire       [35:0]   _zz_5928;
  wire       [17:0]   _zz_5929;
  wire       [35:0]   _zz_5930;
  wire       [35:0]   _zz_5931;
  wire       [35:0]   _zz_5932;
  wire       [17:0]   _zz_5933;
  wire       [35:0]   _zz_5934;
  wire       [35:0]   _zz_5935;
  wire       [35:0]   _zz_5936;
  wire       [35:0]   _zz_5937;
  wire       [35:0]   _zz_5938;
  wire       [35:0]   _zz_5939;
  wire       [26:0]   _zz_5940;
  wire       [35:0]   _zz_5941;
  wire       [17:0]   _zz_5942;
  wire       [35:0]   _zz_5943;
  wire       [35:0]   _zz_5944;
  wire       [35:0]   _zz_5945;
  wire       [35:0]   _zz_5946;
  wire       [35:0]   _zz_5947;
  wire       [26:0]   _zz_5948;
  wire       [35:0]   _zz_5949;
  wire       [17:0]   _zz_5950;
  wire       [35:0]   _zz_5951;
  wire       [35:0]   _zz_5952;
  wire       [35:0]   _zz_5953;
  wire       [35:0]   _zz_5954;
  wire       [35:0]   _zz_5955;
  wire       [26:0]   _zz_5956;
  wire       [35:0]   _zz_5957;
  wire       [17:0]   _zz_5958;
  wire       [35:0]   _zz_5959;
  wire       [35:0]   _zz_5960;
  wire       [35:0]   _zz_5961;
  wire       [35:0]   _zz_5962;
  wire       [35:0]   _zz_5963;
  wire       [26:0]   _zz_5964;
  wire       [35:0]   _zz_5965;
  wire       [17:0]   _zz_5966;
  wire       [17:0]   _zz_5967;
  wire       [35:0]   _zz_5968;
  wire       [35:0]   _zz_5969;
  wire       [17:0]   _zz_5970;
  wire       [35:0]   _zz_5971;
  wire       [35:0]   _zz_5972;
  wire       [35:0]   _zz_5973;
  wire       [17:0]   _zz_5974;
  wire       [35:0]   _zz_5975;
  wire       [35:0]   _zz_5976;
  wire       [35:0]   _zz_5977;
  wire       [35:0]   _zz_5978;
  wire       [35:0]   _zz_5979;
  wire       [35:0]   _zz_5980;
  wire       [26:0]   _zz_5981;
  wire       [35:0]   _zz_5982;
  wire       [17:0]   _zz_5983;
  wire       [35:0]   _zz_5984;
  wire       [35:0]   _zz_5985;
  wire       [35:0]   _zz_5986;
  wire       [35:0]   _zz_5987;
  wire       [35:0]   _zz_5988;
  wire       [26:0]   _zz_5989;
  wire       [35:0]   _zz_5990;
  wire       [17:0]   _zz_5991;
  wire       [35:0]   _zz_5992;
  wire       [35:0]   _zz_5993;
  wire       [35:0]   _zz_5994;
  wire       [35:0]   _zz_5995;
  wire       [35:0]   _zz_5996;
  wire       [26:0]   _zz_5997;
  wire       [35:0]   _zz_5998;
  wire       [17:0]   _zz_5999;
  wire       [35:0]   _zz_6000;
  wire       [35:0]   _zz_6001;
  wire       [35:0]   _zz_6002;
  wire       [35:0]   _zz_6003;
  wire       [35:0]   _zz_6004;
  wire       [26:0]   _zz_6005;
  wire       [35:0]   _zz_6006;
  wire       [17:0]   _zz_6007;
  wire       [17:0]   _zz_6008;
  wire       [35:0]   _zz_6009;
  wire       [35:0]   _zz_6010;
  wire       [17:0]   _zz_6011;
  wire       [35:0]   _zz_6012;
  wire       [35:0]   _zz_6013;
  wire       [35:0]   _zz_6014;
  wire       [17:0]   _zz_6015;
  wire       [35:0]   _zz_6016;
  wire       [35:0]   _zz_6017;
  wire       [35:0]   _zz_6018;
  wire       [35:0]   _zz_6019;
  wire       [35:0]   _zz_6020;
  wire       [35:0]   _zz_6021;
  wire       [26:0]   _zz_6022;
  wire       [35:0]   _zz_6023;
  wire       [17:0]   _zz_6024;
  wire       [35:0]   _zz_6025;
  wire       [35:0]   _zz_6026;
  wire       [35:0]   _zz_6027;
  wire       [35:0]   _zz_6028;
  wire       [35:0]   _zz_6029;
  wire       [26:0]   _zz_6030;
  wire       [35:0]   _zz_6031;
  wire       [17:0]   _zz_6032;
  wire       [35:0]   _zz_6033;
  wire       [35:0]   _zz_6034;
  wire       [35:0]   _zz_6035;
  wire       [35:0]   _zz_6036;
  wire       [35:0]   _zz_6037;
  wire       [26:0]   _zz_6038;
  wire       [35:0]   _zz_6039;
  wire       [17:0]   _zz_6040;
  wire       [35:0]   _zz_6041;
  wire       [35:0]   _zz_6042;
  wire       [35:0]   _zz_6043;
  wire       [35:0]   _zz_6044;
  wire       [35:0]   _zz_6045;
  wire       [26:0]   _zz_6046;
  wire       [35:0]   _zz_6047;
  wire       [17:0]   _zz_6048;
  wire       [17:0]   _zz_6049;
  wire       [35:0]   _zz_6050;
  wire       [35:0]   _zz_6051;
  wire       [17:0]   _zz_6052;
  wire       [35:0]   _zz_6053;
  wire       [35:0]   _zz_6054;
  wire       [35:0]   _zz_6055;
  wire       [17:0]   _zz_6056;
  wire       [35:0]   _zz_6057;
  wire       [35:0]   _zz_6058;
  wire       [35:0]   _zz_6059;
  wire       [35:0]   _zz_6060;
  wire       [35:0]   _zz_6061;
  wire       [35:0]   _zz_6062;
  wire       [26:0]   _zz_6063;
  wire       [35:0]   _zz_6064;
  wire       [17:0]   _zz_6065;
  wire       [35:0]   _zz_6066;
  wire       [35:0]   _zz_6067;
  wire       [35:0]   _zz_6068;
  wire       [35:0]   _zz_6069;
  wire       [35:0]   _zz_6070;
  wire       [26:0]   _zz_6071;
  wire       [35:0]   _zz_6072;
  wire       [17:0]   _zz_6073;
  wire       [35:0]   _zz_6074;
  wire       [35:0]   _zz_6075;
  wire       [35:0]   _zz_6076;
  wire       [35:0]   _zz_6077;
  wire       [35:0]   _zz_6078;
  wire       [26:0]   _zz_6079;
  wire       [35:0]   _zz_6080;
  wire       [17:0]   _zz_6081;
  wire       [35:0]   _zz_6082;
  wire       [35:0]   _zz_6083;
  wire       [35:0]   _zz_6084;
  wire       [35:0]   _zz_6085;
  wire       [35:0]   _zz_6086;
  wire       [26:0]   _zz_6087;
  wire       [35:0]   _zz_6088;
  wire       [17:0]   _zz_6089;
  wire       [17:0]   _zz_6090;
  wire       [35:0]   _zz_6091;
  wire       [35:0]   _zz_6092;
  wire       [17:0]   _zz_6093;
  wire       [35:0]   _zz_6094;
  wire       [35:0]   _zz_6095;
  wire       [35:0]   _zz_6096;
  wire       [17:0]   _zz_6097;
  wire       [35:0]   _zz_6098;
  wire       [35:0]   _zz_6099;
  wire       [35:0]   _zz_6100;
  wire       [35:0]   _zz_6101;
  wire       [35:0]   _zz_6102;
  wire       [35:0]   _zz_6103;
  wire       [26:0]   _zz_6104;
  wire       [35:0]   _zz_6105;
  wire       [17:0]   _zz_6106;
  wire       [35:0]   _zz_6107;
  wire       [35:0]   _zz_6108;
  wire       [35:0]   _zz_6109;
  wire       [35:0]   _zz_6110;
  wire       [35:0]   _zz_6111;
  wire       [26:0]   _zz_6112;
  wire       [35:0]   _zz_6113;
  wire       [17:0]   _zz_6114;
  wire       [35:0]   _zz_6115;
  wire       [35:0]   _zz_6116;
  wire       [35:0]   _zz_6117;
  wire       [35:0]   _zz_6118;
  wire       [35:0]   _zz_6119;
  wire       [26:0]   _zz_6120;
  wire       [35:0]   _zz_6121;
  wire       [17:0]   _zz_6122;
  wire       [35:0]   _zz_6123;
  wire       [35:0]   _zz_6124;
  wire       [35:0]   _zz_6125;
  wire       [35:0]   _zz_6126;
  wire       [35:0]   _zz_6127;
  wire       [26:0]   _zz_6128;
  wire       [35:0]   _zz_6129;
  wire       [17:0]   _zz_6130;
  wire       [17:0]   _zz_6131;
  wire       [35:0]   _zz_6132;
  wire       [35:0]   _zz_6133;
  wire       [17:0]   _zz_6134;
  wire       [35:0]   _zz_6135;
  wire       [35:0]   _zz_6136;
  wire       [35:0]   _zz_6137;
  wire       [17:0]   _zz_6138;
  wire       [35:0]   _zz_6139;
  wire       [35:0]   _zz_6140;
  wire       [35:0]   _zz_6141;
  wire       [35:0]   _zz_6142;
  wire       [35:0]   _zz_6143;
  wire       [35:0]   _zz_6144;
  wire       [26:0]   _zz_6145;
  wire       [35:0]   _zz_6146;
  wire       [17:0]   _zz_6147;
  wire       [35:0]   _zz_6148;
  wire       [35:0]   _zz_6149;
  wire       [35:0]   _zz_6150;
  wire       [35:0]   _zz_6151;
  wire       [35:0]   _zz_6152;
  wire       [26:0]   _zz_6153;
  wire       [35:0]   _zz_6154;
  wire       [17:0]   _zz_6155;
  wire       [35:0]   _zz_6156;
  wire       [35:0]   _zz_6157;
  wire       [35:0]   _zz_6158;
  wire       [35:0]   _zz_6159;
  wire       [35:0]   _zz_6160;
  wire       [26:0]   _zz_6161;
  wire       [35:0]   _zz_6162;
  wire       [17:0]   _zz_6163;
  wire       [35:0]   _zz_6164;
  wire       [35:0]   _zz_6165;
  wire       [35:0]   _zz_6166;
  wire       [35:0]   _zz_6167;
  wire       [35:0]   _zz_6168;
  wire       [26:0]   _zz_6169;
  wire       [35:0]   _zz_6170;
  wire       [17:0]   _zz_6171;
  wire       [17:0]   _zz_6172;
  wire       [35:0]   _zz_6173;
  wire       [35:0]   _zz_6174;
  wire       [17:0]   _zz_6175;
  wire       [35:0]   _zz_6176;
  wire       [35:0]   _zz_6177;
  wire       [35:0]   _zz_6178;
  wire       [17:0]   _zz_6179;
  wire       [35:0]   _zz_6180;
  wire       [35:0]   _zz_6181;
  wire       [35:0]   _zz_6182;
  wire       [35:0]   _zz_6183;
  wire       [35:0]   _zz_6184;
  wire       [35:0]   _zz_6185;
  wire       [26:0]   _zz_6186;
  wire       [35:0]   _zz_6187;
  wire       [17:0]   _zz_6188;
  wire       [35:0]   _zz_6189;
  wire       [35:0]   _zz_6190;
  wire       [35:0]   _zz_6191;
  wire       [35:0]   _zz_6192;
  wire       [35:0]   _zz_6193;
  wire       [26:0]   _zz_6194;
  wire       [35:0]   _zz_6195;
  wire       [17:0]   _zz_6196;
  wire       [35:0]   _zz_6197;
  wire       [35:0]   _zz_6198;
  wire       [35:0]   _zz_6199;
  wire       [35:0]   _zz_6200;
  wire       [35:0]   _zz_6201;
  wire       [26:0]   _zz_6202;
  wire       [35:0]   _zz_6203;
  wire       [17:0]   _zz_6204;
  wire       [35:0]   _zz_6205;
  wire       [35:0]   _zz_6206;
  wire       [35:0]   _zz_6207;
  wire       [35:0]   _zz_6208;
  wire       [35:0]   _zz_6209;
  wire       [26:0]   _zz_6210;
  wire       [35:0]   _zz_6211;
  wire       [17:0]   _zz_6212;
  wire       [17:0]   _zz_6213;
  wire       [35:0]   _zz_6214;
  wire       [35:0]   _zz_6215;
  wire       [17:0]   _zz_6216;
  wire       [35:0]   _zz_6217;
  wire       [35:0]   _zz_6218;
  wire       [35:0]   _zz_6219;
  wire       [17:0]   _zz_6220;
  wire       [35:0]   _zz_6221;
  wire       [35:0]   _zz_6222;
  wire       [35:0]   _zz_6223;
  wire       [35:0]   _zz_6224;
  wire       [35:0]   _zz_6225;
  wire       [35:0]   _zz_6226;
  wire       [26:0]   _zz_6227;
  wire       [35:0]   _zz_6228;
  wire       [17:0]   _zz_6229;
  wire       [35:0]   _zz_6230;
  wire       [35:0]   _zz_6231;
  wire       [35:0]   _zz_6232;
  wire       [35:0]   _zz_6233;
  wire       [35:0]   _zz_6234;
  wire       [26:0]   _zz_6235;
  wire       [35:0]   _zz_6236;
  wire       [17:0]   _zz_6237;
  wire       [35:0]   _zz_6238;
  wire       [35:0]   _zz_6239;
  wire       [35:0]   _zz_6240;
  wire       [35:0]   _zz_6241;
  wire       [35:0]   _zz_6242;
  wire       [26:0]   _zz_6243;
  wire       [35:0]   _zz_6244;
  wire       [17:0]   _zz_6245;
  wire       [35:0]   _zz_6246;
  wire       [35:0]   _zz_6247;
  wire       [35:0]   _zz_6248;
  wire       [35:0]   _zz_6249;
  wire       [35:0]   _zz_6250;
  wire       [26:0]   _zz_6251;
  wire       [35:0]   _zz_6252;
  wire       [17:0]   _zz_6253;
  wire       [17:0]   _zz_6254;
  wire       [35:0]   _zz_6255;
  wire       [35:0]   _zz_6256;
  wire       [17:0]   _zz_6257;
  wire       [35:0]   _zz_6258;
  wire       [35:0]   _zz_6259;
  wire       [35:0]   _zz_6260;
  wire       [17:0]   _zz_6261;
  wire       [35:0]   _zz_6262;
  wire       [35:0]   _zz_6263;
  wire       [35:0]   _zz_6264;
  wire       [35:0]   _zz_6265;
  wire       [35:0]   _zz_6266;
  wire       [35:0]   _zz_6267;
  wire       [26:0]   _zz_6268;
  wire       [35:0]   _zz_6269;
  wire       [17:0]   _zz_6270;
  wire       [35:0]   _zz_6271;
  wire       [35:0]   _zz_6272;
  wire       [35:0]   _zz_6273;
  wire       [35:0]   _zz_6274;
  wire       [35:0]   _zz_6275;
  wire       [26:0]   _zz_6276;
  wire       [35:0]   _zz_6277;
  wire       [17:0]   _zz_6278;
  wire       [35:0]   _zz_6279;
  wire       [35:0]   _zz_6280;
  wire       [35:0]   _zz_6281;
  wire       [35:0]   _zz_6282;
  wire       [35:0]   _zz_6283;
  wire       [26:0]   _zz_6284;
  wire       [35:0]   _zz_6285;
  wire       [17:0]   _zz_6286;
  wire       [35:0]   _zz_6287;
  wire       [35:0]   _zz_6288;
  wire       [35:0]   _zz_6289;
  wire       [35:0]   _zz_6290;
  wire       [35:0]   _zz_6291;
  wire       [26:0]   _zz_6292;
  wire       [35:0]   _zz_6293;
  wire       [17:0]   _zz_6294;
  wire       [17:0]   _zz_6295;
  wire       [35:0]   _zz_6296;
  wire       [35:0]   _zz_6297;
  wire       [17:0]   _zz_6298;
  wire       [35:0]   _zz_6299;
  wire       [35:0]   _zz_6300;
  wire       [35:0]   _zz_6301;
  wire       [17:0]   _zz_6302;
  wire       [35:0]   _zz_6303;
  wire       [35:0]   _zz_6304;
  wire       [35:0]   _zz_6305;
  wire       [35:0]   _zz_6306;
  wire       [35:0]   _zz_6307;
  wire       [35:0]   _zz_6308;
  wire       [26:0]   _zz_6309;
  wire       [35:0]   _zz_6310;
  wire       [17:0]   _zz_6311;
  wire       [35:0]   _zz_6312;
  wire       [35:0]   _zz_6313;
  wire       [35:0]   _zz_6314;
  wire       [35:0]   _zz_6315;
  wire       [35:0]   _zz_6316;
  wire       [26:0]   _zz_6317;
  wire       [35:0]   _zz_6318;
  wire       [17:0]   _zz_6319;
  wire       [35:0]   _zz_6320;
  wire       [35:0]   _zz_6321;
  wire       [35:0]   _zz_6322;
  wire       [35:0]   _zz_6323;
  wire       [35:0]   _zz_6324;
  wire       [26:0]   _zz_6325;
  wire       [35:0]   _zz_6326;
  wire       [17:0]   _zz_6327;
  wire       [35:0]   _zz_6328;
  wire       [35:0]   _zz_6329;
  wire       [35:0]   _zz_6330;
  wire       [35:0]   _zz_6331;
  wire       [35:0]   _zz_6332;
  wire       [26:0]   _zz_6333;
  wire       [35:0]   _zz_6334;
  wire       [17:0]   _zz_6335;
  wire       [17:0]   _zz_6336;
  wire       [35:0]   _zz_6337;
  wire       [35:0]   _zz_6338;
  wire       [17:0]   _zz_6339;
  wire       [35:0]   _zz_6340;
  wire       [35:0]   _zz_6341;
  wire       [35:0]   _zz_6342;
  wire       [17:0]   _zz_6343;
  wire       [35:0]   _zz_6344;
  wire       [35:0]   _zz_6345;
  wire       [35:0]   _zz_6346;
  wire       [35:0]   _zz_6347;
  wire       [35:0]   _zz_6348;
  wire       [35:0]   _zz_6349;
  wire       [26:0]   _zz_6350;
  wire       [35:0]   _zz_6351;
  wire       [17:0]   _zz_6352;
  wire       [35:0]   _zz_6353;
  wire       [35:0]   _zz_6354;
  wire       [35:0]   _zz_6355;
  wire       [35:0]   _zz_6356;
  wire       [35:0]   _zz_6357;
  wire       [26:0]   _zz_6358;
  wire       [35:0]   _zz_6359;
  wire       [17:0]   _zz_6360;
  wire       [35:0]   _zz_6361;
  wire       [35:0]   _zz_6362;
  wire       [35:0]   _zz_6363;
  wire       [35:0]   _zz_6364;
  wire       [35:0]   _zz_6365;
  wire       [26:0]   _zz_6366;
  wire       [35:0]   _zz_6367;
  wire       [17:0]   _zz_6368;
  wire       [35:0]   _zz_6369;
  wire       [35:0]   _zz_6370;
  wire       [35:0]   _zz_6371;
  wire       [35:0]   _zz_6372;
  wire       [35:0]   _zz_6373;
  wire       [26:0]   _zz_6374;
  wire       [35:0]   _zz_6375;
  wire       [17:0]   _zz_6376;
  wire       [17:0]   _zz_6377;
  wire       [35:0]   _zz_6378;
  wire       [35:0]   _zz_6379;
  wire       [17:0]   _zz_6380;
  wire       [35:0]   _zz_6381;
  wire       [35:0]   _zz_6382;
  wire       [35:0]   _zz_6383;
  wire       [17:0]   _zz_6384;
  wire       [35:0]   _zz_6385;
  wire       [35:0]   _zz_6386;
  wire       [35:0]   _zz_6387;
  wire       [35:0]   _zz_6388;
  wire       [35:0]   _zz_6389;
  wire       [35:0]   _zz_6390;
  wire       [26:0]   _zz_6391;
  wire       [35:0]   _zz_6392;
  wire       [17:0]   _zz_6393;
  wire       [35:0]   _zz_6394;
  wire       [35:0]   _zz_6395;
  wire       [35:0]   _zz_6396;
  wire       [35:0]   _zz_6397;
  wire       [35:0]   _zz_6398;
  wire       [26:0]   _zz_6399;
  wire       [35:0]   _zz_6400;
  wire       [17:0]   _zz_6401;
  wire       [35:0]   _zz_6402;
  wire       [35:0]   _zz_6403;
  wire       [35:0]   _zz_6404;
  wire       [35:0]   _zz_6405;
  wire       [35:0]   _zz_6406;
  wire       [26:0]   _zz_6407;
  wire       [35:0]   _zz_6408;
  wire       [17:0]   _zz_6409;
  wire       [35:0]   _zz_6410;
  wire       [35:0]   _zz_6411;
  wire       [35:0]   _zz_6412;
  wire       [35:0]   _zz_6413;
  wire       [35:0]   _zz_6414;
  wire       [26:0]   _zz_6415;
  wire       [35:0]   _zz_6416;
  wire       [17:0]   _zz_6417;
  wire       [17:0]   _zz_6418;
  wire       [35:0]   _zz_6419;
  wire       [35:0]   _zz_6420;
  wire       [17:0]   _zz_6421;
  wire       [35:0]   _zz_6422;
  wire       [35:0]   _zz_6423;
  wire       [35:0]   _zz_6424;
  wire       [17:0]   _zz_6425;
  wire       [35:0]   _zz_6426;
  wire       [35:0]   _zz_6427;
  wire       [35:0]   _zz_6428;
  wire       [35:0]   _zz_6429;
  wire       [35:0]   _zz_6430;
  wire       [35:0]   _zz_6431;
  wire       [26:0]   _zz_6432;
  wire       [35:0]   _zz_6433;
  wire       [17:0]   _zz_6434;
  wire       [35:0]   _zz_6435;
  wire       [35:0]   _zz_6436;
  wire       [35:0]   _zz_6437;
  wire       [35:0]   _zz_6438;
  wire       [35:0]   _zz_6439;
  wire       [26:0]   _zz_6440;
  wire       [35:0]   _zz_6441;
  wire       [17:0]   _zz_6442;
  wire       [35:0]   _zz_6443;
  wire       [35:0]   _zz_6444;
  wire       [35:0]   _zz_6445;
  wire       [35:0]   _zz_6446;
  wire       [35:0]   _zz_6447;
  wire       [26:0]   _zz_6448;
  wire       [35:0]   _zz_6449;
  wire       [17:0]   _zz_6450;
  wire       [35:0]   _zz_6451;
  wire       [35:0]   _zz_6452;
  wire       [35:0]   _zz_6453;
  wire       [35:0]   _zz_6454;
  wire       [35:0]   _zz_6455;
  wire       [26:0]   _zz_6456;
  wire       [35:0]   _zz_6457;
  wire       [17:0]   _zz_6458;
  wire       [17:0]   _zz_6459;
  wire       [35:0]   _zz_6460;
  wire       [35:0]   _zz_6461;
  wire       [17:0]   _zz_6462;
  wire       [35:0]   _zz_6463;
  wire       [35:0]   _zz_6464;
  wire       [35:0]   _zz_6465;
  wire       [17:0]   _zz_6466;
  wire       [35:0]   _zz_6467;
  wire       [35:0]   _zz_6468;
  wire       [35:0]   _zz_6469;
  wire       [35:0]   _zz_6470;
  wire       [35:0]   _zz_6471;
  wire       [35:0]   _zz_6472;
  wire       [26:0]   _zz_6473;
  wire       [35:0]   _zz_6474;
  wire       [17:0]   _zz_6475;
  wire       [35:0]   _zz_6476;
  wire       [35:0]   _zz_6477;
  wire       [35:0]   _zz_6478;
  wire       [35:0]   _zz_6479;
  wire       [35:0]   _zz_6480;
  wire       [26:0]   _zz_6481;
  wire       [35:0]   _zz_6482;
  wire       [17:0]   _zz_6483;
  wire       [35:0]   _zz_6484;
  wire       [35:0]   _zz_6485;
  wire       [35:0]   _zz_6486;
  wire       [35:0]   _zz_6487;
  wire       [35:0]   _zz_6488;
  wire       [26:0]   _zz_6489;
  wire       [35:0]   _zz_6490;
  wire       [17:0]   _zz_6491;
  wire       [35:0]   _zz_6492;
  wire       [35:0]   _zz_6493;
  wire       [35:0]   _zz_6494;
  wire       [35:0]   _zz_6495;
  wire       [35:0]   _zz_6496;
  wire       [26:0]   _zz_6497;
  wire       [35:0]   _zz_6498;
  wire       [17:0]   _zz_6499;
  wire       [17:0]   _zz_6500;
  wire       [35:0]   _zz_6501;
  wire       [35:0]   _zz_6502;
  wire       [17:0]   _zz_6503;
  wire       [35:0]   _zz_6504;
  wire       [35:0]   _zz_6505;
  wire       [35:0]   _zz_6506;
  wire       [17:0]   _zz_6507;
  wire       [35:0]   _zz_6508;
  wire       [35:0]   _zz_6509;
  wire       [35:0]   _zz_6510;
  wire       [35:0]   _zz_6511;
  wire       [35:0]   _zz_6512;
  wire       [35:0]   _zz_6513;
  wire       [26:0]   _zz_6514;
  wire       [35:0]   _zz_6515;
  wire       [17:0]   _zz_6516;
  wire       [35:0]   _zz_6517;
  wire       [35:0]   _zz_6518;
  wire       [35:0]   _zz_6519;
  wire       [35:0]   _zz_6520;
  wire       [35:0]   _zz_6521;
  wire       [26:0]   _zz_6522;
  wire       [35:0]   _zz_6523;
  wire       [17:0]   _zz_6524;
  wire       [35:0]   _zz_6525;
  wire       [35:0]   _zz_6526;
  wire       [35:0]   _zz_6527;
  wire       [35:0]   _zz_6528;
  wire       [35:0]   _zz_6529;
  wire       [26:0]   _zz_6530;
  wire       [35:0]   _zz_6531;
  wire       [17:0]   _zz_6532;
  wire       [35:0]   _zz_6533;
  wire       [35:0]   _zz_6534;
  wire       [35:0]   _zz_6535;
  wire       [35:0]   _zz_6536;
  wire       [35:0]   _zz_6537;
  wire       [26:0]   _zz_6538;
  wire       [35:0]   _zz_6539;
  wire       [17:0]   _zz_6540;
  wire       [17:0]   _zz_6541;
  wire       [35:0]   _zz_6542;
  wire       [35:0]   _zz_6543;
  wire       [17:0]   _zz_6544;
  wire       [35:0]   _zz_6545;
  wire       [35:0]   _zz_6546;
  wire       [35:0]   _zz_6547;
  wire       [17:0]   _zz_6548;
  wire       [35:0]   _zz_6549;
  wire       [35:0]   _zz_6550;
  wire       [35:0]   _zz_6551;
  wire       [35:0]   _zz_6552;
  wire       [35:0]   _zz_6553;
  wire       [35:0]   _zz_6554;
  wire       [26:0]   _zz_6555;
  wire       [35:0]   _zz_6556;
  wire       [17:0]   _zz_6557;
  wire       [35:0]   _zz_6558;
  wire       [35:0]   _zz_6559;
  wire       [35:0]   _zz_6560;
  wire       [35:0]   _zz_6561;
  wire       [35:0]   _zz_6562;
  wire       [26:0]   _zz_6563;
  wire       [35:0]   _zz_6564;
  wire       [17:0]   _zz_6565;
  wire       [35:0]   _zz_6566;
  wire       [35:0]   _zz_6567;
  wire       [35:0]   _zz_6568;
  wire       [35:0]   _zz_6569;
  wire       [35:0]   _zz_6570;
  wire       [26:0]   _zz_6571;
  wire       [35:0]   _zz_6572;
  wire       [17:0]   _zz_6573;
  wire       [35:0]   _zz_6574;
  wire       [35:0]   _zz_6575;
  wire       [35:0]   _zz_6576;
  wire       [35:0]   _zz_6577;
  wire       [35:0]   _zz_6578;
  wire       [26:0]   _zz_6579;
  wire       [35:0]   _zz_6580;
  wire       [17:0]   _zz_6581;
  wire       [17:0]   _zz_6582;
  wire       [35:0]   _zz_6583;
  wire       [35:0]   _zz_6584;
  wire       [17:0]   _zz_6585;
  wire       [35:0]   _zz_6586;
  wire       [35:0]   _zz_6587;
  wire       [35:0]   _zz_6588;
  wire       [17:0]   _zz_6589;
  wire       [35:0]   _zz_6590;
  wire       [35:0]   _zz_6591;
  wire       [35:0]   _zz_6592;
  wire       [35:0]   _zz_6593;
  wire       [35:0]   _zz_6594;
  wire       [35:0]   _zz_6595;
  wire       [26:0]   _zz_6596;
  wire       [35:0]   _zz_6597;
  wire       [17:0]   _zz_6598;
  wire       [35:0]   _zz_6599;
  wire       [35:0]   _zz_6600;
  wire       [35:0]   _zz_6601;
  wire       [35:0]   _zz_6602;
  wire       [35:0]   _zz_6603;
  wire       [26:0]   _zz_6604;
  wire       [35:0]   _zz_6605;
  wire       [17:0]   _zz_6606;
  wire       [35:0]   _zz_6607;
  wire       [35:0]   _zz_6608;
  wire       [35:0]   _zz_6609;
  wire       [35:0]   _zz_6610;
  wire       [35:0]   _zz_6611;
  wire       [26:0]   _zz_6612;
  wire       [35:0]   _zz_6613;
  wire       [17:0]   _zz_6614;
  wire       [35:0]   _zz_6615;
  wire       [35:0]   _zz_6616;
  wire       [35:0]   _zz_6617;
  wire       [35:0]   _zz_6618;
  wire       [35:0]   _zz_6619;
  wire       [26:0]   _zz_6620;
  wire       [35:0]   _zz_6621;
  wire       [17:0]   _zz_6622;
  wire       [17:0]   _zz_6623;
  wire       [35:0]   _zz_6624;
  wire       [35:0]   _zz_6625;
  wire       [17:0]   _zz_6626;
  wire       [35:0]   _zz_6627;
  wire       [35:0]   _zz_6628;
  wire       [35:0]   _zz_6629;
  wire       [17:0]   _zz_6630;
  wire       [35:0]   _zz_6631;
  wire       [35:0]   _zz_6632;
  wire       [35:0]   _zz_6633;
  wire       [35:0]   _zz_6634;
  wire       [35:0]   _zz_6635;
  wire       [35:0]   _zz_6636;
  wire       [26:0]   _zz_6637;
  wire       [35:0]   _zz_6638;
  wire       [17:0]   _zz_6639;
  wire       [35:0]   _zz_6640;
  wire       [35:0]   _zz_6641;
  wire       [35:0]   _zz_6642;
  wire       [35:0]   _zz_6643;
  wire       [35:0]   _zz_6644;
  wire       [26:0]   _zz_6645;
  wire       [35:0]   _zz_6646;
  wire       [17:0]   _zz_6647;
  wire       [35:0]   _zz_6648;
  wire       [35:0]   _zz_6649;
  wire       [35:0]   _zz_6650;
  wire       [35:0]   _zz_6651;
  wire       [35:0]   _zz_6652;
  wire       [26:0]   _zz_6653;
  wire       [35:0]   _zz_6654;
  wire       [17:0]   _zz_6655;
  wire       [35:0]   _zz_6656;
  wire       [35:0]   _zz_6657;
  wire       [35:0]   _zz_6658;
  wire       [35:0]   _zz_6659;
  wire       [35:0]   _zz_6660;
  wire       [26:0]   _zz_6661;
  wire       [35:0]   _zz_6662;
  wire       [17:0]   _zz_6663;
  wire       [17:0]   _zz_6664;
  wire       [35:0]   _zz_6665;
  wire       [35:0]   _zz_6666;
  wire       [17:0]   _zz_6667;
  wire       [35:0]   _zz_6668;
  wire       [35:0]   _zz_6669;
  wire       [35:0]   _zz_6670;
  wire       [17:0]   _zz_6671;
  wire       [35:0]   _zz_6672;
  wire       [35:0]   _zz_6673;
  wire       [35:0]   _zz_6674;
  wire       [35:0]   _zz_6675;
  wire       [35:0]   _zz_6676;
  wire       [35:0]   _zz_6677;
  wire       [26:0]   _zz_6678;
  wire       [35:0]   _zz_6679;
  wire       [17:0]   _zz_6680;
  wire       [35:0]   _zz_6681;
  wire       [35:0]   _zz_6682;
  wire       [35:0]   _zz_6683;
  wire       [35:0]   _zz_6684;
  wire       [35:0]   _zz_6685;
  wire       [26:0]   _zz_6686;
  wire       [35:0]   _zz_6687;
  wire       [17:0]   _zz_6688;
  wire       [35:0]   _zz_6689;
  wire       [35:0]   _zz_6690;
  wire       [35:0]   _zz_6691;
  wire       [35:0]   _zz_6692;
  wire       [35:0]   _zz_6693;
  wire       [26:0]   _zz_6694;
  wire       [35:0]   _zz_6695;
  wire       [17:0]   _zz_6696;
  wire       [35:0]   _zz_6697;
  wire       [35:0]   _zz_6698;
  wire       [35:0]   _zz_6699;
  wire       [35:0]   _zz_6700;
  wire       [35:0]   _zz_6701;
  wire       [26:0]   _zz_6702;
  wire       [35:0]   _zz_6703;
  wire       [17:0]   _zz_6704;
  wire       [17:0]   _zz_6705;
  wire       [35:0]   _zz_6706;
  wire       [35:0]   _zz_6707;
  wire       [17:0]   _zz_6708;
  wire       [35:0]   _zz_6709;
  wire       [35:0]   _zz_6710;
  wire       [35:0]   _zz_6711;
  wire       [17:0]   _zz_6712;
  wire       [35:0]   _zz_6713;
  wire       [35:0]   _zz_6714;
  wire       [35:0]   _zz_6715;
  wire       [35:0]   _zz_6716;
  wire       [35:0]   _zz_6717;
  wire       [35:0]   _zz_6718;
  wire       [26:0]   _zz_6719;
  wire       [35:0]   _zz_6720;
  wire       [17:0]   _zz_6721;
  wire       [35:0]   _zz_6722;
  wire       [35:0]   _zz_6723;
  wire       [35:0]   _zz_6724;
  wire       [35:0]   _zz_6725;
  wire       [35:0]   _zz_6726;
  wire       [26:0]   _zz_6727;
  wire       [35:0]   _zz_6728;
  wire       [17:0]   _zz_6729;
  wire       [35:0]   _zz_6730;
  wire       [35:0]   _zz_6731;
  wire       [35:0]   _zz_6732;
  wire       [35:0]   _zz_6733;
  wire       [35:0]   _zz_6734;
  wire       [26:0]   _zz_6735;
  wire       [35:0]   _zz_6736;
  wire       [17:0]   _zz_6737;
  wire       [35:0]   _zz_6738;
  wire       [35:0]   _zz_6739;
  wire       [35:0]   _zz_6740;
  wire       [35:0]   _zz_6741;
  wire       [35:0]   _zz_6742;
  wire       [26:0]   _zz_6743;
  wire       [35:0]   _zz_6744;
  wire       [17:0]   _zz_6745;
  wire       [17:0]   _zz_6746;
  wire       [35:0]   _zz_6747;
  wire       [35:0]   _zz_6748;
  wire       [17:0]   _zz_6749;
  wire       [35:0]   _zz_6750;
  wire       [35:0]   _zz_6751;
  wire       [35:0]   _zz_6752;
  wire       [17:0]   _zz_6753;
  wire       [35:0]   _zz_6754;
  wire       [35:0]   _zz_6755;
  wire       [35:0]   _zz_6756;
  wire       [35:0]   _zz_6757;
  wire       [35:0]   _zz_6758;
  wire       [35:0]   _zz_6759;
  wire       [26:0]   _zz_6760;
  wire       [35:0]   _zz_6761;
  wire       [17:0]   _zz_6762;
  wire       [35:0]   _zz_6763;
  wire       [35:0]   _zz_6764;
  wire       [35:0]   _zz_6765;
  wire       [35:0]   _zz_6766;
  wire       [35:0]   _zz_6767;
  wire       [26:0]   _zz_6768;
  wire       [35:0]   _zz_6769;
  wire       [17:0]   _zz_6770;
  wire       [35:0]   _zz_6771;
  wire       [35:0]   _zz_6772;
  wire       [35:0]   _zz_6773;
  wire       [35:0]   _zz_6774;
  wire       [35:0]   _zz_6775;
  wire       [26:0]   _zz_6776;
  wire       [35:0]   _zz_6777;
  wire       [17:0]   _zz_6778;
  wire       [35:0]   _zz_6779;
  wire       [35:0]   _zz_6780;
  wire       [35:0]   _zz_6781;
  wire       [35:0]   _zz_6782;
  wire       [35:0]   _zz_6783;
  wire       [26:0]   _zz_6784;
  wire       [35:0]   _zz_6785;
  wire       [17:0]   _zz_6786;
  wire       [17:0]   _zz_6787;
  wire       [35:0]   _zz_6788;
  wire       [35:0]   _zz_6789;
  wire       [17:0]   _zz_6790;
  wire       [35:0]   _zz_6791;
  wire       [35:0]   _zz_6792;
  wire       [35:0]   _zz_6793;
  wire       [17:0]   _zz_6794;
  wire       [35:0]   _zz_6795;
  wire       [35:0]   _zz_6796;
  wire       [35:0]   _zz_6797;
  wire       [35:0]   _zz_6798;
  wire       [35:0]   _zz_6799;
  wire       [35:0]   _zz_6800;
  wire       [26:0]   _zz_6801;
  wire       [35:0]   _zz_6802;
  wire       [17:0]   _zz_6803;
  wire       [35:0]   _zz_6804;
  wire       [35:0]   _zz_6805;
  wire       [35:0]   _zz_6806;
  wire       [35:0]   _zz_6807;
  wire       [35:0]   _zz_6808;
  wire       [26:0]   _zz_6809;
  wire       [35:0]   _zz_6810;
  wire       [17:0]   _zz_6811;
  wire       [35:0]   _zz_6812;
  wire       [35:0]   _zz_6813;
  wire       [35:0]   _zz_6814;
  wire       [35:0]   _zz_6815;
  wire       [35:0]   _zz_6816;
  wire       [26:0]   _zz_6817;
  wire       [35:0]   _zz_6818;
  wire       [17:0]   _zz_6819;
  wire       [35:0]   _zz_6820;
  wire       [35:0]   _zz_6821;
  wire       [35:0]   _zz_6822;
  wire       [35:0]   _zz_6823;
  wire       [35:0]   _zz_6824;
  wire       [26:0]   _zz_6825;
  wire       [35:0]   _zz_6826;
  wire       [17:0]   _zz_6827;
  wire       [17:0]   _zz_6828;
  wire       [35:0]   _zz_6829;
  wire       [35:0]   _zz_6830;
  wire       [17:0]   _zz_6831;
  wire       [35:0]   _zz_6832;
  wire       [35:0]   _zz_6833;
  wire       [35:0]   _zz_6834;
  wire       [17:0]   _zz_6835;
  wire       [35:0]   _zz_6836;
  wire       [35:0]   _zz_6837;
  wire       [35:0]   _zz_6838;
  wire       [35:0]   _zz_6839;
  wire       [35:0]   _zz_6840;
  wire       [35:0]   _zz_6841;
  wire       [26:0]   _zz_6842;
  wire       [35:0]   _zz_6843;
  wire       [17:0]   _zz_6844;
  wire       [35:0]   _zz_6845;
  wire       [35:0]   _zz_6846;
  wire       [35:0]   _zz_6847;
  wire       [35:0]   _zz_6848;
  wire       [35:0]   _zz_6849;
  wire       [26:0]   _zz_6850;
  wire       [35:0]   _zz_6851;
  wire       [17:0]   _zz_6852;
  wire       [35:0]   _zz_6853;
  wire       [35:0]   _zz_6854;
  wire       [35:0]   _zz_6855;
  wire       [35:0]   _zz_6856;
  wire       [35:0]   _zz_6857;
  wire       [26:0]   _zz_6858;
  wire       [35:0]   _zz_6859;
  wire       [17:0]   _zz_6860;
  wire       [35:0]   _zz_6861;
  wire       [35:0]   _zz_6862;
  wire       [35:0]   _zz_6863;
  wire       [35:0]   _zz_6864;
  wire       [35:0]   _zz_6865;
  wire       [26:0]   _zz_6866;
  wire       [35:0]   _zz_6867;
  wire       [17:0]   _zz_6868;
  wire       [17:0]   _zz_6869;
  wire       [35:0]   _zz_6870;
  wire       [35:0]   _zz_6871;
  wire       [17:0]   _zz_6872;
  wire       [35:0]   _zz_6873;
  wire       [35:0]   _zz_6874;
  wire       [35:0]   _zz_6875;
  wire       [17:0]   _zz_6876;
  wire       [35:0]   _zz_6877;
  wire       [35:0]   _zz_6878;
  wire       [35:0]   _zz_6879;
  wire       [35:0]   _zz_6880;
  wire       [35:0]   _zz_6881;
  wire       [35:0]   _zz_6882;
  wire       [26:0]   _zz_6883;
  wire       [35:0]   _zz_6884;
  wire       [17:0]   _zz_6885;
  wire       [35:0]   _zz_6886;
  wire       [35:0]   _zz_6887;
  wire       [35:0]   _zz_6888;
  wire       [35:0]   _zz_6889;
  wire       [35:0]   _zz_6890;
  wire       [26:0]   _zz_6891;
  wire       [35:0]   _zz_6892;
  wire       [17:0]   _zz_6893;
  wire       [35:0]   _zz_6894;
  wire       [35:0]   _zz_6895;
  wire       [35:0]   _zz_6896;
  wire       [35:0]   _zz_6897;
  wire       [35:0]   _zz_6898;
  wire       [26:0]   _zz_6899;
  wire       [35:0]   _zz_6900;
  wire       [17:0]   _zz_6901;
  wire       [35:0]   _zz_6902;
  wire       [35:0]   _zz_6903;
  wire       [35:0]   _zz_6904;
  wire       [35:0]   _zz_6905;
  wire       [35:0]   _zz_6906;
  wire       [26:0]   _zz_6907;
  wire       [35:0]   _zz_6908;
  wire       [17:0]   _zz_6909;
  wire       [17:0]   _zz_6910;
  wire       [35:0]   _zz_6911;
  wire       [35:0]   _zz_6912;
  wire       [17:0]   _zz_6913;
  wire       [35:0]   _zz_6914;
  wire       [35:0]   _zz_6915;
  wire       [35:0]   _zz_6916;
  wire       [17:0]   _zz_6917;
  wire       [35:0]   _zz_6918;
  wire       [35:0]   _zz_6919;
  wire       [35:0]   _zz_6920;
  wire       [35:0]   _zz_6921;
  wire       [35:0]   _zz_6922;
  wire       [35:0]   _zz_6923;
  wire       [26:0]   _zz_6924;
  wire       [35:0]   _zz_6925;
  wire       [17:0]   _zz_6926;
  wire       [35:0]   _zz_6927;
  wire       [35:0]   _zz_6928;
  wire       [35:0]   _zz_6929;
  wire       [35:0]   _zz_6930;
  wire       [35:0]   _zz_6931;
  wire       [26:0]   _zz_6932;
  wire       [35:0]   _zz_6933;
  wire       [17:0]   _zz_6934;
  wire       [35:0]   _zz_6935;
  wire       [35:0]   _zz_6936;
  wire       [35:0]   _zz_6937;
  wire       [35:0]   _zz_6938;
  wire       [35:0]   _zz_6939;
  wire       [26:0]   _zz_6940;
  wire       [35:0]   _zz_6941;
  wire       [17:0]   _zz_6942;
  wire       [35:0]   _zz_6943;
  wire       [35:0]   _zz_6944;
  wire       [35:0]   _zz_6945;
  wire       [35:0]   _zz_6946;
  wire       [35:0]   _zz_6947;
  wire       [26:0]   _zz_6948;
  wire       [35:0]   _zz_6949;
  wire       [17:0]   _zz_6950;
  wire       [17:0]   _zz_6951;
  wire       [35:0]   _zz_6952;
  wire       [35:0]   _zz_6953;
  wire       [17:0]   _zz_6954;
  wire       [35:0]   _zz_6955;
  wire       [35:0]   _zz_6956;
  wire       [35:0]   _zz_6957;
  wire       [17:0]   _zz_6958;
  wire       [35:0]   _zz_6959;
  wire       [35:0]   _zz_6960;
  wire       [35:0]   _zz_6961;
  wire       [35:0]   _zz_6962;
  wire       [35:0]   _zz_6963;
  wire       [35:0]   _zz_6964;
  wire       [26:0]   _zz_6965;
  wire       [35:0]   _zz_6966;
  wire       [17:0]   _zz_6967;
  wire       [35:0]   _zz_6968;
  wire       [35:0]   _zz_6969;
  wire       [35:0]   _zz_6970;
  wire       [35:0]   _zz_6971;
  wire       [35:0]   _zz_6972;
  wire       [26:0]   _zz_6973;
  wire       [35:0]   _zz_6974;
  wire       [17:0]   _zz_6975;
  wire       [35:0]   _zz_6976;
  wire       [35:0]   _zz_6977;
  wire       [35:0]   _zz_6978;
  wire       [35:0]   _zz_6979;
  wire       [35:0]   _zz_6980;
  wire       [26:0]   _zz_6981;
  wire       [35:0]   _zz_6982;
  wire       [17:0]   _zz_6983;
  wire       [35:0]   _zz_6984;
  wire       [35:0]   _zz_6985;
  wire       [35:0]   _zz_6986;
  wire       [35:0]   _zz_6987;
  wire       [35:0]   _zz_6988;
  wire       [26:0]   _zz_6989;
  wire       [35:0]   _zz_6990;
  wire       [17:0]   _zz_6991;
  wire       [17:0]   _zz_6992;
  wire       [35:0]   _zz_6993;
  wire       [35:0]   _zz_6994;
  wire       [17:0]   _zz_6995;
  wire       [35:0]   _zz_6996;
  wire       [35:0]   _zz_6997;
  wire       [35:0]   _zz_6998;
  wire       [17:0]   _zz_6999;
  wire       [35:0]   _zz_7000;
  wire       [35:0]   _zz_7001;
  wire       [35:0]   _zz_7002;
  wire       [35:0]   _zz_7003;
  wire       [35:0]   _zz_7004;
  wire       [35:0]   _zz_7005;
  wire       [26:0]   _zz_7006;
  wire       [35:0]   _zz_7007;
  wire       [17:0]   _zz_7008;
  wire       [35:0]   _zz_7009;
  wire       [35:0]   _zz_7010;
  wire       [35:0]   _zz_7011;
  wire       [35:0]   _zz_7012;
  wire       [35:0]   _zz_7013;
  wire       [26:0]   _zz_7014;
  wire       [35:0]   _zz_7015;
  wire       [17:0]   _zz_7016;
  wire       [35:0]   _zz_7017;
  wire       [35:0]   _zz_7018;
  wire       [35:0]   _zz_7019;
  wire       [35:0]   _zz_7020;
  wire       [35:0]   _zz_7021;
  wire       [26:0]   _zz_7022;
  wire       [35:0]   _zz_7023;
  wire       [17:0]   _zz_7024;
  wire       [35:0]   _zz_7025;
  wire       [35:0]   _zz_7026;
  wire       [35:0]   _zz_7027;
  wire       [35:0]   _zz_7028;
  wire       [35:0]   _zz_7029;
  wire       [26:0]   _zz_7030;
  wire       [35:0]   _zz_7031;
  wire       [17:0]   _zz_7032;
  wire       [17:0]   _zz_7033;
  wire       [35:0]   _zz_7034;
  wire       [35:0]   _zz_7035;
  wire       [17:0]   _zz_7036;
  wire       [35:0]   _zz_7037;
  wire       [35:0]   _zz_7038;
  wire       [35:0]   _zz_7039;
  wire       [17:0]   _zz_7040;
  wire       [35:0]   _zz_7041;
  wire       [35:0]   _zz_7042;
  wire       [35:0]   _zz_7043;
  wire       [35:0]   _zz_7044;
  wire       [35:0]   _zz_7045;
  wire       [35:0]   _zz_7046;
  wire       [26:0]   _zz_7047;
  wire       [35:0]   _zz_7048;
  wire       [17:0]   _zz_7049;
  wire       [35:0]   _zz_7050;
  wire       [35:0]   _zz_7051;
  wire       [35:0]   _zz_7052;
  wire       [35:0]   _zz_7053;
  wire       [35:0]   _zz_7054;
  wire       [26:0]   _zz_7055;
  wire       [35:0]   _zz_7056;
  wire       [17:0]   _zz_7057;
  wire       [35:0]   _zz_7058;
  wire       [35:0]   _zz_7059;
  wire       [35:0]   _zz_7060;
  wire       [35:0]   _zz_7061;
  wire       [35:0]   _zz_7062;
  wire       [26:0]   _zz_7063;
  wire       [35:0]   _zz_7064;
  wire       [17:0]   _zz_7065;
  wire       [35:0]   _zz_7066;
  wire       [35:0]   _zz_7067;
  wire       [35:0]   _zz_7068;
  wire       [35:0]   _zz_7069;
  wire       [35:0]   _zz_7070;
  wire       [26:0]   _zz_7071;
  wire       [35:0]   _zz_7072;
  wire       [17:0]   _zz_7073;
  wire       [17:0]   _zz_7074;
  wire       [35:0]   _zz_7075;
  wire       [35:0]   _zz_7076;
  wire       [17:0]   _zz_7077;
  wire       [35:0]   _zz_7078;
  wire       [35:0]   _zz_7079;
  wire       [35:0]   _zz_7080;
  wire       [17:0]   _zz_7081;
  wire       [35:0]   _zz_7082;
  wire       [35:0]   _zz_7083;
  wire       [35:0]   _zz_7084;
  wire       [35:0]   _zz_7085;
  wire       [35:0]   _zz_7086;
  wire       [35:0]   _zz_7087;
  wire       [26:0]   _zz_7088;
  wire       [35:0]   _zz_7089;
  wire       [17:0]   _zz_7090;
  wire       [35:0]   _zz_7091;
  wire       [35:0]   _zz_7092;
  wire       [35:0]   _zz_7093;
  wire       [35:0]   _zz_7094;
  wire       [35:0]   _zz_7095;
  wire       [26:0]   _zz_7096;
  wire       [35:0]   _zz_7097;
  wire       [17:0]   _zz_7098;
  wire       [35:0]   _zz_7099;
  wire       [35:0]   _zz_7100;
  wire       [35:0]   _zz_7101;
  wire       [35:0]   _zz_7102;
  wire       [35:0]   _zz_7103;
  wire       [26:0]   _zz_7104;
  wire       [35:0]   _zz_7105;
  wire       [17:0]   _zz_7106;
  wire       [35:0]   _zz_7107;
  wire       [35:0]   _zz_7108;
  wire       [35:0]   _zz_7109;
  wire       [35:0]   _zz_7110;
  wire       [35:0]   _zz_7111;
  wire       [26:0]   _zz_7112;
  wire       [35:0]   _zz_7113;
  wire       [17:0]   _zz_7114;
  wire       [17:0]   _zz_7115;
  wire       [35:0]   _zz_7116;
  wire       [35:0]   _zz_7117;
  wire       [17:0]   _zz_7118;
  wire       [35:0]   _zz_7119;
  wire       [35:0]   _zz_7120;
  wire       [35:0]   _zz_7121;
  wire       [17:0]   _zz_7122;
  wire       [35:0]   _zz_7123;
  wire       [35:0]   _zz_7124;
  wire       [35:0]   _zz_7125;
  wire       [35:0]   _zz_7126;
  wire       [35:0]   _zz_7127;
  wire       [35:0]   _zz_7128;
  wire       [26:0]   _zz_7129;
  wire       [35:0]   _zz_7130;
  wire       [17:0]   _zz_7131;
  wire       [35:0]   _zz_7132;
  wire       [35:0]   _zz_7133;
  wire       [35:0]   _zz_7134;
  wire       [35:0]   _zz_7135;
  wire       [35:0]   _zz_7136;
  wire       [26:0]   _zz_7137;
  wire       [35:0]   _zz_7138;
  wire       [17:0]   _zz_7139;
  wire       [35:0]   _zz_7140;
  wire       [35:0]   _zz_7141;
  wire       [35:0]   _zz_7142;
  wire       [35:0]   _zz_7143;
  wire       [35:0]   _zz_7144;
  wire       [26:0]   _zz_7145;
  wire       [35:0]   _zz_7146;
  wire       [17:0]   _zz_7147;
  wire       [35:0]   _zz_7148;
  wire       [35:0]   _zz_7149;
  wire       [35:0]   _zz_7150;
  wire       [35:0]   _zz_7151;
  wire       [35:0]   _zz_7152;
  wire       [26:0]   _zz_7153;
  wire       [35:0]   _zz_7154;
  wire       [17:0]   _zz_7155;
  wire       [17:0]   _zz_7156;
  wire       [35:0]   _zz_7157;
  wire       [35:0]   _zz_7158;
  wire       [17:0]   _zz_7159;
  wire       [35:0]   _zz_7160;
  wire       [35:0]   _zz_7161;
  wire       [35:0]   _zz_7162;
  wire       [17:0]   _zz_7163;
  wire       [35:0]   _zz_7164;
  wire       [35:0]   _zz_7165;
  wire       [35:0]   _zz_7166;
  wire       [35:0]   _zz_7167;
  wire       [35:0]   _zz_7168;
  wire       [35:0]   _zz_7169;
  wire       [26:0]   _zz_7170;
  wire       [35:0]   _zz_7171;
  wire       [17:0]   _zz_7172;
  wire       [35:0]   _zz_7173;
  wire       [35:0]   _zz_7174;
  wire       [35:0]   _zz_7175;
  wire       [35:0]   _zz_7176;
  wire       [35:0]   _zz_7177;
  wire       [26:0]   _zz_7178;
  wire       [35:0]   _zz_7179;
  wire       [17:0]   _zz_7180;
  wire       [35:0]   _zz_7181;
  wire       [35:0]   _zz_7182;
  wire       [35:0]   _zz_7183;
  wire       [35:0]   _zz_7184;
  wire       [35:0]   _zz_7185;
  wire       [26:0]   _zz_7186;
  wire       [35:0]   _zz_7187;
  wire       [17:0]   _zz_7188;
  wire       [35:0]   _zz_7189;
  wire       [35:0]   _zz_7190;
  wire       [35:0]   _zz_7191;
  wire       [35:0]   _zz_7192;
  wire       [35:0]   _zz_7193;
  wire       [26:0]   _zz_7194;
  wire       [35:0]   _zz_7195;
  wire       [17:0]   _zz_7196;
  wire       [17:0]   _zz_7197;
  wire       [35:0]   _zz_7198;
  wire       [35:0]   _zz_7199;
  wire       [17:0]   _zz_7200;
  wire       [35:0]   _zz_7201;
  wire       [35:0]   _zz_7202;
  wire       [35:0]   _zz_7203;
  wire       [17:0]   _zz_7204;
  wire       [35:0]   _zz_7205;
  wire       [35:0]   _zz_7206;
  wire       [35:0]   _zz_7207;
  wire       [35:0]   _zz_7208;
  wire       [35:0]   _zz_7209;
  wire       [35:0]   _zz_7210;
  wire       [26:0]   _zz_7211;
  wire       [35:0]   _zz_7212;
  wire       [17:0]   _zz_7213;
  wire       [35:0]   _zz_7214;
  wire       [35:0]   _zz_7215;
  wire       [35:0]   _zz_7216;
  wire       [35:0]   _zz_7217;
  wire       [35:0]   _zz_7218;
  wire       [26:0]   _zz_7219;
  wire       [35:0]   _zz_7220;
  wire       [17:0]   _zz_7221;
  wire       [35:0]   _zz_7222;
  wire       [35:0]   _zz_7223;
  wire       [35:0]   _zz_7224;
  wire       [35:0]   _zz_7225;
  wire       [35:0]   _zz_7226;
  wire       [26:0]   _zz_7227;
  wire       [35:0]   _zz_7228;
  wire       [17:0]   _zz_7229;
  wire       [35:0]   _zz_7230;
  wire       [35:0]   _zz_7231;
  wire       [35:0]   _zz_7232;
  wire       [35:0]   _zz_7233;
  wire       [35:0]   _zz_7234;
  wire       [26:0]   _zz_7235;
  wire       [35:0]   _zz_7236;
  wire       [17:0]   _zz_7237;
  wire       [17:0]   _zz_7238;
  wire       [35:0]   _zz_7239;
  wire       [35:0]   _zz_7240;
  wire       [17:0]   _zz_7241;
  wire       [35:0]   _zz_7242;
  wire       [35:0]   _zz_7243;
  wire       [35:0]   _zz_7244;
  wire       [17:0]   _zz_7245;
  wire       [35:0]   _zz_7246;
  wire       [35:0]   _zz_7247;
  wire       [35:0]   _zz_7248;
  wire       [35:0]   _zz_7249;
  wire       [35:0]   _zz_7250;
  wire       [35:0]   _zz_7251;
  wire       [26:0]   _zz_7252;
  wire       [35:0]   _zz_7253;
  wire       [17:0]   _zz_7254;
  wire       [35:0]   _zz_7255;
  wire       [35:0]   _zz_7256;
  wire       [35:0]   _zz_7257;
  wire       [35:0]   _zz_7258;
  wire       [35:0]   _zz_7259;
  wire       [26:0]   _zz_7260;
  wire       [35:0]   _zz_7261;
  wire       [17:0]   _zz_7262;
  wire       [35:0]   _zz_7263;
  wire       [35:0]   _zz_7264;
  wire       [35:0]   _zz_7265;
  wire       [35:0]   _zz_7266;
  wire       [35:0]   _zz_7267;
  wire       [26:0]   _zz_7268;
  wire       [35:0]   _zz_7269;
  wire       [17:0]   _zz_7270;
  wire       [35:0]   _zz_7271;
  wire       [35:0]   _zz_7272;
  wire       [35:0]   _zz_7273;
  wire       [35:0]   _zz_7274;
  wire       [35:0]   _zz_7275;
  wire       [26:0]   _zz_7276;
  wire       [35:0]   _zz_7277;
  wire       [17:0]   _zz_7278;
  wire       [17:0]   _zz_7279;
  wire       [35:0]   _zz_7280;
  wire       [35:0]   _zz_7281;
  wire       [17:0]   _zz_7282;
  wire       [35:0]   _zz_7283;
  wire       [35:0]   _zz_7284;
  wire       [35:0]   _zz_7285;
  wire       [17:0]   _zz_7286;
  wire       [35:0]   _zz_7287;
  wire       [35:0]   _zz_7288;
  wire       [35:0]   _zz_7289;
  wire       [35:0]   _zz_7290;
  wire       [35:0]   _zz_7291;
  wire       [35:0]   _zz_7292;
  wire       [26:0]   _zz_7293;
  wire       [35:0]   _zz_7294;
  wire       [17:0]   _zz_7295;
  wire       [35:0]   _zz_7296;
  wire       [35:0]   _zz_7297;
  wire       [35:0]   _zz_7298;
  wire       [35:0]   _zz_7299;
  wire       [35:0]   _zz_7300;
  wire       [26:0]   _zz_7301;
  wire       [35:0]   _zz_7302;
  wire       [17:0]   _zz_7303;
  wire       [35:0]   _zz_7304;
  wire       [35:0]   _zz_7305;
  wire       [35:0]   _zz_7306;
  wire       [35:0]   _zz_7307;
  wire       [35:0]   _zz_7308;
  wire       [26:0]   _zz_7309;
  wire       [35:0]   _zz_7310;
  wire       [17:0]   _zz_7311;
  wire       [35:0]   _zz_7312;
  wire       [35:0]   _zz_7313;
  wire       [35:0]   _zz_7314;
  wire       [35:0]   _zz_7315;
  wire       [35:0]   _zz_7316;
  wire       [26:0]   _zz_7317;
  wire       [35:0]   _zz_7318;
  wire       [17:0]   _zz_7319;
  wire       [17:0]   _zz_7320;
  wire       [35:0]   _zz_7321;
  wire       [35:0]   _zz_7322;
  wire       [17:0]   _zz_7323;
  wire       [35:0]   _zz_7324;
  wire       [35:0]   _zz_7325;
  wire       [35:0]   _zz_7326;
  wire       [17:0]   _zz_7327;
  wire       [35:0]   _zz_7328;
  wire       [35:0]   _zz_7329;
  wire       [35:0]   _zz_7330;
  wire       [35:0]   _zz_7331;
  wire       [35:0]   _zz_7332;
  wire       [35:0]   _zz_7333;
  wire       [26:0]   _zz_7334;
  wire       [35:0]   _zz_7335;
  wire       [17:0]   _zz_7336;
  wire       [35:0]   _zz_7337;
  wire       [35:0]   _zz_7338;
  wire       [35:0]   _zz_7339;
  wire       [35:0]   _zz_7340;
  wire       [35:0]   _zz_7341;
  wire       [26:0]   _zz_7342;
  wire       [35:0]   _zz_7343;
  wire       [17:0]   _zz_7344;
  wire       [35:0]   _zz_7345;
  wire       [35:0]   _zz_7346;
  wire       [35:0]   _zz_7347;
  wire       [35:0]   _zz_7348;
  wire       [35:0]   _zz_7349;
  wire       [26:0]   _zz_7350;
  wire       [35:0]   _zz_7351;
  wire       [17:0]   _zz_7352;
  wire       [35:0]   _zz_7353;
  wire       [35:0]   _zz_7354;
  wire       [35:0]   _zz_7355;
  wire       [35:0]   _zz_7356;
  wire       [35:0]   _zz_7357;
  wire       [26:0]   _zz_7358;
  wire       [35:0]   _zz_7359;
  wire       [17:0]   _zz_7360;
  wire       [17:0]   _zz_7361;
  wire       [35:0]   _zz_7362;
  wire       [35:0]   _zz_7363;
  wire       [17:0]   _zz_7364;
  wire       [35:0]   _zz_7365;
  wire       [35:0]   _zz_7366;
  wire       [35:0]   _zz_7367;
  wire       [17:0]   _zz_7368;
  wire       [35:0]   _zz_7369;
  wire       [35:0]   _zz_7370;
  wire       [35:0]   _zz_7371;
  wire       [35:0]   _zz_7372;
  wire       [35:0]   _zz_7373;
  wire       [35:0]   _zz_7374;
  wire       [26:0]   _zz_7375;
  wire       [35:0]   _zz_7376;
  wire       [17:0]   _zz_7377;
  wire       [35:0]   _zz_7378;
  wire       [35:0]   _zz_7379;
  wire       [35:0]   _zz_7380;
  wire       [35:0]   _zz_7381;
  wire       [35:0]   _zz_7382;
  wire       [26:0]   _zz_7383;
  wire       [35:0]   _zz_7384;
  wire       [17:0]   _zz_7385;
  wire       [35:0]   _zz_7386;
  wire       [35:0]   _zz_7387;
  wire       [35:0]   _zz_7388;
  wire       [35:0]   _zz_7389;
  wire       [35:0]   _zz_7390;
  wire       [26:0]   _zz_7391;
  wire       [35:0]   _zz_7392;
  wire       [17:0]   _zz_7393;
  wire       [35:0]   _zz_7394;
  wire       [35:0]   _zz_7395;
  wire       [35:0]   _zz_7396;
  wire       [35:0]   _zz_7397;
  wire       [35:0]   _zz_7398;
  wire       [26:0]   _zz_7399;
  wire       [35:0]   _zz_7400;
  wire       [17:0]   _zz_7401;
  wire       [17:0]   _zz_7402;
  wire       [35:0]   _zz_7403;
  wire       [35:0]   _zz_7404;
  wire       [17:0]   _zz_7405;
  wire       [35:0]   _zz_7406;
  wire       [35:0]   _zz_7407;
  wire       [35:0]   _zz_7408;
  wire       [17:0]   _zz_7409;
  wire       [35:0]   _zz_7410;
  wire       [35:0]   _zz_7411;
  wire       [35:0]   _zz_7412;
  wire       [35:0]   _zz_7413;
  wire       [35:0]   _zz_7414;
  wire       [35:0]   _zz_7415;
  wire       [26:0]   _zz_7416;
  wire       [35:0]   _zz_7417;
  wire       [17:0]   _zz_7418;
  wire       [35:0]   _zz_7419;
  wire       [35:0]   _zz_7420;
  wire       [35:0]   _zz_7421;
  wire       [35:0]   _zz_7422;
  wire       [35:0]   _zz_7423;
  wire       [26:0]   _zz_7424;
  wire       [35:0]   _zz_7425;
  wire       [17:0]   _zz_7426;
  wire       [35:0]   _zz_7427;
  wire       [35:0]   _zz_7428;
  wire       [35:0]   _zz_7429;
  wire       [35:0]   _zz_7430;
  wire       [35:0]   _zz_7431;
  wire       [26:0]   _zz_7432;
  wire       [35:0]   _zz_7433;
  wire       [17:0]   _zz_7434;
  wire       [35:0]   _zz_7435;
  wire       [35:0]   _zz_7436;
  wire       [35:0]   _zz_7437;
  wire       [35:0]   _zz_7438;
  wire       [35:0]   _zz_7439;
  wire       [26:0]   _zz_7440;
  wire       [35:0]   _zz_7441;
  wire       [17:0]   _zz_7442;
  wire       [17:0]   _zz_7443;
  wire       [35:0]   _zz_7444;
  wire       [35:0]   _zz_7445;
  wire       [17:0]   _zz_7446;
  wire       [35:0]   _zz_7447;
  wire       [35:0]   _zz_7448;
  wire       [35:0]   _zz_7449;
  wire       [17:0]   _zz_7450;
  wire       [35:0]   _zz_7451;
  wire       [35:0]   _zz_7452;
  wire       [35:0]   _zz_7453;
  wire       [35:0]   _zz_7454;
  wire       [35:0]   _zz_7455;
  wire       [35:0]   _zz_7456;
  wire       [26:0]   _zz_7457;
  wire       [35:0]   _zz_7458;
  wire       [17:0]   _zz_7459;
  wire       [35:0]   _zz_7460;
  wire       [35:0]   _zz_7461;
  wire       [35:0]   _zz_7462;
  wire       [35:0]   _zz_7463;
  wire       [35:0]   _zz_7464;
  wire       [26:0]   _zz_7465;
  wire       [35:0]   _zz_7466;
  wire       [17:0]   _zz_7467;
  wire       [35:0]   _zz_7468;
  wire       [35:0]   _zz_7469;
  wire       [35:0]   _zz_7470;
  wire       [35:0]   _zz_7471;
  wire       [35:0]   _zz_7472;
  wire       [26:0]   _zz_7473;
  wire       [35:0]   _zz_7474;
  wire       [17:0]   _zz_7475;
  wire       [35:0]   _zz_7476;
  wire       [35:0]   _zz_7477;
  wire       [35:0]   _zz_7478;
  wire       [35:0]   _zz_7479;
  wire       [35:0]   _zz_7480;
  wire       [26:0]   _zz_7481;
  wire       [35:0]   _zz_7482;
  wire       [17:0]   _zz_7483;
  wire       [17:0]   _zz_7484;
  wire       [35:0]   _zz_7485;
  wire       [35:0]   _zz_7486;
  wire       [17:0]   _zz_7487;
  wire       [35:0]   _zz_7488;
  wire       [35:0]   _zz_7489;
  wire       [35:0]   _zz_7490;
  wire       [17:0]   _zz_7491;
  wire       [35:0]   _zz_7492;
  wire       [35:0]   _zz_7493;
  wire       [35:0]   _zz_7494;
  wire       [35:0]   _zz_7495;
  wire       [35:0]   _zz_7496;
  wire       [35:0]   _zz_7497;
  wire       [26:0]   _zz_7498;
  wire       [35:0]   _zz_7499;
  wire       [17:0]   _zz_7500;
  wire       [35:0]   _zz_7501;
  wire       [35:0]   _zz_7502;
  wire       [35:0]   _zz_7503;
  wire       [35:0]   _zz_7504;
  wire       [35:0]   _zz_7505;
  wire       [26:0]   _zz_7506;
  wire       [35:0]   _zz_7507;
  wire       [17:0]   _zz_7508;
  wire       [35:0]   _zz_7509;
  wire       [35:0]   _zz_7510;
  wire       [35:0]   _zz_7511;
  wire       [35:0]   _zz_7512;
  wire       [35:0]   _zz_7513;
  wire       [26:0]   _zz_7514;
  wire       [35:0]   _zz_7515;
  wire       [17:0]   _zz_7516;
  wire       [35:0]   _zz_7517;
  wire       [35:0]   _zz_7518;
  wire       [35:0]   _zz_7519;
  wire       [35:0]   _zz_7520;
  wire       [35:0]   _zz_7521;
  wire       [26:0]   _zz_7522;
  wire       [35:0]   _zz_7523;
  wire       [17:0]   _zz_7524;
  wire       [17:0]   _zz_7525;
  wire       [35:0]   _zz_7526;
  wire       [35:0]   _zz_7527;
  wire       [17:0]   _zz_7528;
  wire       [35:0]   _zz_7529;
  wire       [35:0]   _zz_7530;
  wire       [35:0]   _zz_7531;
  wire       [17:0]   _zz_7532;
  wire       [35:0]   _zz_7533;
  wire       [35:0]   _zz_7534;
  wire       [35:0]   _zz_7535;
  wire       [35:0]   _zz_7536;
  wire       [35:0]   _zz_7537;
  wire       [35:0]   _zz_7538;
  wire       [26:0]   _zz_7539;
  wire       [35:0]   _zz_7540;
  wire       [17:0]   _zz_7541;
  wire       [35:0]   _zz_7542;
  wire       [35:0]   _zz_7543;
  wire       [35:0]   _zz_7544;
  wire       [35:0]   _zz_7545;
  wire       [35:0]   _zz_7546;
  wire       [26:0]   _zz_7547;
  wire       [35:0]   _zz_7548;
  wire       [17:0]   _zz_7549;
  wire       [35:0]   _zz_7550;
  wire       [35:0]   _zz_7551;
  wire       [35:0]   _zz_7552;
  wire       [35:0]   _zz_7553;
  wire       [35:0]   _zz_7554;
  wire       [26:0]   _zz_7555;
  wire       [35:0]   _zz_7556;
  wire       [17:0]   _zz_7557;
  wire       [35:0]   _zz_7558;
  wire       [35:0]   _zz_7559;
  wire       [35:0]   _zz_7560;
  wire       [35:0]   _zz_7561;
  wire       [35:0]   _zz_7562;
  wire       [26:0]   _zz_7563;
  wire       [35:0]   _zz_7564;
  wire       [17:0]   _zz_7565;
  wire       [17:0]   _zz_7566;
  wire       [35:0]   _zz_7567;
  wire       [35:0]   _zz_7568;
  wire       [17:0]   _zz_7569;
  wire       [35:0]   _zz_7570;
  wire       [35:0]   _zz_7571;
  wire       [35:0]   _zz_7572;
  wire       [17:0]   _zz_7573;
  wire       [35:0]   _zz_7574;
  wire       [35:0]   _zz_7575;
  wire       [35:0]   _zz_7576;
  wire       [35:0]   _zz_7577;
  wire       [35:0]   _zz_7578;
  wire       [35:0]   _zz_7579;
  wire       [26:0]   _zz_7580;
  wire       [35:0]   _zz_7581;
  wire       [17:0]   _zz_7582;
  wire       [35:0]   _zz_7583;
  wire       [35:0]   _zz_7584;
  wire       [35:0]   _zz_7585;
  wire       [35:0]   _zz_7586;
  wire       [35:0]   _zz_7587;
  wire       [26:0]   _zz_7588;
  wire       [35:0]   _zz_7589;
  wire       [17:0]   _zz_7590;
  wire       [35:0]   _zz_7591;
  wire       [35:0]   _zz_7592;
  wire       [35:0]   _zz_7593;
  wire       [35:0]   _zz_7594;
  wire       [35:0]   _zz_7595;
  wire       [26:0]   _zz_7596;
  wire       [35:0]   _zz_7597;
  wire       [17:0]   _zz_7598;
  wire       [35:0]   _zz_7599;
  wire       [35:0]   _zz_7600;
  wire       [35:0]   _zz_7601;
  wire       [35:0]   _zz_7602;
  wire       [35:0]   _zz_7603;
  wire       [26:0]   _zz_7604;
  wire       [35:0]   _zz_7605;
  wire       [17:0]   _zz_7606;
  wire       [17:0]   _zz_7607;
  wire       [35:0]   _zz_7608;
  wire       [35:0]   _zz_7609;
  wire       [17:0]   _zz_7610;
  wire       [35:0]   _zz_7611;
  wire       [35:0]   _zz_7612;
  wire       [35:0]   _zz_7613;
  wire       [17:0]   _zz_7614;
  wire       [35:0]   _zz_7615;
  wire       [35:0]   _zz_7616;
  wire       [35:0]   _zz_7617;
  wire       [35:0]   _zz_7618;
  wire       [35:0]   _zz_7619;
  wire       [35:0]   _zz_7620;
  wire       [26:0]   _zz_7621;
  wire       [35:0]   _zz_7622;
  wire       [17:0]   _zz_7623;
  wire       [35:0]   _zz_7624;
  wire       [35:0]   _zz_7625;
  wire       [35:0]   _zz_7626;
  wire       [35:0]   _zz_7627;
  wire       [35:0]   _zz_7628;
  wire       [26:0]   _zz_7629;
  wire       [35:0]   _zz_7630;
  wire       [17:0]   _zz_7631;
  wire       [35:0]   _zz_7632;
  wire       [35:0]   _zz_7633;
  wire       [35:0]   _zz_7634;
  wire       [35:0]   _zz_7635;
  wire       [35:0]   _zz_7636;
  wire       [26:0]   _zz_7637;
  wire       [35:0]   _zz_7638;
  wire       [17:0]   _zz_7639;
  wire       [35:0]   _zz_7640;
  wire       [35:0]   _zz_7641;
  wire       [35:0]   _zz_7642;
  wire       [35:0]   _zz_7643;
  wire       [35:0]   _zz_7644;
  wire       [26:0]   _zz_7645;
  wire       [35:0]   _zz_7646;
  wire       [17:0]   _zz_7647;
  wire       [17:0]   _zz_7648;
  wire       [35:0]   _zz_7649;
  wire       [35:0]   _zz_7650;
  wire       [17:0]   _zz_7651;
  wire       [35:0]   _zz_7652;
  wire       [35:0]   _zz_7653;
  wire       [35:0]   _zz_7654;
  wire       [17:0]   _zz_7655;
  wire       [35:0]   _zz_7656;
  wire       [35:0]   _zz_7657;
  wire       [35:0]   _zz_7658;
  wire       [35:0]   _zz_7659;
  wire       [35:0]   _zz_7660;
  wire       [35:0]   _zz_7661;
  wire       [26:0]   _zz_7662;
  wire       [35:0]   _zz_7663;
  wire       [17:0]   _zz_7664;
  wire       [35:0]   _zz_7665;
  wire       [35:0]   _zz_7666;
  wire       [35:0]   _zz_7667;
  wire       [35:0]   _zz_7668;
  wire       [35:0]   _zz_7669;
  wire       [26:0]   _zz_7670;
  wire       [35:0]   _zz_7671;
  wire       [17:0]   _zz_7672;
  wire       [35:0]   _zz_7673;
  wire       [35:0]   _zz_7674;
  wire       [35:0]   _zz_7675;
  wire       [35:0]   _zz_7676;
  wire       [35:0]   _zz_7677;
  wire       [26:0]   _zz_7678;
  wire       [35:0]   _zz_7679;
  wire       [17:0]   _zz_7680;
  wire       [35:0]   _zz_7681;
  wire       [35:0]   _zz_7682;
  wire       [35:0]   _zz_7683;
  wire       [35:0]   _zz_7684;
  wire       [35:0]   _zz_7685;
  wire       [26:0]   _zz_7686;
  wire       [35:0]   _zz_7687;
  wire       [17:0]   _zz_7688;
  wire       [17:0]   _zz_7689;
  wire       [35:0]   _zz_7690;
  wire       [35:0]   _zz_7691;
  wire       [17:0]   _zz_7692;
  wire       [35:0]   _zz_7693;
  wire       [35:0]   _zz_7694;
  wire       [35:0]   _zz_7695;
  wire       [17:0]   _zz_7696;
  wire       [35:0]   _zz_7697;
  wire       [35:0]   _zz_7698;
  wire       [35:0]   _zz_7699;
  wire       [35:0]   _zz_7700;
  wire       [35:0]   _zz_7701;
  wire       [35:0]   _zz_7702;
  wire       [26:0]   _zz_7703;
  wire       [35:0]   _zz_7704;
  wire       [17:0]   _zz_7705;
  wire       [35:0]   _zz_7706;
  wire       [35:0]   _zz_7707;
  wire       [35:0]   _zz_7708;
  wire       [35:0]   _zz_7709;
  wire       [35:0]   _zz_7710;
  wire       [26:0]   _zz_7711;
  wire       [35:0]   _zz_7712;
  wire       [17:0]   _zz_7713;
  wire       [35:0]   _zz_7714;
  wire       [35:0]   _zz_7715;
  wire       [35:0]   _zz_7716;
  wire       [35:0]   _zz_7717;
  wire       [35:0]   _zz_7718;
  wire       [26:0]   _zz_7719;
  wire       [35:0]   _zz_7720;
  wire       [17:0]   _zz_7721;
  wire       [35:0]   _zz_7722;
  wire       [35:0]   _zz_7723;
  wire       [35:0]   _zz_7724;
  wire       [35:0]   _zz_7725;
  wire       [35:0]   _zz_7726;
  wire       [26:0]   _zz_7727;
  wire       [35:0]   _zz_7728;
  wire       [17:0]   _zz_7729;
  wire       [17:0]   _zz_7730;
  wire       [35:0]   _zz_7731;
  wire       [35:0]   _zz_7732;
  wire       [17:0]   _zz_7733;
  wire       [35:0]   _zz_7734;
  wire       [35:0]   _zz_7735;
  wire       [35:0]   _zz_7736;
  wire       [17:0]   _zz_7737;
  wire       [35:0]   _zz_7738;
  wire       [35:0]   _zz_7739;
  wire       [35:0]   _zz_7740;
  wire       [35:0]   _zz_7741;
  wire       [35:0]   _zz_7742;
  wire       [35:0]   _zz_7743;
  wire       [26:0]   _zz_7744;
  wire       [35:0]   _zz_7745;
  wire       [17:0]   _zz_7746;
  wire       [35:0]   _zz_7747;
  wire       [35:0]   _zz_7748;
  wire       [35:0]   _zz_7749;
  wire       [35:0]   _zz_7750;
  wire       [35:0]   _zz_7751;
  wire       [26:0]   _zz_7752;
  wire       [35:0]   _zz_7753;
  wire       [17:0]   _zz_7754;
  wire       [35:0]   _zz_7755;
  wire       [35:0]   _zz_7756;
  wire       [35:0]   _zz_7757;
  wire       [35:0]   _zz_7758;
  wire       [35:0]   _zz_7759;
  wire       [26:0]   _zz_7760;
  wire       [35:0]   _zz_7761;
  wire       [17:0]   _zz_7762;
  wire       [35:0]   _zz_7763;
  wire       [35:0]   _zz_7764;
  wire       [35:0]   _zz_7765;
  wire       [35:0]   _zz_7766;
  wire       [35:0]   _zz_7767;
  wire       [26:0]   _zz_7768;
  wire       [35:0]   _zz_7769;
  wire       [17:0]   _zz_7770;
  wire       [17:0]   _zz_7771;
  wire       [35:0]   _zz_7772;
  wire       [35:0]   _zz_7773;
  wire       [17:0]   _zz_7774;
  wire       [35:0]   _zz_7775;
  wire       [35:0]   _zz_7776;
  wire       [35:0]   _zz_7777;
  wire       [17:0]   _zz_7778;
  wire       [35:0]   _zz_7779;
  wire       [35:0]   _zz_7780;
  wire       [35:0]   _zz_7781;
  wire       [35:0]   _zz_7782;
  wire       [35:0]   _zz_7783;
  wire       [35:0]   _zz_7784;
  wire       [26:0]   _zz_7785;
  wire       [35:0]   _zz_7786;
  wire       [17:0]   _zz_7787;
  wire       [35:0]   _zz_7788;
  wire       [35:0]   _zz_7789;
  wire       [35:0]   _zz_7790;
  wire       [35:0]   _zz_7791;
  wire       [35:0]   _zz_7792;
  wire       [26:0]   _zz_7793;
  wire       [35:0]   _zz_7794;
  wire       [17:0]   _zz_7795;
  wire       [35:0]   _zz_7796;
  wire       [35:0]   _zz_7797;
  wire       [35:0]   _zz_7798;
  wire       [35:0]   _zz_7799;
  wire       [35:0]   _zz_7800;
  wire       [26:0]   _zz_7801;
  wire       [35:0]   _zz_7802;
  wire       [17:0]   _zz_7803;
  wire       [35:0]   _zz_7804;
  wire       [35:0]   _zz_7805;
  wire       [35:0]   _zz_7806;
  wire       [35:0]   _zz_7807;
  wire       [35:0]   _zz_7808;
  wire       [26:0]   _zz_7809;
  wire       [35:0]   _zz_7810;
  wire       [17:0]   _zz_7811;
  wire       [17:0]   _zz_7812;
  wire       [35:0]   _zz_7813;
  wire       [35:0]   _zz_7814;
  wire       [17:0]   _zz_7815;
  wire       [35:0]   _zz_7816;
  wire       [35:0]   _zz_7817;
  wire       [35:0]   _zz_7818;
  wire       [17:0]   _zz_7819;
  wire       [35:0]   _zz_7820;
  wire       [35:0]   _zz_7821;
  wire       [35:0]   _zz_7822;
  wire       [35:0]   _zz_7823;
  wire       [35:0]   _zz_7824;
  wire       [35:0]   _zz_7825;
  wire       [26:0]   _zz_7826;
  wire       [35:0]   _zz_7827;
  wire       [17:0]   _zz_7828;
  wire       [35:0]   _zz_7829;
  wire       [35:0]   _zz_7830;
  wire       [35:0]   _zz_7831;
  wire       [35:0]   _zz_7832;
  wire       [35:0]   _zz_7833;
  wire       [26:0]   _zz_7834;
  wire       [35:0]   _zz_7835;
  wire       [17:0]   _zz_7836;
  wire       [35:0]   _zz_7837;
  wire       [35:0]   _zz_7838;
  wire       [35:0]   _zz_7839;
  wire       [35:0]   _zz_7840;
  wire       [35:0]   _zz_7841;
  wire       [26:0]   _zz_7842;
  wire       [35:0]   _zz_7843;
  wire       [17:0]   _zz_7844;
  wire       [35:0]   _zz_7845;
  wire       [35:0]   _zz_7846;
  wire       [35:0]   _zz_7847;
  wire       [35:0]   _zz_7848;
  wire       [35:0]   _zz_7849;
  wire       [26:0]   _zz_7850;
  wire       [35:0]   _zz_7851;
  wire       [17:0]   _zz_7852;
  wire       [17:0]   _zz_7853;
  wire       [35:0]   _zz_7854;
  wire       [35:0]   _zz_7855;
  wire       [17:0]   _zz_7856;
  wire       [35:0]   _zz_7857;
  wire       [35:0]   _zz_7858;
  wire       [35:0]   _zz_7859;
  wire       [17:0]   _zz_7860;
  wire       [35:0]   _zz_7861;
  wire       [35:0]   _zz_7862;
  wire       [35:0]   _zz_7863;
  wire       [35:0]   _zz_7864;
  wire       [35:0]   _zz_7865;
  wire       [35:0]   _zz_7866;
  wire       [26:0]   _zz_7867;
  wire       [35:0]   _zz_7868;
  wire       [17:0]   _zz_7869;
  wire       [35:0]   _zz_7870;
  wire       [35:0]   _zz_7871;
  wire       [35:0]   _zz_7872;
  wire       [35:0]   _zz_7873;
  wire       [35:0]   _zz_7874;
  wire       [26:0]   _zz_7875;
  wire       [35:0]   _zz_7876;
  wire       [17:0]   _zz_7877;
  wire       [35:0]   _zz_7878;
  wire       [35:0]   _zz_7879;
  wire       [35:0]   _zz_7880;
  wire       [35:0]   _zz_7881;
  wire       [35:0]   _zz_7882;
  wire       [26:0]   _zz_7883;
  wire       [35:0]   _zz_7884;
  wire       [17:0]   _zz_7885;
  wire       [35:0]   _zz_7886;
  wire       [35:0]   _zz_7887;
  wire       [35:0]   _zz_7888;
  wire       [35:0]   _zz_7889;
  wire       [35:0]   _zz_7890;
  wire       [26:0]   _zz_7891;
  wire       [35:0]   _zz_7892;
  wire       [17:0]   _zz_7893;
  wire       [17:0]   _zz_7894;
  wire       [35:0]   _zz_7895;
  wire       [35:0]   _zz_7896;
  wire       [17:0]   _zz_7897;
  wire       [35:0]   _zz_7898;
  wire       [35:0]   _zz_7899;
  wire       [35:0]   _zz_7900;
  wire       [17:0]   _zz_7901;
  wire       [35:0]   _zz_7902;
  wire       [35:0]   _zz_7903;
  wire       [35:0]   _zz_7904;
  wire       [35:0]   _zz_7905;
  wire       [35:0]   _zz_7906;
  wire       [35:0]   _zz_7907;
  wire       [26:0]   _zz_7908;
  wire       [35:0]   _zz_7909;
  wire       [17:0]   _zz_7910;
  wire       [35:0]   _zz_7911;
  wire       [35:0]   _zz_7912;
  wire       [35:0]   _zz_7913;
  wire       [35:0]   _zz_7914;
  wire       [35:0]   _zz_7915;
  wire       [26:0]   _zz_7916;
  wire       [35:0]   _zz_7917;
  wire       [17:0]   _zz_7918;
  wire       [35:0]   _zz_7919;
  wire       [35:0]   _zz_7920;
  wire       [35:0]   _zz_7921;
  wire       [35:0]   _zz_7922;
  wire       [35:0]   _zz_7923;
  wire       [26:0]   _zz_7924;
  wire       [35:0]   _zz_7925;
  wire       [17:0]   _zz_7926;
  wire       [35:0]   _zz_7927;
  wire       [35:0]   _zz_7928;
  wire       [35:0]   _zz_7929;
  wire       [35:0]   _zz_7930;
  wire       [35:0]   _zz_7931;
  wire       [26:0]   _zz_7932;
  wire       [35:0]   _zz_7933;
  wire       [17:0]   _zz_7934;
  wire       [17:0]   _zz_7935;
  wire       [35:0]   _zz_7936;
  wire       [35:0]   _zz_7937;
  wire       [17:0]   _zz_7938;
  wire       [35:0]   _zz_7939;
  wire       [35:0]   _zz_7940;
  wire       [35:0]   _zz_7941;
  wire       [17:0]   _zz_7942;
  wire       [35:0]   _zz_7943;
  wire       [35:0]   _zz_7944;
  wire       [35:0]   _zz_7945;
  wire       [35:0]   _zz_7946;
  wire       [35:0]   _zz_7947;
  wire       [35:0]   _zz_7948;
  wire       [26:0]   _zz_7949;
  wire       [35:0]   _zz_7950;
  wire       [17:0]   _zz_7951;
  wire       [35:0]   _zz_7952;
  wire       [35:0]   _zz_7953;
  wire       [35:0]   _zz_7954;
  wire       [35:0]   _zz_7955;
  wire       [35:0]   _zz_7956;
  wire       [26:0]   _zz_7957;
  wire       [35:0]   _zz_7958;
  wire       [17:0]   _zz_7959;
  wire       [35:0]   _zz_7960;
  wire       [35:0]   _zz_7961;
  wire       [35:0]   _zz_7962;
  wire       [35:0]   _zz_7963;
  wire       [35:0]   _zz_7964;
  wire       [26:0]   _zz_7965;
  wire       [35:0]   _zz_7966;
  wire       [17:0]   _zz_7967;
  wire       [35:0]   _zz_7968;
  wire       [35:0]   _zz_7969;
  wire       [35:0]   _zz_7970;
  wire       [35:0]   _zz_7971;
  wire       [35:0]   _zz_7972;
  wire       [26:0]   _zz_7973;
  wire       [35:0]   _zz_7974;
  wire       [17:0]   _zz_7975;
  wire       [17:0]   _zz_7976;
  wire       [35:0]   _zz_7977;
  wire       [35:0]   _zz_7978;
  wire       [17:0]   _zz_7979;
  wire       [35:0]   _zz_7980;
  wire       [35:0]   _zz_7981;
  wire       [35:0]   _zz_7982;
  wire       [17:0]   _zz_7983;
  wire       [35:0]   _zz_7984;
  wire       [35:0]   _zz_7985;
  wire       [35:0]   _zz_7986;
  wire       [35:0]   _zz_7987;
  wire       [35:0]   _zz_7988;
  wire       [35:0]   _zz_7989;
  wire       [26:0]   _zz_7990;
  wire       [35:0]   _zz_7991;
  wire       [17:0]   _zz_7992;
  wire       [35:0]   _zz_7993;
  wire       [35:0]   _zz_7994;
  wire       [35:0]   _zz_7995;
  wire       [35:0]   _zz_7996;
  wire       [35:0]   _zz_7997;
  wire       [26:0]   _zz_7998;
  wire       [35:0]   _zz_7999;
  wire       [17:0]   _zz_8000;
  wire       [35:0]   _zz_8001;
  wire       [35:0]   _zz_8002;
  wire       [35:0]   _zz_8003;
  wire       [35:0]   _zz_8004;
  wire       [35:0]   _zz_8005;
  wire       [26:0]   _zz_8006;
  wire       [35:0]   _zz_8007;
  wire       [17:0]   _zz_8008;
  wire       [35:0]   _zz_8009;
  wire       [35:0]   _zz_8010;
  wire       [35:0]   _zz_8011;
  wire       [35:0]   _zz_8012;
  wire       [35:0]   _zz_8013;
  wire       [26:0]   _zz_8014;
  wire       [35:0]   _zz_8015;
  wire       [17:0]   _zz_8016;
  wire       [17:0]   _zz_8017;
  wire       [35:0]   _zz_8018;
  wire       [35:0]   _zz_8019;
  wire       [17:0]   _zz_8020;
  wire       [35:0]   _zz_8021;
  wire       [35:0]   _zz_8022;
  wire       [35:0]   _zz_8023;
  wire       [17:0]   _zz_8024;
  wire       [35:0]   _zz_8025;
  wire       [35:0]   _zz_8026;
  wire       [35:0]   _zz_8027;
  wire       [35:0]   _zz_8028;
  wire       [35:0]   _zz_8029;
  wire       [35:0]   _zz_8030;
  wire       [26:0]   _zz_8031;
  wire       [35:0]   _zz_8032;
  wire       [17:0]   _zz_8033;
  wire       [35:0]   _zz_8034;
  wire       [35:0]   _zz_8035;
  wire       [35:0]   _zz_8036;
  wire       [35:0]   _zz_8037;
  wire       [35:0]   _zz_8038;
  wire       [26:0]   _zz_8039;
  wire       [35:0]   _zz_8040;
  wire       [17:0]   _zz_8041;
  wire       [35:0]   _zz_8042;
  wire       [35:0]   _zz_8043;
  wire       [35:0]   _zz_8044;
  wire       [35:0]   _zz_8045;
  wire       [35:0]   _zz_8046;
  wire       [26:0]   _zz_8047;
  wire       [35:0]   _zz_8048;
  wire       [17:0]   _zz_8049;
  wire       [35:0]   _zz_8050;
  wire       [35:0]   _zz_8051;
  wire       [35:0]   _zz_8052;
  wire       [35:0]   _zz_8053;
  wire       [35:0]   _zz_8054;
  wire       [26:0]   _zz_8055;
  wire       [35:0]   _zz_8056;
  wire       [17:0]   _zz_8057;
  wire       [17:0]   _zz_8058;
  wire       [35:0]   _zz_8059;
  wire       [35:0]   _zz_8060;
  wire       [17:0]   _zz_8061;
  wire       [35:0]   _zz_8062;
  wire       [35:0]   _zz_8063;
  wire       [35:0]   _zz_8064;
  wire       [17:0]   _zz_8065;
  wire       [35:0]   _zz_8066;
  wire       [35:0]   _zz_8067;
  wire       [35:0]   _zz_8068;
  wire       [35:0]   _zz_8069;
  wire       [35:0]   _zz_8070;
  wire       [35:0]   _zz_8071;
  wire       [26:0]   _zz_8072;
  wire       [35:0]   _zz_8073;
  wire       [17:0]   _zz_8074;
  wire       [35:0]   _zz_8075;
  wire       [35:0]   _zz_8076;
  wire       [35:0]   _zz_8077;
  wire       [35:0]   _zz_8078;
  wire       [35:0]   _zz_8079;
  wire       [26:0]   _zz_8080;
  wire       [35:0]   _zz_8081;
  wire       [17:0]   _zz_8082;
  wire       [35:0]   _zz_8083;
  wire       [35:0]   _zz_8084;
  wire       [35:0]   _zz_8085;
  wire       [35:0]   _zz_8086;
  wire       [35:0]   _zz_8087;
  wire       [26:0]   _zz_8088;
  wire       [35:0]   _zz_8089;
  wire       [17:0]   _zz_8090;
  wire       [35:0]   _zz_8091;
  wire       [35:0]   _zz_8092;
  wire       [35:0]   _zz_8093;
  wire       [35:0]   _zz_8094;
  wire       [35:0]   _zz_8095;
  wire       [26:0]   _zz_8096;
  wire       [35:0]   _zz_8097;
  wire       [17:0]   _zz_8098;
  wire       [17:0]   _zz_8099;
  wire       [35:0]   _zz_8100;
  wire       [35:0]   _zz_8101;
  wire       [17:0]   _zz_8102;
  wire       [35:0]   _zz_8103;
  wire       [35:0]   _zz_8104;
  wire       [35:0]   _zz_8105;
  wire       [17:0]   _zz_8106;
  wire       [35:0]   _zz_8107;
  wire       [35:0]   _zz_8108;
  wire       [35:0]   _zz_8109;
  wire       [35:0]   _zz_8110;
  wire       [35:0]   _zz_8111;
  wire       [35:0]   _zz_8112;
  wire       [26:0]   _zz_8113;
  wire       [35:0]   _zz_8114;
  wire       [17:0]   _zz_8115;
  wire       [35:0]   _zz_8116;
  wire       [35:0]   _zz_8117;
  wire       [35:0]   _zz_8118;
  wire       [35:0]   _zz_8119;
  wire       [35:0]   _zz_8120;
  wire       [26:0]   _zz_8121;
  wire       [35:0]   _zz_8122;
  wire       [17:0]   _zz_8123;
  wire       [35:0]   _zz_8124;
  wire       [35:0]   _zz_8125;
  wire       [35:0]   _zz_8126;
  wire       [35:0]   _zz_8127;
  wire       [35:0]   _zz_8128;
  wire       [26:0]   _zz_8129;
  wire       [35:0]   _zz_8130;
  wire       [17:0]   _zz_8131;
  wire       [35:0]   _zz_8132;
  wire       [35:0]   _zz_8133;
  wire       [35:0]   _zz_8134;
  wire       [35:0]   _zz_8135;
  wire       [35:0]   _zz_8136;
  wire       [26:0]   _zz_8137;
  wire       [35:0]   _zz_8138;
  wire       [17:0]   _zz_8139;
  wire       [17:0]   _zz_8140;
  wire       [35:0]   _zz_8141;
  wire       [35:0]   _zz_8142;
  wire       [17:0]   _zz_8143;
  wire       [35:0]   _zz_8144;
  wire       [35:0]   _zz_8145;
  wire       [35:0]   _zz_8146;
  wire       [17:0]   _zz_8147;
  wire       [35:0]   _zz_8148;
  wire       [35:0]   _zz_8149;
  wire       [35:0]   _zz_8150;
  wire       [35:0]   _zz_8151;
  wire       [35:0]   _zz_8152;
  wire       [35:0]   _zz_8153;
  wire       [26:0]   _zz_8154;
  wire       [35:0]   _zz_8155;
  wire       [17:0]   _zz_8156;
  wire       [35:0]   _zz_8157;
  wire       [35:0]   _zz_8158;
  wire       [35:0]   _zz_8159;
  wire       [35:0]   _zz_8160;
  wire       [35:0]   _zz_8161;
  wire       [26:0]   _zz_8162;
  wire       [35:0]   _zz_8163;
  wire       [17:0]   _zz_8164;
  wire       [35:0]   _zz_8165;
  wire       [35:0]   _zz_8166;
  wire       [35:0]   _zz_8167;
  wire       [35:0]   _zz_8168;
  wire       [35:0]   _zz_8169;
  wire       [26:0]   _zz_8170;
  wire       [35:0]   _zz_8171;
  wire       [17:0]   _zz_8172;
  wire       [35:0]   _zz_8173;
  wire       [35:0]   _zz_8174;
  wire       [35:0]   _zz_8175;
  wire       [35:0]   _zz_8176;
  wire       [35:0]   _zz_8177;
  wire       [26:0]   _zz_8178;
  wire       [35:0]   _zz_8179;
  wire       [17:0]   _zz_8180;
  wire       [17:0]   _zz_8181;
  wire       [35:0]   _zz_8182;
  wire       [35:0]   _zz_8183;
  wire       [17:0]   _zz_8184;
  wire       [35:0]   _zz_8185;
  wire       [35:0]   _zz_8186;
  wire       [35:0]   _zz_8187;
  wire       [17:0]   _zz_8188;
  wire       [35:0]   _zz_8189;
  wire       [35:0]   _zz_8190;
  wire       [35:0]   _zz_8191;
  wire       [35:0]   _zz_8192;
  wire       [35:0]   _zz_8193;
  wire       [35:0]   _zz_8194;
  wire       [26:0]   _zz_8195;
  wire       [35:0]   _zz_8196;
  wire       [17:0]   _zz_8197;
  wire       [35:0]   _zz_8198;
  wire       [35:0]   _zz_8199;
  wire       [35:0]   _zz_8200;
  wire       [35:0]   _zz_8201;
  wire       [35:0]   _zz_8202;
  wire       [26:0]   _zz_8203;
  wire       [35:0]   _zz_8204;
  wire       [17:0]   _zz_8205;
  wire       [35:0]   _zz_8206;
  wire       [35:0]   _zz_8207;
  wire       [35:0]   _zz_8208;
  wire       [35:0]   _zz_8209;
  wire       [35:0]   _zz_8210;
  wire       [26:0]   _zz_8211;
  wire       [35:0]   _zz_8212;
  wire       [17:0]   _zz_8213;
  wire       [35:0]   _zz_8214;
  wire       [35:0]   _zz_8215;
  wire       [35:0]   _zz_8216;
  wire       [35:0]   _zz_8217;
  wire       [35:0]   _zz_8218;
  wire       [26:0]   _zz_8219;
  wire       [35:0]   _zz_8220;
  wire       [17:0]   _zz_8221;
  wire       [17:0]   _zz_8222;
  wire       [35:0]   _zz_8223;
  wire       [35:0]   _zz_8224;
  wire       [17:0]   _zz_8225;
  wire       [35:0]   _zz_8226;
  wire       [35:0]   _zz_8227;
  wire       [35:0]   _zz_8228;
  wire       [17:0]   _zz_8229;
  wire       [35:0]   _zz_8230;
  wire       [35:0]   _zz_8231;
  wire       [35:0]   _zz_8232;
  wire       [35:0]   _zz_8233;
  wire       [35:0]   _zz_8234;
  wire       [35:0]   _zz_8235;
  wire       [26:0]   _zz_8236;
  wire       [35:0]   _zz_8237;
  wire       [17:0]   _zz_8238;
  wire       [35:0]   _zz_8239;
  wire       [35:0]   _zz_8240;
  wire       [35:0]   _zz_8241;
  wire       [35:0]   _zz_8242;
  wire       [35:0]   _zz_8243;
  wire       [26:0]   _zz_8244;
  wire       [35:0]   _zz_8245;
  wire       [17:0]   _zz_8246;
  wire       [35:0]   _zz_8247;
  wire       [35:0]   _zz_8248;
  wire       [35:0]   _zz_8249;
  wire       [35:0]   _zz_8250;
  wire       [35:0]   _zz_8251;
  wire       [26:0]   _zz_8252;
  wire       [35:0]   _zz_8253;
  wire       [17:0]   _zz_8254;
  wire       [35:0]   _zz_8255;
  wire       [35:0]   _zz_8256;
  wire       [35:0]   _zz_8257;
  wire       [35:0]   _zz_8258;
  wire       [35:0]   _zz_8259;
  wire       [26:0]   _zz_8260;
  wire       [35:0]   _zz_8261;
  wire       [17:0]   _zz_8262;
  wire       [17:0]   _zz_8263;
  wire       [35:0]   _zz_8264;
  wire       [35:0]   _zz_8265;
  wire       [17:0]   _zz_8266;
  wire       [35:0]   _zz_8267;
  wire       [35:0]   _zz_8268;
  wire       [35:0]   _zz_8269;
  wire       [17:0]   _zz_8270;
  wire       [35:0]   _zz_8271;
  wire       [35:0]   _zz_8272;
  wire       [35:0]   _zz_8273;
  wire       [35:0]   _zz_8274;
  wire       [35:0]   _zz_8275;
  wire       [35:0]   _zz_8276;
  wire       [26:0]   _zz_8277;
  wire       [35:0]   _zz_8278;
  wire       [17:0]   _zz_8279;
  wire       [35:0]   _zz_8280;
  wire       [35:0]   _zz_8281;
  wire       [35:0]   _zz_8282;
  wire       [35:0]   _zz_8283;
  wire       [35:0]   _zz_8284;
  wire       [26:0]   _zz_8285;
  wire       [35:0]   _zz_8286;
  wire       [17:0]   _zz_8287;
  wire       [35:0]   _zz_8288;
  wire       [35:0]   _zz_8289;
  wire       [35:0]   _zz_8290;
  wire       [35:0]   _zz_8291;
  wire       [35:0]   _zz_8292;
  wire       [26:0]   _zz_8293;
  wire       [35:0]   _zz_8294;
  wire       [17:0]   _zz_8295;
  wire       [35:0]   _zz_8296;
  wire       [35:0]   _zz_8297;
  wire       [35:0]   _zz_8298;
  wire       [35:0]   _zz_8299;
  wire       [35:0]   _zz_8300;
  wire       [26:0]   _zz_8301;
  wire       [35:0]   _zz_8302;
  wire       [17:0]   _zz_8303;
  wire       [17:0]   _zz_8304;
  wire       [35:0]   _zz_8305;
  wire       [35:0]   _zz_8306;
  wire       [17:0]   _zz_8307;
  wire       [35:0]   _zz_8308;
  wire       [35:0]   _zz_8309;
  wire       [35:0]   _zz_8310;
  wire       [17:0]   _zz_8311;
  wire       [35:0]   _zz_8312;
  wire       [35:0]   _zz_8313;
  wire       [35:0]   _zz_8314;
  wire       [35:0]   _zz_8315;
  wire       [35:0]   _zz_8316;
  wire       [35:0]   _zz_8317;
  wire       [26:0]   _zz_8318;
  wire       [35:0]   _zz_8319;
  wire       [17:0]   _zz_8320;
  wire       [35:0]   _zz_8321;
  wire       [35:0]   _zz_8322;
  wire       [35:0]   _zz_8323;
  wire       [35:0]   _zz_8324;
  wire       [35:0]   _zz_8325;
  wire       [26:0]   _zz_8326;
  wire       [35:0]   _zz_8327;
  wire       [17:0]   _zz_8328;
  wire       [35:0]   _zz_8329;
  wire       [35:0]   _zz_8330;
  wire       [35:0]   _zz_8331;
  wire       [35:0]   _zz_8332;
  wire       [35:0]   _zz_8333;
  wire       [26:0]   _zz_8334;
  wire       [35:0]   _zz_8335;
  wire       [17:0]   _zz_8336;
  wire       [35:0]   _zz_8337;
  wire       [35:0]   _zz_8338;
  wire       [35:0]   _zz_8339;
  wire       [35:0]   _zz_8340;
  wire       [35:0]   _zz_8341;
  wire       [26:0]   _zz_8342;
  wire       [35:0]   _zz_8343;
  wire       [17:0]   _zz_8344;
  wire       [17:0]   _zz_8345;
  wire       [35:0]   _zz_8346;
  wire       [35:0]   _zz_8347;
  wire       [17:0]   _zz_8348;
  wire       [35:0]   _zz_8349;
  wire       [35:0]   _zz_8350;
  wire       [35:0]   _zz_8351;
  wire       [17:0]   _zz_8352;
  wire       [35:0]   _zz_8353;
  wire       [35:0]   _zz_8354;
  wire       [35:0]   _zz_8355;
  wire       [35:0]   _zz_8356;
  wire       [35:0]   _zz_8357;
  wire       [35:0]   _zz_8358;
  wire       [26:0]   _zz_8359;
  wire       [35:0]   _zz_8360;
  wire       [17:0]   _zz_8361;
  wire       [35:0]   _zz_8362;
  wire       [35:0]   _zz_8363;
  wire       [35:0]   _zz_8364;
  wire       [35:0]   _zz_8365;
  wire       [35:0]   _zz_8366;
  wire       [26:0]   _zz_8367;
  wire       [35:0]   _zz_8368;
  wire       [17:0]   _zz_8369;
  wire       [35:0]   _zz_8370;
  wire       [35:0]   _zz_8371;
  wire       [35:0]   _zz_8372;
  wire       [35:0]   _zz_8373;
  wire       [35:0]   _zz_8374;
  wire       [26:0]   _zz_8375;
  wire       [35:0]   _zz_8376;
  wire       [17:0]   _zz_8377;
  wire       [35:0]   _zz_8378;
  wire       [35:0]   _zz_8379;
  wire       [35:0]   _zz_8380;
  wire       [35:0]   _zz_8381;
  wire       [35:0]   _zz_8382;
  wire       [26:0]   _zz_8383;
  wire       [35:0]   _zz_8384;
  wire       [17:0]   _zz_8385;
  wire       [17:0]   _zz_8386;
  wire       [35:0]   _zz_8387;
  wire       [35:0]   _zz_8388;
  wire       [17:0]   _zz_8389;
  wire       [35:0]   _zz_8390;
  wire       [35:0]   _zz_8391;
  wire       [35:0]   _zz_8392;
  wire       [17:0]   _zz_8393;
  wire       [35:0]   _zz_8394;
  wire       [35:0]   _zz_8395;
  wire       [35:0]   _zz_8396;
  wire       [35:0]   _zz_8397;
  wire       [35:0]   _zz_8398;
  wire       [35:0]   _zz_8399;
  wire       [26:0]   _zz_8400;
  wire       [35:0]   _zz_8401;
  wire       [17:0]   _zz_8402;
  wire       [35:0]   _zz_8403;
  wire       [35:0]   _zz_8404;
  wire       [35:0]   _zz_8405;
  wire       [35:0]   _zz_8406;
  wire       [35:0]   _zz_8407;
  wire       [26:0]   _zz_8408;
  wire       [35:0]   _zz_8409;
  wire       [17:0]   _zz_8410;
  wire       [35:0]   _zz_8411;
  wire       [35:0]   _zz_8412;
  wire       [35:0]   _zz_8413;
  wire       [35:0]   _zz_8414;
  wire       [35:0]   _zz_8415;
  wire       [26:0]   _zz_8416;
  wire       [35:0]   _zz_8417;
  wire       [17:0]   _zz_8418;
  wire       [35:0]   _zz_8419;
  wire       [35:0]   _zz_8420;
  wire       [35:0]   _zz_8421;
  wire       [35:0]   _zz_8422;
  wire       [35:0]   _zz_8423;
  wire       [26:0]   _zz_8424;
  wire       [35:0]   _zz_8425;
  wire       [17:0]   _zz_8426;
  wire       [17:0]   _zz_8427;
  wire       [35:0]   _zz_8428;
  wire       [35:0]   _zz_8429;
  wire       [17:0]   _zz_8430;
  wire       [35:0]   _zz_8431;
  wire       [35:0]   _zz_8432;
  wire       [35:0]   _zz_8433;
  wire       [17:0]   _zz_8434;
  wire       [35:0]   _zz_8435;
  wire       [35:0]   _zz_8436;
  wire       [35:0]   _zz_8437;
  wire       [35:0]   _zz_8438;
  wire       [35:0]   _zz_8439;
  wire       [35:0]   _zz_8440;
  wire       [26:0]   _zz_8441;
  wire       [35:0]   _zz_8442;
  wire       [17:0]   _zz_8443;
  wire       [35:0]   _zz_8444;
  wire       [35:0]   _zz_8445;
  wire       [35:0]   _zz_8446;
  wire       [35:0]   _zz_8447;
  wire       [35:0]   _zz_8448;
  wire       [26:0]   _zz_8449;
  wire       [35:0]   _zz_8450;
  wire       [17:0]   _zz_8451;
  wire       [35:0]   _zz_8452;
  wire       [35:0]   _zz_8453;
  wire       [35:0]   _zz_8454;
  wire       [35:0]   _zz_8455;
  wire       [35:0]   _zz_8456;
  wire       [26:0]   _zz_8457;
  wire       [35:0]   _zz_8458;
  wire       [17:0]   _zz_8459;
  wire       [35:0]   _zz_8460;
  wire       [35:0]   _zz_8461;
  wire       [35:0]   _zz_8462;
  wire       [35:0]   _zz_8463;
  wire       [35:0]   _zz_8464;
  wire       [26:0]   _zz_8465;
  wire       [35:0]   _zz_8466;
  wire       [17:0]   _zz_8467;
  wire       [17:0]   _zz_8468;
  wire       [35:0]   _zz_8469;
  wire       [35:0]   _zz_8470;
  wire       [17:0]   _zz_8471;
  wire       [35:0]   _zz_8472;
  wire       [35:0]   _zz_8473;
  wire       [35:0]   _zz_8474;
  wire       [17:0]   _zz_8475;
  wire       [35:0]   _zz_8476;
  wire       [35:0]   _zz_8477;
  wire       [35:0]   _zz_8478;
  wire       [35:0]   _zz_8479;
  wire       [35:0]   _zz_8480;
  wire       [35:0]   _zz_8481;
  wire       [26:0]   _zz_8482;
  wire       [35:0]   _zz_8483;
  wire       [17:0]   _zz_8484;
  wire       [35:0]   _zz_8485;
  wire       [35:0]   _zz_8486;
  wire       [35:0]   _zz_8487;
  wire       [35:0]   _zz_8488;
  wire       [35:0]   _zz_8489;
  wire       [26:0]   _zz_8490;
  wire       [35:0]   _zz_8491;
  wire       [17:0]   _zz_8492;
  wire       [35:0]   _zz_8493;
  wire       [35:0]   _zz_8494;
  wire       [35:0]   _zz_8495;
  wire       [35:0]   _zz_8496;
  wire       [35:0]   _zz_8497;
  wire       [26:0]   _zz_8498;
  wire       [35:0]   _zz_8499;
  wire       [17:0]   _zz_8500;
  wire       [35:0]   _zz_8501;
  wire       [35:0]   _zz_8502;
  wire       [35:0]   _zz_8503;
  wire       [35:0]   _zz_8504;
  wire       [35:0]   _zz_8505;
  wire       [26:0]   _zz_8506;
  wire       [35:0]   _zz_8507;
  wire       [17:0]   _zz_8508;
  wire       [17:0]   _zz_8509;
  wire       [35:0]   _zz_8510;
  wire       [35:0]   _zz_8511;
  wire       [17:0]   _zz_8512;
  wire       [35:0]   _zz_8513;
  wire       [35:0]   _zz_8514;
  wire       [35:0]   _zz_8515;
  wire       [17:0]   _zz_8516;
  wire       [35:0]   _zz_8517;
  wire       [35:0]   _zz_8518;
  wire       [35:0]   _zz_8519;
  wire       [35:0]   _zz_8520;
  wire       [35:0]   _zz_8521;
  wire       [35:0]   _zz_8522;
  wire       [26:0]   _zz_8523;
  wire       [35:0]   _zz_8524;
  wire       [17:0]   _zz_8525;
  wire       [35:0]   _zz_8526;
  wire       [35:0]   _zz_8527;
  wire       [35:0]   _zz_8528;
  wire       [35:0]   _zz_8529;
  wire       [35:0]   _zz_8530;
  wire       [26:0]   _zz_8531;
  wire       [35:0]   _zz_8532;
  wire       [17:0]   _zz_8533;
  wire       [35:0]   _zz_8534;
  wire       [35:0]   _zz_8535;
  wire       [35:0]   _zz_8536;
  wire       [35:0]   _zz_8537;
  wire       [35:0]   _zz_8538;
  wire       [26:0]   _zz_8539;
  wire       [35:0]   _zz_8540;
  wire       [17:0]   _zz_8541;
  wire       [35:0]   _zz_8542;
  wire       [35:0]   _zz_8543;
  wire       [35:0]   _zz_8544;
  wire       [35:0]   _zz_8545;
  wire       [35:0]   _zz_8546;
  wire       [26:0]   _zz_8547;
  wire       [35:0]   _zz_8548;
  wire       [17:0]   _zz_8549;
  wire       [17:0]   _zz_8550;
  wire       [35:0]   _zz_8551;
  wire       [35:0]   _zz_8552;
  wire       [17:0]   _zz_8553;
  wire       [35:0]   _zz_8554;
  wire       [35:0]   _zz_8555;
  wire       [35:0]   _zz_8556;
  wire       [17:0]   _zz_8557;
  wire       [35:0]   _zz_8558;
  wire       [35:0]   _zz_8559;
  wire       [35:0]   _zz_8560;
  wire       [35:0]   _zz_8561;
  wire       [35:0]   _zz_8562;
  wire       [35:0]   _zz_8563;
  wire       [26:0]   _zz_8564;
  wire       [35:0]   _zz_8565;
  wire       [17:0]   _zz_8566;
  wire       [35:0]   _zz_8567;
  wire       [35:0]   _zz_8568;
  wire       [35:0]   _zz_8569;
  wire       [35:0]   _zz_8570;
  wire       [35:0]   _zz_8571;
  wire       [26:0]   _zz_8572;
  wire       [35:0]   _zz_8573;
  wire       [17:0]   _zz_8574;
  wire       [35:0]   _zz_8575;
  wire       [35:0]   _zz_8576;
  wire       [35:0]   _zz_8577;
  wire       [35:0]   _zz_8578;
  wire       [35:0]   _zz_8579;
  wire       [26:0]   _zz_8580;
  wire       [35:0]   _zz_8581;
  wire       [17:0]   _zz_8582;
  wire       [35:0]   _zz_8583;
  wire       [35:0]   _zz_8584;
  wire       [35:0]   _zz_8585;
  wire       [35:0]   _zz_8586;
  wire       [35:0]   _zz_8587;
  wire       [26:0]   _zz_8588;
  wire       [35:0]   _zz_8589;
  wire       [17:0]   _zz_8590;
  wire       [17:0]   _zz_8591;
  wire       [35:0]   _zz_8592;
  wire       [35:0]   _zz_8593;
  wire       [17:0]   _zz_8594;
  wire       [35:0]   _zz_8595;
  wire       [35:0]   _zz_8596;
  wire       [35:0]   _zz_8597;
  wire       [17:0]   _zz_8598;
  wire       [35:0]   _zz_8599;
  wire       [35:0]   _zz_8600;
  wire       [35:0]   _zz_8601;
  wire       [35:0]   _zz_8602;
  wire       [35:0]   _zz_8603;
  wire       [35:0]   _zz_8604;
  wire       [26:0]   _zz_8605;
  wire       [35:0]   _zz_8606;
  wire       [17:0]   _zz_8607;
  wire       [35:0]   _zz_8608;
  wire       [35:0]   _zz_8609;
  wire       [35:0]   _zz_8610;
  wire       [35:0]   _zz_8611;
  wire       [35:0]   _zz_8612;
  wire       [26:0]   _zz_8613;
  wire       [35:0]   _zz_8614;
  wire       [17:0]   _zz_8615;
  wire       [35:0]   _zz_8616;
  wire       [35:0]   _zz_8617;
  wire       [35:0]   _zz_8618;
  wire       [35:0]   _zz_8619;
  wire       [35:0]   _zz_8620;
  wire       [26:0]   _zz_8621;
  wire       [35:0]   _zz_8622;
  wire       [17:0]   _zz_8623;
  wire       [35:0]   _zz_8624;
  wire       [35:0]   _zz_8625;
  wire       [35:0]   _zz_8626;
  wire       [35:0]   _zz_8627;
  wire       [35:0]   _zz_8628;
  wire       [26:0]   _zz_8629;
  wire       [35:0]   _zz_8630;
  wire       [17:0]   _zz_8631;
  wire       [17:0]   _zz_8632;
  wire       [35:0]   _zz_8633;
  wire       [35:0]   _zz_8634;
  wire       [17:0]   _zz_8635;
  wire       [35:0]   _zz_8636;
  wire       [35:0]   _zz_8637;
  wire       [35:0]   _zz_8638;
  wire       [17:0]   _zz_8639;
  wire       [35:0]   _zz_8640;
  wire       [35:0]   _zz_8641;
  wire       [35:0]   _zz_8642;
  wire       [35:0]   _zz_8643;
  wire       [35:0]   _zz_8644;
  wire       [35:0]   _zz_8645;
  wire       [26:0]   _zz_8646;
  wire       [35:0]   _zz_8647;
  wire       [17:0]   _zz_8648;
  wire       [35:0]   _zz_8649;
  wire       [35:0]   _zz_8650;
  wire       [35:0]   _zz_8651;
  wire       [35:0]   _zz_8652;
  wire       [35:0]   _zz_8653;
  wire       [26:0]   _zz_8654;
  wire       [35:0]   _zz_8655;
  wire       [17:0]   _zz_8656;
  wire       [35:0]   _zz_8657;
  wire       [35:0]   _zz_8658;
  wire       [35:0]   _zz_8659;
  wire       [35:0]   _zz_8660;
  wire       [35:0]   _zz_8661;
  wire       [26:0]   _zz_8662;
  wire       [35:0]   _zz_8663;
  wire       [17:0]   _zz_8664;
  wire       [35:0]   _zz_8665;
  wire       [35:0]   _zz_8666;
  wire       [35:0]   _zz_8667;
  wire       [35:0]   _zz_8668;
  wire       [35:0]   _zz_8669;
  wire       [26:0]   _zz_8670;
  wire       [35:0]   _zz_8671;
  wire       [17:0]   _zz_8672;
  wire       [17:0]   _zz_8673;
  wire       [35:0]   _zz_8674;
  wire       [35:0]   _zz_8675;
  wire       [17:0]   _zz_8676;
  wire       [35:0]   _zz_8677;
  wire       [35:0]   _zz_8678;
  wire       [35:0]   _zz_8679;
  wire       [17:0]   _zz_8680;
  wire       [35:0]   _zz_8681;
  wire       [35:0]   _zz_8682;
  wire       [35:0]   _zz_8683;
  wire       [35:0]   _zz_8684;
  wire       [35:0]   _zz_8685;
  wire       [35:0]   _zz_8686;
  wire       [26:0]   _zz_8687;
  wire       [35:0]   _zz_8688;
  wire       [17:0]   _zz_8689;
  wire       [35:0]   _zz_8690;
  wire       [35:0]   _zz_8691;
  wire       [35:0]   _zz_8692;
  wire       [35:0]   _zz_8693;
  wire       [35:0]   _zz_8694;
  wire       [26:0]   _zz_8695;
  wire       [35:0]   _zz_8696;
  wire       [17:0]   _zz_8697;
  wire       [35:0]   _zz_8698;
  wire       [35:0]   _zz_8699;
  wire       [35:0]   _zz_8700;
  wire       [35:0]   _zz_8701;
  wire       [35:0]   _zz_8702;
  wire       [26:0]   _zz_8703;
  wire       [35:0]   _zz_8704;
  wire       [17:0]   _zz_8705;
  wire       [35:0]   _zz_8706;
  wire       [35:0]   _zz_8707;
  wire       [35:0]   _zz_8708;
  wire       [35:0]   _zz_8709;
  wire       [35:0]   _zz_8710;
  wire       [26:0]   _zz_8711;
  wire       [35:0]   _zz_8712;
  wire       [17:0]   _zz_8713;
  wire       [17:0]   _zz_8714;
  wire       [35:0]   _zz_8715;
  wire       [35:0]   _zz_8716;
  wire       [17:0]   _zz_8717;
  wire       [35:0]   _zz_8718;
  wire       [35:0]   _zz_8719;
  wire       [35:0]   _zz_8720;
  wire       [17:0]   _zz_8721;
  wire       [35:0]   _zz_8722;
  wire       [35:0]   _zz_8723;
  wire       [35:0]   _zz_8724;
  wire       [35:0]   _zz_8725;
  wire       [35:0]   _zz_8726;
  wire       [35:0]   _zz_8727;
  wire       [26:0]   _zz_8728;
  wire       [35:0]   _zz_8729;
  wire       [17:0]   _zz_8730;
  wire       [35:0]   _zz_8731;
  wire       [35:0]   _zz_8732;
  wire       [35:0]   _zz_8733;
  wire       [35:0]   _zz_8734;
  wire       [35:0]   _zz_8735;
  wire       [26:0]   _zz_8736;
  wire       [35:0]   _zz_8737;
  wire       [17:0]   _zz_8738;
  wire       [35:0]   _zz_8739;
  wire       [35:0]   _zz_8740;
  wire       [35:0]   _zz_8741;
  wire       [35:0]   _zz_8742;
  wire       [35:0]   _zz_8743;
  wire       [26:0]   _zz_8744;
  wire       [35:0]   _zz_8745;
  wire       [17:0]   _zz_8746;
  wire       [35:0]   _zz_8747;
  wire       [35:0]   _zz_8748;
  wire       [35:0]   _zz_8749;
  wire       [35:0]   _zz_8750;
  wire       [35:0]   _zz_8751;
  wire       [26:0]   _zz_8752;
  wire       [35:0]   _zz_8753;
  wire       [17:0]   _zz_8754;
  wire       [17:0]   _zz_8755;
  wire       [35:0]   _zz_8756;
  wire       [35:0]   _zz_8757;
  wire       [17:0]   _zz_8758;
  wire       [35:0]   _zz_8759;
  wire       [35:0]   _zz_8760;
  wire       [35:0]   _zz_8761;
  wire       [17:0]   _zz_8762;
  wire       [35:0]   _zz_8763;
  wire       [35:0]   _zz_8764;
  wire       [35:0]   _zz_8765;
  wire       [35:0]   _zz_8766;
  wire       [35:0]   _zz_8767;
  wire       [35:0]   _zz_8768;
  wire       [26:0]   _zz_8769;
  wire       [35:0]   _zz_8770;
  wire       [17:0]   _zz_8771;
  wire       [35:0]   _zz_8772;
  wire       [35:0]   _zz_8773;
  wire       [35:0]   _zz_8774;
  wire       [35:0]   _zz_8775;
  wire       [35:0]   _zz_8776;
  wire       [26:0]   _zz_8777;
  wire       [35:0]   _zz_8778;
  wire       [17:0]   _zz_8779;
  wire       [35:0]   _zz_8780;
  wire       [35:0]   _zz_8781;
  wire       [35:0]   _zz_8782;
  wire       [35:0]   _zz_8783;
  wire       [35:0]   _zz_8784;
  wire       [26:0]   _zz_8785;
  wire       [35:0]   _zz_8786;
  wire       [17:0]   _zz_8787;
  wire       [35:0]   _zz_8788;
  wire       [35:0]   _zz_8789;
  wire       [35:0]   _zz_8790;
  wire       [35:0]   _zz_8791;
  wire       [35:0]   _zz_8792;
  wire       [26:0]   _zz_8793;
  wire       [35:0]   _zz_8794;
  wire       [17:0]   _zz_8795;
  wire       [17:0]   _zz_8796;
  wire       [35:0]   _zz_8797;
  wire       [35:0]   _zz_8798;
  wire       [17:0]   _zz_8799;
  wire       [35:0]   _zz_8800;
  wire       [35:0]   _zz_8801;
  wire       [35:0]   _zz_8802;
  wire       [17:0]   _zz_8803;
  wire       [35:0]   _zz_8804;
  wire       [35:0]   _zz_8805;
  wire       [35:0]   _zz_8806;
  wire       [35:0]   _zz_8807;
  wire       [35:0]   _zz_8808;
  wire       [35:0]   _zz_8809;
  wire       [26:0]   _zz_8810;
  wire       [35:0]   _zz_8811;
  wire       [17:0]   _zz_8812;
  wire       [35:0]   _zz_8813;
  wire       [35:0]   _zz_8814;
  wire       [35:0]   _zz_8815;
  wire       [35:0]   _zz_8816;
  wire       [35:0]   _zz_8817;
  wire       [26:0]   _zz_8818;
  wire       [35:0]   _zz_8819;
  wire       [17:0]   _zz_8820;
  wire       [35:0]   _zz_8821;
  wire       [35:0]   _zz_8822;
  wire       [35:0]   _zz_8823;
  wire       [35:0]   _zz_8824;
  wire       [35:0]   _zz_8825;
  wire       [26:0]   _zz_8826;
  wire       [35:0]   _zz_8827;
  wire       [17:0]   _zz_8828;
  wire       [35:0]   _zz_8829;
  wire       [35:0]   _zz_8830;
  wire       [35:0]   _zz_8831;
  wire       [35:0]   _zz_8832;
  wire       [35:0]   _zz_8833;
  wire       [26:0]   _zz_8834;
  wire       [35:0]   _zz_8835;
  wire       [17:0]   _zz_8836;
  wire       [17:0]   _zz_8837;
  wire       [35:0]   _zz_8838;
  wire       [35:0]   _zz_8839;
  wire       [17:0]   _zz_8840;
  wire       [35:0]   _zz_8841;
  wire       [35:0]   _zz_8842;
  wire       [35:0]   _zz_8843;
  wire       [17:0]   _zz_8844;
  wire       [35:0]   _zz_8845;
  wire       [35:0]   _zz_8846;
  wire       [35:0]   _zz_8847;
  wire       [35:0]   _zz_8848;
  wire       [35:0]   _zz_8849;
  wire       [35:0]   _zz_8850;
  wire       [26:0]   _zz_8851;
  wire       [35:0]   _zz_8852;
  wire       [17:0]   _zz_8853;
  wire       [35:0]   _zz_8854;
  wire       [35:0]   _zz_8855;
  wire       [35:0]   _zz_8856;
  wire       [35:0]   _zz_8857;
  wire       [35:0]   _zz_8858;
  wire       [26:0]   _zz_8859;
  wire       [35:0]   _zz_8860;
  wire       [17:0]   _zz_8861;
  wire       [35:0]   _zz_8862;
  wire       [35:0]   _zz_8863;
  wire       [35:0]   _zz_8864;
  wire       [35:0]   _zz_8865;
  wire       [35:0]   _zz_8866;
  wire       [26:0]   _zz_8867;
  wire       [35:0]   _zz_8868;
  wire       [17:0]   _zz_8869;
  wire       [35:0]   _zz_8870;
  wire       [35:0]   _zz_8871;
  wire       [35:0]   _zz_8872;
  wire       [35:0]   _zz_8873;
  wire       [35:0]   _zz_8874;
  wire       [26:0]   _zz_8875;
  wire       [35:0]   _zz_8876;
  wire       [17:0]   _zz_8877;
  wire       [17:0]   _zz_8878;
  wire       [35:0]   _zz_8879;
  wire       [35:0]   _zz_8880;
  wire       [17:0]   _zz_8881;
  wire       [35:0]   _zz_8882;
  wire       [35:0]   _zz_8883;
  wire       [35:0]   _zz_8884;
  wire       [17:0]   _zz_8885;
  wire       [35:0]   _zz_8886;
  wire       [35:0]   _zz_8887;
  wire       [35:0]   _zz_8888;
  wire       [35:0]   _zz_8889;
  wire       [35:0]   _zz_8890;
  wire       [35:0]   _zz_8891;
  wire       [26:0]   _zz_8892;
  wire       [35:0]   _zz_8893;
  wire       [17:0]   _zz_8894;
  wire       [35:0]   _zz_8895;
  wire       [35:0]   _zz_8896;
  wire       [35:0]   _zz_8897;
  wire       [35:0]   _zz_8898;
  wire       [35:0]   _zz_8899;
  wire       [26:0]   _zz_8900;
  wire       [35:0]   _zz_8901;
  wire       [17:0]   _zz_8902;
  wire       [35:0]   _zz_8903;
  wire       [35:0]   _zz_8904;
  wire       [35:0]   _zz_8905;
  wire       [35:0]   _zz_8906;
  wire       [35:0]   _zz_8907;
  wire       [26:0]   _zz_8908;
  wire       [35:0]   _zz_8909;
  wire       [17:0]   _zz_8910;
  wire       [35:0]   _zz_8911;
  wire       [35:0]   _zz_8912;
  wire       [35:0]   _zz_8913;
  wire       [35:0]   _zz_8914;
  wire       [35:0]   _zz_8915;
  wire       [26:0]   _zz_8916;
  wire       [35:0]   _zz_8917;
  wire       [17:0]   _zz_8918;
  wire       [17:0]   _zz_8919;
  wire       [35:0]   _zz_8920;
  wire       [35:0]   _zz_8921;
  wire       [17:0]   _zz_8922;
  wire       [35:0]   _zz_8923;
  wire       [35:0]   _zz_8924;
  wire       [35:0]   _zz_8925;
  wire       [17:0]   _zz_8926;
  wire       [35:0]   _zz_8927;
  wire       [35:0]   _zz_8928;
  wire       [35:0]   _zz_8929;
  wire       [35:0]   _zz_8930;
  wire       [35:0]   _zz_8931;
  wire       [35:0]   _zz_8932;
  wire       [26:0]   _zz_8933;
  wire       [35:0]   _zz_8934;
  wire       [17:0]   _zz_8935;
  wire       [35:0]   _zz_8936;
  wire       [35:0]   _zz_8937;
  wire       [35:0]   _zz_8938;
  wire       [35:0]   _zz_8939;
  wire       [35:0]   _zz_8940;
  wire       [26:0]   _zz_8941;
  wire       [35:0]   _zz_8942;
  wire       [17:0]   _zz_8943;
  wire       [35:0]   _zz_8944;
  wire       [35:0]   _zz_8945;
  wire       [35:0]   _zz_8946;
  wire       [35:0]   _zz_8947;
  wire       [35:0]   _zz_8948;
  wire       [26:0]   _zz_8949;
  wire       [35:0]   _zz_8950;
  wire       [17:0]   _zz_8951;
  wire       [35:0]   _zz_8952;
  wire       [35:0]   _zz_8953;
  wire       [35:0]   _zz_8954;
  wire       [35:0]   _zz_8955;
  wire       [35:0]   _zz_8956;
  wire       [26:0]   _zz_8957;
  wire       [35:0]   _zz_8958;
  wire       [17:0]   _zz_8959;
  wire       [17:0]   _zz_8960;
  wire       [35:0]   _zz_8961;
  wire       [35:0]   _zz_8962;
  wire       [17:0]   _zz_8963;
  wire       [35:0]   _zz_8964;
  wire       [35:0]   _zz_8965;
  wire       [35:0]   _zz_8966;
  wire       [17:0]   _zz_8967;
  wire       [35:0]   _zz_8968;
  wire       [35:0]   _zz_8969;
  wire       [35:0]   _zz_8970;
  wire       [35:0]   _zz_8971;
  wire       [35:0]   _zz_8972;
  wire       [35:0]   _zz_8973;
  wire       [26:0]   _zz_8974;
  wire       [35:0]   _zz_8975;
  wire       [17:0]   _zz_8976;
  wire       [35:0]   _zz_8977;
  wire       [35:0]   _zz_8978;
  wire       [35:0]   _zz_8979;
  wire       [35:0]   _zz_8980;
  wire       [35:0]   _zz_8981;
  wire       [26:0]   _zz_8982;
  wire       [35:0]   _zz_8983;
  wire       [17:0]   _zz_8984;
  wire       [35:0]   _zz_8985;
  wire       [35:0]   _zz_8986;
  wire       [35:0]   _zz_8987;
  wire       [35:0]   _zz_8988;
  wire       [35:0]   _zz_8989;
  wire       [26:0]   _zz_8990;
  wire       [35:0]   _zz_8991;
  wire       [17:0]   _zz_8992;
  wire       [35:0]   _zz_8993;
  wire       [35:0]   _zz_8994;
  wire       [35:0]   _zz_8995;
  wire       [35:0]   _zz_8996;
  wire       [35:0]   _zz_8997;
  wire       [26:0]   _zz_8998;
  wire       [35:0]   _zz_8999;
  wire       [17:0]   _zz_9000;
  wire       [17:0]   _zz_9001;
  wire       [35:0]   _zz_9002;
  wire       [35:0]   _zz_9003;
  wire       [17:0]   _zz_9004;
  wire       [35:0]   _zz_9005;
  wire       [35:0]   _zz_9006;
  wire       [35:0]   _zz_9007;
  wire       [17:0]   _zz_9008;
  wire       [35:0]   _zz_9009;
  wire       [35:0]   _zz_9010;
  wire       [35:0]   _zz_9011;
  wire       [35:0]   _zz_9012;
  wire       [35:0]   _zz_9013;
  wire       [35:0]   _zz_9014;
  wire       [26:0]   _zz_9015;
  wire       [35:0]   _zz_9016;
  wire       [17:0]   _zz_9017;
  wire       [35:0]   _zz_9018;
  wire       [35:0]   _zz_9019;
  wire       [35:0]   _zz_9020;
  wire       [35:0]   _zz_9021;
  wire       [35:0]   _zz_9022;
  wire       [26:0]   _zz_9023;
  wire       [35:0]   _zz_9024;
  wire       [17:0]   _zz_9025;
  wire       [35:0]   _zz_9026;
  wire       [35:0]   _zz_9027;
  wire       [35:0]   _zz_9028;
  wire       [35:0]   _zz_9029;
  wire       [35:0]   _zz_9030;
  wire       [26:0]   _zz_9031;
  wire       [35:0]   _zz_9032;
  wire       [17:0]   _zz_9033;
  wire       [35:0]   _zz_9034;
  wire       [35:0]   _zz_9035;
  wire       [35:0]   _zz_9036;
  wire       [35:0]   _zz_9037;
  wire       [35:0]   _zz_9038;
  wire       [26:0]   _zz_9039;
  wire       [35:0]   _zz_9040;
  wire       [17:0]   _zz_9041;
  wire       [17:0]   _zz_9042;
  wire       [35:0]   _zz_9043;
  wire       [35:0]   _zz_9044;
  wire       [17:0]   _zz_9045;
  wire       [35:0]   _zz_9046;
  wire       [35:0]   _zz_9047;
  wire       [35:0]   _zz_9048;
  wire       [17:0]   _zz_9049;
  wire       [35:0]   _zz_9050;
  wire       [35:0]   _zz_9051;
  wire       [35:0]   _zz_9052;
  wire       [35:0]   _zz_9053;
  wire       [35:0]   _zz_9054;
  wire       [35:0]   _zz_9055;
  wire       [26:0]   _zz_9056;
  wire       [35:0]   _zz_9057;
  wire       [17:0]   _zz_9058;
  wire       [35:0]   _zz_9059;
  wire       [35:0]   _zz_9060;
  wire       [35:0]   _zz_9061;
  wire       [35:0]   _zz_9062;
  wire       [35:0]   _zz_9063;
  wire       [26:0]   _zz_9064;
  wire       [35:0]   _zz_9065;
  wire       [17:0]   _zz_9066;
  wire       [35:0]   _zz_9067;
  wire       [35:0]   _zz_9068;
  wire       [35:0]   _zz_9069;
  wire       [35:0]   _zz_9070;
  wire       [35:0]   _zz_9071;
  wire       [26:0]   _zz_9072;
  wire       [35:0]   _zz_9073;
  wire       [17:0]   _zz_9074;
  wire       [35:0]   _zz_9075;
  wire       [35:0]   _zz_9076;
  wire       [35:0]   _zz_9077;
  wire       [35:0]   _zz_9078;
  wire       [35:0]   _zz_9079;
  wire       [26:0]   _zz_9080;
  wire       [35:0]   _zz_9081;
  wire       [17:0]   _zz_9082;
  wire       [17:0]   _zz_9083;
  wire       [35:0]   _zz_9084;
  wire       [35:0]   _zz_9085;
  wire       [17:0]   _zz_9086;
  wire       [35:0]   _zz_9087;
  wire       [35:0]   _zz_9088;
  wire       [35:0]   _zz_9089;
  wire       [17:0]   _zz_9090;
  wire       [35:0]   _zz_9091;
  wire       [35:0]   _zz_9092;
  wire       [35:0]   _zz_9093;
  wire       [35:0]   _zz_9094;
  wire       [35:0]   _zz_9095;
  wire       [35:0]   _zz_9096;
  wire       [26:0]   _zz_9097;
  wire       [35:0]   _zz_9098;
  wire       [17:0]   _zz_9099;
  wire       [35:0]   _zz_9100;
  wire       [35:0]   _zz_9101;
  wire       [35:0]   _zz_9102;
  wire       [35:0]   _zz_9103;
  wire       [35:0]   _zz_9104;
  wire       [26:0]   _zz_9105;
  wire       [35:0]   _zz_9106;
  wire       [17:0]   _zz_9107;
  wire       [35:0]   _zz_9108;
  wire       [35:0]   _zz_9109;
  wire       [35:0]   _zz_9110;
  wire       [35:0]   _zz_9111;
  wire       [35:0]   _zz_9112;
  wire       [26:0]   _zz_9113;
  wire       [35:0]   _zz_9114;
  wire       [17:0]   _zz_9115;
  wire       [35:0]   _zz_9116;
  wire       [35:0]   _zz_9117;
  wire       [35:0]   _zz_9118;
  wire       [35:0]   _zz_9119;
  wire       [35:0]   _zz_9120;
  wire       [26:0]   _zz_9121;
  wire       [35:0]   _zz_9122;
  wire       [17:0]   _zz_9123;
  wire       [17:0]   _zz_9124;
  wire       [35:0]   _zz_9125;
  wire       [35:0]   _zz_9126;
  wire       [17:0]   _zz_9127;
  wire       [35:0]   _zz_9128;
  wire       [35:0]   _zz_9129;
  wire       [35:0]   _zz_9130;
  wire       [17:0]   _zz_9131;
  wire       [35:0]   _zz_9132;
  wire       [35:0]   _zz_9133;
  wire       [35:0]   _zz_9134;
  wire       [35:0]   _zz_9135;
  wire       [35:0]   _zz_9136;
  wire       [35:0]   _zz_9137;
  wire       [26:0]   _zz_9138;
  wire       [35:0]   _zz_9139;
  wire       [17:0]   _zz_9140;
  wire       [35:0]   _zz_9141;
  wire       [35:0]   _zz_9142;
  wire       [35:0]   _zz_9143;
  wire       [35:0]   _zz_9144;
  wire       [35:0]   _zz_9145;
  wire       [26:0]   _zz_9146;
  wire       [35:0]   _zz_9147;
  wire       [17:0]   _zz_9148;
  wire       [35:0]   _zz_9149;
  wire       [35:0]   _zz_9150;
  wire       [35:0]   _zz_9151;
  wire       [35:0]   _zz_9152;
  wire       [35:0]   _zz_9153;
  wire       [26:0]   _zz_9154;
  wire       [35:0]   _zz_9155;
  wire       [17:0]   _zz_9156;
  wire       [35:0]   _zz_9157;
  wire       [35:0]   _zz_9158;
  wire       [35:0]   _zz_9159;
  wire       [35:0]   _zz_9160;
  wire       [35:0]   _zz_9161;
  wire       [26:0]   _zz_9162;
  wire       [35:0]   _zz_9163;
  wire       [17:0]   _zz_9164;
  wire       [17:0]   _zz_9165;
  wire       [35:0]   _zz_9166;
  wire       [35:0]   _zz_9167;
  wire       [17:0]   _zz_9168;
  wire       [35:0]   _zz_9169;
  wire       [35:0]   _zz_9170;
  wire       [35:0]   _zz_9171;
  wire       [17:0]   _zz_9172;
  wire       [35:0]   _zz_9173;
  wire       [35:0]   _zz_9174;
  wire       [35:0]   _zz_9175;
  wire       [35:0]   _zz_9176;
  wire       [35:0]   _zz_9177;
  wire       [35:0]   _zz_9178;
  wire       [26:0]   _zz_9179;
  wire       [35:0]   _zz_9180;
  wire       [17:0]   _zz_9181;
  wire       [35:0]   _zz_9182;
  wire       [35:0]   _zz_9183;
  wire       [35:0]   _zz_9184;
  wire       [35:0]   _zz_9185;
  wire       [35:0]   _zz_9186;
  wire       [26:0]   _zz_9187;
  wire       [35:0]   _zz_9188;
  wire       [17:0]   _zz_9189;
  wire       [35:0]   _zz_9190;
  wire       [35:0]   _zz_9191;
  wire       [35:0]   _zz_9192;
  wire       [35:0]   _zz_9193;
  wire       [35:0]   _zz_9194;
  wire       [26:0]   _zz_9195;
  wire       [35:0]   _zz_9196;
  wire       [17:0]   _zz_9197;
  wire       [35:0]   _zz_9198;
  wire       [35:0]   _zz_9199;
  wire       [35:0]   _zz_9200;
  wire       [35:0]   _zz_9201;
  wire       [35:0]   _zz_9202;
  wire       [26:0]   _zz_9203;
  wire       [35:0]   _zz_9204;
  wire       [17:0]   _zz_9205;
  wire       [17:0]   _zz_9206;
  wire       [35:0]   _zz_9207;
  wire       [35:0]   _zz_9208;
  wire       [17:0]   _zz_9209;
  wire       [35:0]   _zz_9210;
  wire       [35:0]   _zz_9211;
  wire       [35:0]   _zz_9212;
  wire       [17:0]   _zz_9213;
  wire       [35:0]   _zz_9214;
  wire       [35:0]   _zz_9215;
  wire       [35:0]   _zz_9216;
  wire       [35:0]   _zz_9217;
  wire       [35:0]   _zz_9218;
  wire       [35:0]   _zz_9219;
  wire       [26:0]   _zz_9220;
  wire       [35:0]   _zz_9221;
  wire       [17:0]   _zz_9222;
  wire       [35:0]   _zz_9223;
  wire       [35:0]   _zz_9224;
  wire       [35:0]   _zz_9225;
  wire       [35:0]   _zz_9226;
  wire       [35:0]   _zz_9227;
  wire       [26:0]   _zz_9228;
  wire       [35:0]   _zz_9229;
  wire       [17:0]   _zz_9230;
  wire       [35:0]   _zz_9231;
  wire       [35:0]   _zz_9232;
  wire       [35:0]   _zz_9233;
  wire       [35:0]   _zz_9234;
  wire       [35:0]   _zz_9235;
  wire       [26:0]   _zz_9236;
  wire       [35:0]   _zz_9237;
  wire       [17:0]   _zz_9238;
  wire       [35:0]   _zz_9239;
  wire       [35:0]   _zz_9240;
  wire       [35:0]   _zz_9241;
  wire       [35:0]   _zz_9242;
  wire       [35:0]   _zz_9243;
  wire       [26:0]   _zz_9244;
  wire       [35:0]   _zz_9245;
  wire       [17:0]   _zz_9246;
  wire       [17:0]   _zz_9247;
  wire       [35:0]   _zz_9248;
  wire       [35:0]   _zz_9249;
  wire       [17:0]   _zz_9250;
  wire       [35:0]   _zz_9251;
  wire       [35:0]   _zz_9252;
  wire       [35:0]   _zz_9253;
  wire       [17:0]   _zz_9254;
  wire       [35:0]   _zz_9255;
  wire       [35:0]   _zz_9256;
  wire       [35:0]   _zz_9257;
  wire       [35:0]   _zz_9258;
  wire       [35:0]   _zz_9259;
  wire       [35:0]   _zz_9260;
  wire       [26:0]   _zz_9261;
  wire       [35:0]   _zz_9262;
  wire       [17:0]   _zz_9263;
  wire       [35:0]   _zz_9264;
  wire       [35:0]   _zz_9265;
  wire       [35:0]   _zz_9266;
  wire       [35:0]   _zz_9267;
  wire       [35:0]   _zz_9268;
  wire       [26:0]   _zz_9269;
  wire       [35:0]   _zz_9270;
  wire       [17:0]   _zz_9271;
  wire       [35:0]   _zz_9272;
  wire       [35:0]   _zz_9273;
  wire       [35:0]   _zz_9274;
  wire       [35:0]   _zz_9275;
  wire       [35:0]   _zz_9276;
  wire       [26:0]   _zz_9277;
  wire       [35:0]   _zz_9278;
  wire       [17:0]   _zz_9279;
  wire       [35:0]   _zz_9280;
  wire       [35:0]   _zz_9281;
  wire       [35:0]   _zz_9282;
  wire       [35:0]   _zz_9283;
  wire       [35:0]   _zz_9284;
  wire       [26:0]   _zz_9285;
  wire       [35:0]   _zz_9286;
  wire       [17:0]   _zz_9287;
  wire       [17:0]   _zz_9288;
  wire       [35:0]   _zz_9289;
  wire       [35:0]   _zz_9290;
  wire       [17:0]   _zz_9291;
  wire       [35:0]   _zz_9292;
  wire       [35:0]   _zz_9293;
  wire       [35:0]   _zz_9294;
  wire       [17:0]   _zz_9295;
  wire       [35:0]   _zz_9296;
  wire       [35:0]   _zz_9297;
  wire       [35:0]   _zz_9298;
  wire       [35:0]   _zz_9299;
  wire       [35:0]   _zz_9300;
  wire       [35:0]   _zz_9301;
  wire       [26:0]   _zz_9302;
  wire       [35:0]   _zz_9303;
  wire       [17:0]   _zz_9304;
  wire       [35:0]   _zz_9305;
  wire       [35:0]   _zz_9306;
  wire       [35:0]   _zz_9307;
  wire       [35:0]   _zz_9308;
  wire       [35:0]   _zz_9309;
  wire       [26:0]   _zz_9310;
  wire       [35:0]   _zz_9311;
  wire       [17:0]   _zz_9312;
  wire       [35:0]   _zz_9313;
  wire       [35:0]   _zz_9314;
  wire       [35:0]   _zz_9315;
  wire       [35:0]   _zz_9316;
  wire       [35:0]   _zz_9317;
  wire       [26:0]   _zz_9318;
  wire       [35:0]   _zz_9319;
  wire       [17:0]   _zz_9320;
  wire       [35:0]   _zz_9321;
  wire       [35:0]   _zz_9322;
  wire       [35:0]   _zz_9323;
  wire       [35:0]   _zz_9324;
  wire       [35:0]   _zz_9325;
  wire       [26:0]   _zz_9326;
  wire       [35:0]   _zz_9327;
  wire       [17:0]   _zz_9328;
  wire       [17:0]   _zz_9329;
  wire       [35:0]   _zz_9330;
  wire       [35:0]   _zz_9331;
  wire       [17:0]   _zz_9332;
  wire       [35:0]   _zz_9333;
  wire       [35:0]   _zz_9334;
  wire       [35:0]   _zz_9335;
  wire       [17:0]   _zz_9336;
  wire       [35:0]   _zz_9337;
  wire       [35:0]   _zz_9338;
  wire       [35:0]   _zz_9339;
  wire       [35:0]   _zz_9340;
  wire       [35:0]   _zz_9341;
  wire       [35:0]   _zz_9342;
  wire       [26:0]   _zz_9343;
  wire       [35:0]   _zz_9344;
  wire       [17:0]   _zz_9345;
  wire       [35:0]   _zz_9346;
  wire       [35:0]   _zz_9347;
  wire       [35:0]   _zz_9348;
  wire       [35:0]   _zz_9349;
  wire       [35:0]   _zz_9350;
  wire       [26:0]   _zz_9351;
  wire       [35:0]   _zz_9352;
  wire       [17:0]   _zz_9353;
  wire       [35:0]   _zz_9354;
  wire       [35:0]   _zz_9355;
  wire       [35:0]   _zz_9356;
  wire       [35:0]   _zz_9357;
  wire       [35:0]   _zz_9358;
  wire       [26:0]   _zz_9359;
  wire       [35:0]   _zz_9360;
  wire       [17:0]   _zz_9361;
  wire       [35:0]   _zz_9362;
  wire       [35:0]   _zz_9363;
  wire       [35:0]   _zz_9364;
  wire       [35:0]   _zz_9365;
  wire       [35:0]   _zz_9366;
  wire       [26:0]   _zz_9367;
  wire       [35:0]   _zz_9368;
  wire       [17:0]   _zz_9369;
  wire       [17:0]   _zz_9370;
  wire       [35:0]   _zz_9371;
  wire       [35:0]   _zz_9372;
  wire       [17:0]   _zz_9373;
  wire       [35:0]   _zz_9374;
  wire       [35:0]   _zz_9375;
  wire       [35:0]   _zz_9376;
  wire       [17:0]   _zz_9377;
  wire       [35:0]   _zz_9378;
  wire       [35:0]   _zz_9379;
  wire       [35:0]   _zz_9380;
  wire       [35:0]   _zz_9381;
  wire       [35:0]   _zz_9382;
  wire       [35:0]   _zz_9383;
  wire       [26:0]   _zz_9384;
  wire       [35:0]   _zz_9385;
  wire       [17:0]   _zz_9386;
  wire       [35:0]   _zz_9387;
  wire       [35:0]   _zz_9388;
  wire       [35:0]   _zz_9389;
  wire       [35:0]   _zz_9390;
  wire       [35:0]   _zz_9391;
  wire       [26:0]   _zz_9392;
  wire       [35:0]   _zz_9393;
  wire       [17:0]   _zz_9394;
  wire       [35:0]   _zz_9395;
  wire       [35:0]   _zz_9396;
  wire       [35:0]   _zz_9397;
  wire       [35:0]   _zz_9398;
  wire       [35:0]   _zz_9399;
  wire       [26:0]   _zz_9400;
  wire       [35:0]   _zz_9401;
  wire       [17:0]   _zz_9402;
  wire       [35:0]   _zz_9403;
  wire       [35:0]   _zz_9404;
  wire       [35:0]   _zz_9405;
  wire       [35:0]   _zz_9406;
  wire       [35:0]   _zz_9407;
  wire       [26:0]   _zz_9408;
  wire       [35:0]   _zz_9409;
  wire       [17:0]   _zz_9410;
  wire       [17:0]   _zz_9411;
  wire       [35:0]   _zz_9412;
  wire       [35:0]   _zz_9413;
  wire       [17:0]   _zz_9414;
  wire       [35:0]   _zz_9415;
  wire       [35:0]   _zz_9416;
  wire       [35:0]   _zz_9417;
  wire       [17:0]   _zz_9418;
  wire       [35:0]   _zz_9419;
  wire       [35:0]   _zz_9420;
  wire       [35:0]   _zz_9421;
  wire       [35:0]   _zz_9422;
  wire       [35:0]   _zz_9423;
  wire       [35:0]   _zz_9424;
  wire       [26:0]   _zz_9425;
  wire       [35:0]   _zz_9426;
  wire       [17:0]   _zz_9427;
  wire       [35:0]   _zz_9428;
  wire       [35:0]   _zz_9429;
  wire       [35:0]   _zz_9430;
  wire       [35:0]   _zz_9431;
  wire       [35:0]   _zz_9432;
  wire       [26:0]   _zz_9433;
  wire       [35:0]   _zz_9434;
  wire       [17:0]   _zz_9435;
  wire       [35:0]   _zz_9436;
  wire       [35:0]   _zz_9437;
  wire       [35:0]   _zz_9438;
  wire       [35:0]   _zz_9439;
  wire       [35:0]   _zz_9440;
  wire       [26:0]   _zz_9441;
  wire       [35:0]   _zz_9442;
  wire       [17:0]   _zz_9443;
  wire       [35:0]   _zz_9444;
  wire       [35:0]   _zz_9445;
  wire       [35:0]   _zz_9446;
  wire       [35:0]   _zz_9447;
  wire       [35:0]   _zz_9448;
  wire       [26:0]   _zz_9449;
  wire       [35:0]   _zz_9450;
  wire       [17:0]   _zz_9451;
  wire       [17:0]   _zz_9452;
  wire       [35:0]   _zz_9453;
  wire       [35:0]   _zz_9454;
  wire       [17:0]   _zz_9455;
  wire       [35:0]   _zz_9456;
  wire       [35:0]   _zz_9457;
  wire       [35:0]   _zz_9458;
  wire       [17:0]   _zz_9459;
  wire       [35:0]   _zz_9460;
  wire       [35:0]   _zz_9461;
  wire       [35:0]   _zz_9462;
  wire       [35:0]   _zz_9463;
  wire       [35:0]   _zz_9464;
  wire       [35:0]   _zz_9465;
  wire       [26:0]   _zz_9466;
  wire       [35:0]   _zz_9467;
  wire       [17:0]   _zz_9468;
  wire       [35:0]   _zz_9469;
  wire       [35:0]   _zz_9470;
  wire       [35:0]   _zz_9471;
  wire       [35:0]   _zz_9472;
  wire       [35:0]   _zz_9473;
  wire       [26:0]   _zz_9474;
  wire       [35:0]   _zz_9475;
  wire       [17:0]   _zz_9476;
  wire       [35:0]   _zz_9477;
  wire       [35:0]   _zz_9478;
  wire       [35:0]   _zz_9479;
  wire       [35:0]   _zz_9480;
  wire       [35:0]   _zz_9481;
  wire       [26:0]   _zz_9482;
  wire       [35:0]   _zz_9483;
  wire       [17:0]   _zz_9484;
  wire       [35:0]   _zz_9485;
  wire       [35:0]   _zz_9486;
  wire       [35:0]   _zz_9487;
  wire       [35:0]   _zz_9488;
  wire       [35:0]   _zz_9489;
  wire       [26:0]   _zz_9490;
  wire       [35:0]   _zz_9491;
  wire       [17:0]   _zz_9492;
  wire       [17:0]   _zz_9493;
  wire       [35:0]   _zz_9494;
  wire       [35:0]   _zz_9495;
  wire       [17:0]   _zz_9496;
  wire       [35:0]   _zz_9497;
  wire       [35:0]   _zz_9498;
  wire       [35:0]   _zz_9499;
  wire       [17:0]   _zz_9500;
  wire       [35:0]   _zz_9501;
  wire       [35:0]   _zz_9502;
  wire       [35:0]   _zz_9503;
  wire       [35:0]   _zz_9504;
  wire       [35:0]   _zz_9505;
  wire       [35:0]   _zz_9506;
  wire       [26:0]   _zz_9507;
  wire       [35:0]   _zz_9508;
  wire       [17:0]   _zz_9509;
  wire       [35:0]   _zz_9510;
  wire       [35:0]   _zz_9511;
  wire       [35:0]   _zz_9512;
  wire       [35:0]   _zz_9513;
  wire       [35:0]   _zz_9514;
  wire       [26:0]   _zz_9515;
  wire       [35:0]   _zz_9516;
  wire       [17:0]   _zz_9517;
  wire       [35:0]   _zz_9518;
  wire       [35:0]   _zz_9519;
  wire       [35:0]   _zz_9520;
  wire       [35:0]   _zz_9521;
  wire       [35:0]   _zz_9522;
  wire       [26:0]   _zz_9523;
  wire       [35:0]   _zz_9524;
  wire       [17:0]   _zz_9525;
  wire       [35:0]   _zz_9526;
  wire       [35:0]   _zz_9527;
  wire       [35:0]   _zz_9528;
  wire       [35:0]   _zz_9529;
  wire       [35:0]   _zz_9530;
  wire       [26:0]   _zz_9531;
  wire       [35:0]   _zz_9532;
  wire       [17:0]   _zz_9533;
  wire       [17:0]   _zz_9534;
  wire       [35:0]   _zz_9535;
  wire       [35:0]   _zz_9536;
  wire       [17:0]   _zz_9537;
  wire       [35:0]   _zz_9538;
  wire       [35:0]   _zz_9539;
  wire       [35:0]   _zz_9540;
  wire       [17:0]   _zz_9541;
  wire       [35:0]   _zz_9542;
  wire       [35:0]   _zz_9543;
  wire       [35:0]   _zz_9544;
  wire       [35:0]   _zz_9545;
  wire       [35:0]   _zz_9546;
  wire       [35:0]   _zz_9547;
  wire       [26:0]   _zz_9548;
  wire       [35:0]   _zz_9549;
  wire       [17:0]   _zz_9550;
  wire       [35:0]   _zz_9551;
  wire       [35:0]   _zz_9552;
  wire       [35:0]   _zz_9553;
  wire       [35:0]   _zz_9554;
  wire       [35:0]   _zz_9555;
  wire       [26:0]   _zz_9556;
  wire       [35:0]   _zz_9557;
  wire       [17:0]   _zz_9558;
  wire       [35:0]   _zz_9559;
  wire       [35:0]   _zz_9560;
  wire       [35:0]   _zz_9561;
  wire       [35:0]   _zz_9562;
  wire       [35:0]   _zz_9563;
  wire       [26:0]   _zz_9564;
  wire       [35:0]   _zz_9565;
  wire       [17:0]   _zz_9566;
  wire       [35:0]   _zz_9567;
  wire       [35:0]   _zz_9568;
  wire       [35:0]   _zz_9569;
  wire       [35:0]   _zz_9570;
  wire       [35:0]   _zz_9571;
  wire       [26:0]   _zz_9572;
  wire       [35:0]   _zz_9573;
  wire       [17:0]   _zz_9574;
  wire       [17:0]   _zz_9575;
  wire       [35:0]   _zz_9576;
  wire       [35:0]   _zz_9577;
  wire       [17:0]   _zz_9578;
  wire       [35:0]   _zz_9579;
  wire       [35:0]   _zz_9580;
  wire       [35:0]   _zz_9581;
  wire       [17:0]   _zz_9582;
  wire       [35:0]   _zz_9583;
  wire       [35:0]   _zz_9584;
  wire       [35:0]   _zz_9585;
  wire       [35:0]   _zz_9586;
  wire       [35:0]   _zz_9587;
  wire       [35:0]   _zz_9588;
  wire       [26:0]   _zz_9589;
  wire       [35:0]   _zz_9590;
  wire       [17:0]   _zz_9591;
  wire       [35:0]   _zz_9592;
  wire       [35:0]   _zz_9593;
  wire       [35:0]   _zz_9594;
  wire       [35:0]   _zz_9595;
  wire       [35:0]   _zz_9596;
  wire       [26:0]   _zz_9597;
  wire       [35:0]   _zz_9598;
  wire       [17:0]   _zz_9599;
  wire       [35:0]   _zz_9600;
  wire       [35:0]   _zz_9601;
  wire       [35:0]   _zz_9602;
  wire       [35:0]   _zz_9603;
  wire       [35:0]   _zz_9604;
  wire       [26:0]   _zz_9605;
  wire       [35:0]   _zz_9606;
  wire       [17:0]   _zz_9607;
  wire       [35:0]   _zz_9608;
  wire       [35:0]   _zz_9609;
  wire       [35:0]   _zz_9610;
  wire       [35:0]   _zz_9611;
  wire       [35:0]   _zz_9612;
  wire       [26:0]   _zz_9613;
  wire       [35:0]   _zz_9614;
  wire       [17:0]   _zz_9615;
  wire       [17:0]   _zz_9616;
  wire       [35:0]   _zz_9617;
  wire       [35:0]   _zz_9618;
  wire       [17:0]   _zz_9619;
  wire       [35:0]   _zz_9620;
  wire       [35:0]   _zz_9621;
  wire       [35:0]   _zz_9622;
  wire       [17:0]   _zz_9623;
  wire       [35:0]   _zz_9624;
  wire       [35:0]   _zz_9625;
  wire       [35:0]   _zz_9626;
  wire       [35:0]   _zz_9627;
  wire       [35:0]   _zz_9628;
  wire       [35:0]   _zz_9629;
  wire       [26:0]   _zz_9630;
  wire       [35:0]   _zz_9631;
  wire       [17:0]   _zz_9632;
  wire       [35:0]   _zz_9633;
  wire       [35:0]   _zz_9634;
  wire       [35:0]   _zz_9635;
  wire       [35:0]   _zz_9636;
  wire       [35:0]   _zz_9637;
  wire       [26:0]   _zz_9638;
  wire       [35:0]   _zz_9639;
  wire       [17:0]   _zz_9640;
  wire       [35:0]   _zz_9641;
  wire       [35:0]   _zz_9642;
  wire       [35:0]   _zz_9643;
  wire       [35:0]   _zz_9644;
  wire       [35:0]   _zz_9645;
  wire       [26:0]   _zz_9646;
  wire       [35:0]   _zz_9647;
  wire       [17:0]   _zz_9648;
  wire       [35:0]   _zz_9649;
  wire       [35:0]   _zz_9650;
  wire       [35:0]   _zz_9651;
  wire       [35:0]   _zz_9652;
  wire       [35:0]   _zz_9653;
  wire       [26:0]   _zz_9654;
  wire       [35:0]   _zz_9655;
  wire       [17:0]   _zz_9656;
  wire       [17:0]   _zz_9657;
  wire       [35:0]   _zz_9658;
  wire       [35:0]   _zz_9659;
  wire       [17:0]   _zz_9660;
  wire       [35:0]   _zz_9661;
  wire       [35:0]   _zz_9662;
  wire       [35:0]   _zz_9663;
  wire       [17:0]   _zz_9664;
  wire       [35:0]   _zz_9665;
  wire       [35:0]   _zz_9666;
  wire       [35:0]   _zz_9667;
  wire       [35:0]   _zz_9668;
  wire       [35:0]   _zz_9669;
  wire       [35:0]   _zz_9670;
  wire       [26:0]   _zz_9671;
  wire       [35:0]   _zz_9672;
  wire       [17:0]   _zz_9673;
  wire       [35:0]   _zz_9674;
  wire       [35:0]   _zz_9675;
  wire       [35:0]   _zz_9676;
  wire       [35:0]   _zz_9677;
  wire       [35:0]   _zz_9678;
  wire       [26:0]   _zz_9679;
  wire       [35:0]   _zz_9680;
  wire       [17:0]   _zz_9681;
  wire       [35:0]   _zz_9682;
  wire       [35:0]   _zz_9683;
  wire       [35:0]   _zz_9684;
  wire       [35:0]   _zz_9685;
  wire       [35:0]   _zz_9686;
  wire       [26:0]   _zz_9687;
  wire       [35:0]   _zz_9688;
  wire       [17:0]   _zz_9689;
  wire       [35:0]   _zz_9690;
  wire       [35:0]   _zz_9691;
  wire       [35:0]   _zz_9692;
  wire       [35:0]   _zz_9693;
  wire       [35:0]   _zz_9694;
  wire       [26:0]   _zz_9695;
  wire       [35:0]   _zz_9696;
  wire       [17:0]   _zz_9697;
  wire       [17:0]   _zz_9698;
  wire       [35:0]   _zz_9699;
  wire       [35:0]   _zz_9700;
  wire       [17:0]   _zz_9701;
  wire       [35:0]   _zz_9702;
  wire       [35:0]   _zz_9703;
  wire       [35:0]   _zz_9704;
  wire       [17:0]   _zz_9705;
  wire       [35:0]   _zz_9706;
  wire       [35:0]   _zz_9707;
  wire       [35:0]   _zz_9708;
  wire       [35:0]   _zz_9709;
  wire       [35:0]   _zz_9710;
  wire       [35:0]   _zz_9711;
  wire       [26:0]   _zz_9712;
  wire       [35:0]   _zz_9713;
  wire       [17:0]   _zz_9714;
  wire       [35:0]   _zz_9715;
  wire       [35:0]   _zz_9716;
  wire       [35:0]   _zz_9717;
  wire       [35:0]   _zz_9718;
  wire       [35:0]   _zz_9719;
  wire       [26:0]   _zz_9720;
  wire       [35:0]   _zz_9721;
  wire       [17:0]   _zz_9722;
  wire       [35:0]   _zz_9723;
  wire       [35:0]   _zz_9724;
  wire       [35:0]   _zz_9725;
  wire       [35:0]   _zz_9726;
  wire       [35:0]   _zz_9727;
  wire       [26:0]   _zz_9728;
  wire       [35:0]   _zz_9729;
  wire       [17:0]   _zz_9730;
  wire       [35:0]   _zz_9731;
  wire       [35:0]   _zz_9732;
  wire       [35:0]   _zz_9733;
  wire       [35:0]   _zz_9734;
  wire       [35:0]   _zz_9735;
  wire       [26:0]   _zz_9736;
  wire       [35:0]   _zz_9737;
  wire       [17:0]   _zz_9738;
  wire       [17:0]   _zz_9739;
  wire       [35:0]   _zz_9740;
  wire       [35:0]   _zz_9741;
  wire       [17:0]   _zz_9742;
  wire       [35:0]   _zz_9743;
  wire       [35:0]   _zz_9744;
  wire       [35:0]   _zz_9745;
  wire       [17:0]   _zz_9746;
  wire       [35:0]   _zz_9747;
  wire       [35:0]   _zz_9748;
  wire       [35:0]   _zz_9749;
  wire       [35:0]   _zz_9750;
  wire       [35:0]   _zz_9751;
  wire       [35:0]   _zz_9752;
  wire       [26:0]   _zz_9753;
  wire       [35:0]   _zz_9754;
  wire       [17:0]   _zz_9755;
  wire       [35:0]   _zz_9756;
  wire       [35:0]   _zz_9757;
  wire       [35:0]   _zz_9758;
  wire       [35:0]   _zz_9759;
  wire       [35:0]   _zz_9760;
  wire       [26:0]   _zz_9761;
  wire       [35:0]   _zz_9762;
  wire       [17:0]   _zz_9763;
  wire       [35:0]   _zz_9764;
  wire       [35:0]   _zz_9765;
  wire       [35:0]   _zz_9766;
  wire       [35:0]   _zz_9767;
  wire       [35:0]   _zz_9768;
  wire       [26:0]   _zz_9769;
  wire       [35:0]   _zz_9770;
  wire       [17:0]   _zz_9771;
  wire       [35:0]   _zz_9772;
  wire       [35:0]   _zz_9773;
  wire       [35:0]   _zz_9774;
  wire       [35:0]   _zz_9775;
  wire       [35:0]   _zz_9776;
  wire       [26:0]   _zz_9777;
  wire       [35:0]   _zz_9778;
  wire       [17:0]   _zz_9779;
  wire       [17:0]   _zz_9780;
  wire       [35:0]   _zz_9781;
  wire       [35:0]   _zz_9782;
  wire       [17:0]   _zz_9783;
  wire       [35:0]   _zz_9784;
  wire       [35:0]   _zz_9785;
  wire       [35:0]   _zz_9786;
  wire       [17:0]   _zz_9787;
  wire       [35:0]   _zz_9788;
  wire       [35:0]   _zz_9789;
  wire       [35:0]   _zz_9790;
  wire       [35:0]   _zz_9791;
  wire       [35:0]   _zz_9792;
  wire       [35:0]   _zz_9793;
  wire       [26:0]   _zz_9794;
  wire       [35:0]   _zz_9795;
  wire       [17:0]   _zz_9796;
  wire       [35:0]   _zz_9797;
  wire       [35:0]   _zz_9798;
  wire       [35:0]   _zz_9799;
  wire       [35:0]   _zz_9800;
  wire       [35:0]   _zz_9801;
  wire       [26:0]   _zz_9802;
  wire       [35:0]   _zz_9803;
  wire       [17:0]   _zz_9804;
  wire       [35:0]   _zz_9805;
  wire       [35:0]   _zz_9806;
  wire       [35:0]   _zz_9807;
  wire       [35:0]   _zz_9808;
  wire       [35:0]   _zz_9809;
  wire       [26:0]   _zz_9810;
  wire       [35:0]   _zz_9811;
  wire       [17:0]   _zz_9812;
  wire       [35:0]   _zz_9813;
  wire       [35:0]   _zz_9814;
  wire       [35:0]   _zz_9815;
  wire       [35:0]   _zz_9816;
  wire       [35:0]   _zz_9817;
  wire       [26:0]   _zz_9818;
  wire       [35:0]   _zz_9819;
  wire       [17:0]   _zz_9820;
  wire       [17:0]   _zz_9821;
  wire       [35:0]   _zz_9822;
  wire       [35:0]   _zz_9823;
  wire       [17:0]   _zz_9824;
  wire       [35:0]   _zz_9825;
  wire       [35:0]   _zz_9826;
  wire       [35:0]   _zz_9827;
  wire       [17:0]   _zz_9828;
  wire       [35:0]   _zz_9829;
  wire       [35:0]   _zz_9830;
  wire       [35:0]   _zz_9831;
  wire       [35:0]   _zz_9832;
  wire       [35:0]   _zz_9833;
  wire       [35:0]   _zz_9834;
  wire       [26:0]   _zz_9835;
  wire       [35:0]   _zz_9836;
  wire       [17:0]   _zz_9837;
  wire       [35:0]   _zz_9838;
  wire       [35:0]   _zz_9839;
  wire       [35:0]   _zz_9840;
  wire       [35:0]   _zz_9841;
  wire       [35:0]   _zz_9842;
  wire       [26:0]   _zz_9843;
  wire       [35:0]   _zz_9844;
  wire       [17:0]   _zz_9845;
  wire       [35:0]   _zz_9846;
  wire       [35:0]   _zz_9847;
  wire       [35:0]   _zz_9848;
  wire       [35:0]   _zz_9849;
  wire       [35:0]   _zz_9850;
  wire       [26:0]   _zz_9851;
  wire       [35:0]   _zz_9852;
  wire       [17:0]   _zz_9853;
  wire       [35:0]   _zz_9854;
  wire       [35:0]   _zz_9855;
  wire       [35:0]   _zz_9856;
  wire       [35:0]   _zz_9857;
  wire       [35:0]   _zz_9858;
  wire       [26:0]   _zz_9859;
  wire       [35:0]   _zz_9860;
  wire       [17:0]   _zz_9861;
  wire       [17:0]   _zz_9862;
  wire       [35:0]   _zz_9863;
  wire       [35:0]   _zz_9864;
  wire       [17:0]   _zz_9865;
  wire       [35:0]   _zz_9866;
  wire       [35:0]   _zz_9867;
  wire       [35:0]   _zz_9868;
  wire       [17:0]   _zz_9869;
  wire       [35:0]   _zz_9870;
  wire       [35:0]   _zz_9871;
  wire       [35:0]   _zz_9872;
  wire       [35:0]   _zz_9873;
  wire       [35:0]   _zz_9874;
  wire       [35:0]   _zz_9875;
  wire       [26:0]   _zz_9876;
  wire       [35:0]   _zz_9877;
  wire       [17:0]   _zz_9878;
  wire       [35:0]   _zz_9879;
  wire       [35:0]   _zz_9880;
  wire       [35:0]   _zz_9881;
  wire       [35:0]   _zz_9882;
  wire       [35:0]   _zz_9883;
  wire       [26:0]   _zz_9884;
  wire       [35:0]   _zz_9885;
  wire       [17:0]   _zz_9886;
  wire       [35:0]   _zz_9887;
  wire       [35:0]   _zz_9888;
  wire       [35:0]   _zz_9889;
  wire       [35:0]   _zz_9890;
  wire       [35:0]   _zz_9891;
  wire       [26:0]   _zz_9892;
  wire       [35:0]   _zz_9893;
  wire       [17:0]   _zz_9894;
  wire       [35:0]   _zz_9895;
  wire       [35:0]   _zz_9896;
  wire       [35:0]   _zz_9897;
  wire       [35:0]   _zz_9898;
  wire       [35:0]   _zz_9899;
  wire       [26:0]   _zz_9900;
  wire       [35:0]   _zz_9901;
  wire       [17:0]   _zz_9902;
  wire       [17:0]   _zz_9903;
  wire       [35:0]   _zz_9904;
  wire       [35:0]   _zz_9905;
  wire       [17:0]   _zz_9906;
  wire       [35:0]   _zz_9907;
  wire       [35:0]   _zz_9908;
  wire       [35:0]   _zz_9909;
  wire       [17:0]   _zz_9910;
  wire       [35:0]   _zz_9911;
  wire       [35:0]   _zz_9912;
  wire       [35:0]   _zz_9913;
  wire       [35:0]   _zz_9914;
  wire       [35:0]   _zz_9915;
  wire       [35:0]   _zz_9916;
  wire       [26:0]   _zz_9917;
  wire       [35:0]   _zz_9918;
  wire       [17:0]   _zz_9919;
  wire       [35:0]   _zz_9920;
  wire       [35:0]   _zz_9921;
  wire       [35:0]   _zz_9922;
  wire       [35:0]   _zz_9923;
  wire       [35:0]   _zz_9924;
  wire       [26:0]   _zz_9925;
  wire       [35:0]   _zz_9926;
  wire       [17:0]   _zz_9927;
  wire       [35:0]   _zz_9928;
  wire       [35:0]   _zz_9929;
  wire       [35:0]   _zz_9930;
  wire       [35:0]   _zz_9931;
  wire       [35:0]   _zz_9932;
  wire       [26:0]   _zz_9933;
  wire       [35:0]   _zz_9934;
  wire       [17:0]   _zz_9935;
  wire       [35:0]   _zz_9936;
  wire       [35:0]   _zz_9937;
  wire       [35:0]   _zz_9938;
  wire       [35:0]   _zz_9939;
  wire       [35:0]   _zz_9940;
  wire       [26:0]   _zz_9941;
  wire       [35:0]   _zz_9942;
  wire       [17:0]   _zz_9943;
  wire       [17:0]   _zz_9944;
  wire       [35:0]   _zz_9945;
  wire       [35:0]   _zz_9946;
  wire       [17:0]   _zz_9947;
  wire       [35:0]   _zz_9948;
  wire       [35:0]   _zz_9949;
  wire       [35:0]   _zz_9950;
  wire       [17:0]   _zz_9951;
  wire       [35:0]   _zz_9952;
  wire       [35:0]   _zz_9953;
  wire       [35:0]   _zz_9954;
  wire       [35:0]   _zz_9955;
  wire       [35:0]   _zz_9956;
  wire       [35:0]   _zz_9957;
  wire       [26:0]   _zz_9958;
  wire       [35:0]   _zz_9959;
  wire       [17:0]   _zz_9960;
  wire       [35:0]   _zz_9961;
  wire       [35:0]   _zz_9962;
  wire       [35:0]   _zz_9963;
  wire       [35:0]   _zz_9964;
  wire       [35:0]   _zz_9965;
  wire       [26:0]   _zz_9966;
  wire       [35:0]   _zz_9967;
  wire       [17:0]   _zz_9968;
  wire       [35:0]   _zz_9969;
  wire       [35:0]   _zz_9970;
  wire       [35:0]   _zz_9971;
  wire       [35:0]   _zz_9972;
  wire       [35:0]   _zz_9973;
  wire       [26:0]   _zz_9974;
  wire       [35:0]   _zz_9975;
  wire       [17:0]   _zz_9976;
  wire       [35:0]   _zz_9977;
  wire       [35:0]   _zz_9978;
  wire       [35:0]   _zz_9979;
  wire       [35:0]   _zz_9980;
  wire       [35:0]   _zz_9981;
  wire       [26:0]   _zz_9982;
  wire       [35:0]   _zz_9983;
  wire       [17:0]   _zz_9984;
  reg        [17:0]   data_in_0_real;
  reg        [17:0]   data_in_0_imag;
  reg        [17:0]   data_in_1_real;
  reg        [17:0]   data_in_1_imag;
  reg        [17:0]   data_in_2_real;
  reg        [17:0]   data_in_2_imag;
  reg        [17:0]   data_in_3_real;
  reg        [17:0]   data_in_3_imag;
  reg        [17:0]   data_in_4_real;
  reg        [17:0]   data_in_4_imag;
  reg        [17:0]   data_in_5_real;
  reg        [17:0]   data_in_5_imag;
  reg        [17:0]   data_in_6_real;
  reg        [17:0]   data_in_6_imag;
  reg        [17:0]   data_in_7_real;
  reg        [17:0]   data_in_7_imag;
  reg        [17:0]   data_in_8_real;
  reg        [17:0]   data_in_8_imag;
  reg        [17:0]   data_in_9_real;
  reg        [17:0]   data_in_9_imag;
  reg        [17:0]   data_in_10_real;
  reg        [17:0]   data_in_10_imag;
  reg        [17:0]   data_in_11_real;
  reg        [17:0]   data_in_11_imag;
  reg        [17:0]   data_in_12_real;
  reg        [17:0]   data_in_12_imag;
  reg        [17:0]   data_in_13_real;
  reg        [17:0]   data_in_13_imag;
  reg        [17:0]   data_in_14_real;
  reg        [17:0]   data_in_14_imag;
  reg        [17:0]   data_in_15_real;
  reg        [17:0]   data_in_15_imag;
  reg        [17:0]   data_in_16_real;
  reg        [17:0]   data_in_16_imag;
  reg        [17:0]   data_in_17_real;
  reg        [17:0]   data_in_17_imag;
  reg        [17:0]   data_in_18_real;
  reg        [17:0]   data_in_18_imag;
  reg        [17:0]   data_in_19_real;
  reg        [17:0]   data_in_19_imag;
  reg        [17:0]   data_in_20_real;
  reg        [17:0]   data_in_20_imag;
  reg        [17:0]   data_in_21_real;
  reg        [17:0]   data_in_21_imag;
  reg        [17:0]   data_in_22_real;
  reg        [17:0]   data_in_22_imag;
  reg        [17:0]   data_in_23_real;
  reg        [17:0]   data_in_23_imag;
  reg        [17:0]   data_in_24_real;
  reg        [17:0]   data_in_24_imag;
  reg        [17:0]   data_in_25_real;
  reg        [17:0]   data_in_25_imag;
  reg        [17:0]   data_in_26_real;
  reg        [17:0]   data_in_26_imag;
  reg        [17:0]   data_in_27_real;
  reg        [17:0]   data_in_27_imag;
  reg        [17:0]   data_in_28_real;
  reg        [17:0]   data_in_28_imag;
  reg        [17:0]   data_in_29_real;
  reg        [17:0]   data_in_29_imag;
  reg        [17:0]   data_in_30_real;
  reg        [17:0]   data_in_30_imag;
  reg        [17:0]   data_in_31_real;
  reg        [17:0]   data_in_31_imag;
  reg        [17:0]   data_in_32_real;
  reg        [17:0]   data_in_32_imag;
  reg        [17:0]   data_in_33_real;
  reg        [17:0]   data_in_33_imag;
  reg        [17:0]   data_in_34_real;
  reg        [17:0]   data_in_34_imag;
  reg        [17:0]   data_in_35_real;
  reg        [17:0]   data_in_35_imag;
  reg        [17:0]   data_in_36_real;
  reg        [17:0]   data_in_36_imag;
  reg        [17:0]   data_in_37_real;
  reg        [17:0]   data_in_37_imag;
  reg        [17:0]   data_in_38_real;
  reg        [17:0]   data_in_38_imag;
  reg        [17:0]   data_in_39_real;
  reg        [17:0]   data_in_39_imag;
  reg        [17:0]   data_in_40_real;
  reg        [17:0]   data_in_40_imag;
  reg        [17:0]   data_in_41_real;
  reg        [17:0]   data_in_41_imag;
  reg        [17:0]   data_in_42_real;
  reg        [17:0]   data_in_42_imag;
  reg        [17:0]   data_in_43_real;
  reg        [17:0]   data_in_43_imag;
  reg        [17:0]   data_in_44_real;
  reg        [17:0]   data_in_44_imag;
  reg        [17:0]   data_in_45_real;
  reg        [17:0]   data_in_45_imag;
  reg        [17:0]   data_in_46_real;
  reg        [17:0]   data_in_46_imag;
  reg        [17:0]   data_in_47_real;
  reg        [17:0]   data_in_47_imag;
  reg        [17:0]   data_in_48_real;
  reg        [17:0]   data_in_48_imag;
  reg        [17:0]   data_in_49_real;
  reg        [17:0]   data_in_49_imag;
  reg        [17:0]   data_in_50_real;
  reg        [17:0]   data_in_50_imag;
  reg        [17:0]   data_in_51_real;
  reg        [17:0]   data_in_51_imag;
  reg        [17:0]   data_in_52_real;
  reg        [17:0]   data_in_52_imag;
  reg        [17:0]   data_in_53_real;
  reg        [17:0]   data_in_53_imag;
  reg        [17:0]   data_in_54_real;
  reg        [17:0]   data_in_54_imag;
  reg        [17:0]   data_in_55_real;
  reg        [17:0]   data_in_55_imag;
  reg        [17:0]   data_in_56_real;
  reg        [17:0]   data_in_56_imag;
  reg        [17:0]   data_in_57_real;
  reg        [17:0]   data_in_57_imag;
  reg        [17:0]   data_in_58_real;
  reg        [17:0]   data_in_58_imag;
  reg        [17:0]   data_in_59_real;
  reg        [17:0]   data_in_59_imag;
  reg        [17:0]   data_in_60_real;
  reg        [17:0]   data_in_60_imag;
  reg        [17:0]   data_in_61_real;
  reg        [17:0]   data_in_61_imag;
  reg        [17:0]   data_in_62_real;
  reg        [17:0]   data_in_62_imag;
  reg        [17:0]   data_in_63_real;
  reg        [17:0]   data_in_63_imag;
  wire       [17:0]   twiddle_factor_table_0_real;
  wire       [17:0]   twiddle_factor_table_0_imag;
  wire       [17:0]   twiddle_factor_table_1_real;
  wire       [17:0]   twiddle_factor_table_1_imag;
  wire       [17:0]   twiddle_factor_table_2_real;
  wire       [17:0]   twiddle_factor_table_2_imag;
  wire       [17:0]   twiddle_factor_table_3_real;
  wire       [17:0]   twiddle_factor_table_3_imag;
  wire       [17:0]   twiddle_factor_table_4_real;
  wire       [17:0]   twiddle_factor_table_4_imag;
  wire       [17:0]   twiddle_factor_table_5_real;
  wire       [17:0]   twiddle_factor_table_5_imag;
  wire       [17:0]   twiddle_factor_table_6_real;
  wire       [17:0]   twiddle_factor_table_6_imag;
  wire       [17:0]   twiddle_factor_table_7_real;
  wire       [17:0]   twiddle_factor_table_7_imag;
  wire       [17:0]   twiddle_factor_table_8_real;
  wire       [17:0]   twiddle_factor_table_8_imag;
  wire       [17:0]   twiddle_factor_table_9_real;
  wire       [17:0]   twiddle_factor_table_9_imag;
  wire       [17:0]   twiddle_factor_table_10_real;
  wire       [17:0]   twiddle_factor_table_10_imag;
  wire       [17:0]   twiddle_factor_table_11_real;
  wire       [17:0]   twiddle_factor_table_11_imag;
  wire       [17:0]   twiddle_factor_table_12_real;
  wire       [17:0]   twiddle_factor_table_12_imag;
  wire       [17:0]   twiddle_factor_table_13_real;
  wire       [17:0]   twiddle_factor_table_13_imag;
  wire       [17:0]   twiddle_factor_table_14_real;
  wire       [17:0]   twiddle_factor_table_14_imag;
  wire       [17:0]   twiddle_factor_table_15_real;
  wire       [17:0]   twiddle_factor_table_15_imag;
  wire       [17:0]   twiddle_factor_table_16_real;
  wire       [17:0]   twiddle_factor_table_16_imag;
  wire       [17:0]   twiddle_factor_table_17_real;
  wire       [17:0]   twiddle_factor_table_17_imag;
  wire       [17:0]   twiddle_factor_table_18_real;
  wire       [17:0]   twiddle_factor_table_18_imag;
  wire       [17:0]   twiddle_factor_table_19_real;
  wire       [17:0]   twiddle_factor_table_19_imag;
  wire       [17:0]   twiddle_factor_table_20_real;
  wire       [17:0]   twiddle_factor_table_20_imag;
  wire       [17:0]   twiddle_factor_table_21_real;
  wire       [17:0]   twiddle_factor_table_21_imag;
  wire       [17:0]   twiddle_factor_table_22_real;
  wire       [17:0]   twiddle_factor_table_22_imag;
  wire       [17:0]   twiddle_factor_table_23_real;
  wire       [17:0]   twiddle_factor_table_23_imag;
  wire       [17:0]   twiddle_factor_table_24_real;
  wire       [17:0]   twiddle_factor_table_24_imag;
  wire       [17:0]   twiddle_factor_table_25_real;
  wire       [17:0]   twiddle_factor_table_25_imag;
  wire       [17:0]   twiddle_factor_table_26_real;
  wire       [17:0]   twiddle_factor_table_26_imag;
  wire       [17:0]   twiddle_factor_table_27_real;
  wire       [17:0]   twiddle_factor_table_27_imag;
  wire       [17:0]   twiddle_factor_table_28_real;
  wire       [17:0]   twiddle_factor_table_28_imag;
  wire       [17:0]   twiddle_factor_table_29_real;
  wire       [17:0]   twiddle_factor_table_29_imag;
  wire       [17:0]   twiddle_factor_table_30_real;
  wire       [17:0]   twiddle_factor_table_30_imag;
  wire       [17:0]   twiddle_factor_table_31_real;
  wire       [17:0]   twiddle_factor_table_31_imag;
  wire       [17:0]   twiddle_factor_table_32_real;
  wire       [17:0]   twiddle_factor_table_32_imag;
  wire       [17:0]   twiddle_factor_table_33_real;
  wire       [17:0]   twiddle_factor_table_33_imag;
  wire       [17:0]   twiddle_factor_table_34_real;
  wire       [17:0]   twiddle_factor_table_34_imag;
  wire       [17:0]   twiddle_factor_table_35_real;
  wire       [17:0]   twiddle_factor_table_35_imag;
  wire       [17:0]   twiddle_factor_table_36_real;
  wire       [17:0]   twiddle_factor_table_36_imag;
  wire       [17:0]   twiddle_factor_table_37_real;
  wire       [17:0]   twiddle_factor_table_37_imag;
  wire       [17:0]   twiddle_factor_table_38_real;
  wire       [17:0]   twiddle_factor_table_38_imag;
  wire       [17:0]   twiddle_factor_table_39_real;
  wire       [17:0]   twiddle_factor_table_39_imag;
  wire       [17:0]   twiddle_factor_table_40_real;
  wire       [17:0]   twiddle_factor_table_40_imag;
  wire       [17:0]   twiddle_factor_table_41_real;
  wire       [17:0]   twiddle_factor_table_41_imag;
  wire       [17:0]   twiddle_factor_table_42_real;
  wire       [17:0]   twiddle_factor_table_42_imag;
  wire       [17:0]   twiddle_factor_table_43_real;
  wire       [17:0]   twiddle_factor_table_43_imag;
  wire       [17:0]   twiddle_factor_table_44_real;
  wire       [17:0]   twiddle_factor_table_44_imag;
  wire       [17:0]   twiddle_factor_table_45_real;
  wire       [17:0]   twiddle_factor_table_45_imag;
  wire       [17:0]   twiddle_factor_table_46_real;
  wire       [17:0]   twiddle_factor_table_46_imag;
  wire       [17:0]   twiddle_factor_table_47_real;
  wire       [17:0]   twiddle_factor_table_47_imag;
  wire       [17:0]   twiddle_factor_table_48_real;
  wire       [17:0]   twiddle_factor_table_48_imag;
  wire       [17:0]   twiddle_factor_table_49_real;
  wire       [17:0]   twiddle_factor_table_49_imag;
  wire       [17:0]   twiddle_factor_table_50_real;
  wire       [17:0]   twiddle_factor_table_50_imag;
  wire       [17:0]   twiddle_factor_table_51_real;
  wire       [17:0]   twiddle_factor_table_51_imag;
  wire       [17:0]   twiddle_factor_table_52_real;
  wire       [17:0]   twiddle_factor_table_52_imag;
  wire       [17:0]   twiddle_factor_table_53_real;
  wire       [17:0]   twiddle_factor_table_53_imag;
  wire       [17:0]   twiddle_factor_table_54_real;
  wire       [17:0]   twiddle_factor_table_54_imag;
  wire       [17:0]   twiddle_factor_table_55_real;
  wire       [17:0]   twiddle_factor_table_55_imag;
  wire       [17:0]   twiddle_factor_table_56_real;
  wire       [17:0]   twiddle_factor_table_56_imag;
  wire       [17:0]   twiddle_factor_table_57_real;
  wire       [17:0]   twiddle_factor_table_57_imag;
  wire       [17:0]   twiddle_factor_table_58_real;
  wire       [17:0]   twiddle_factor_table_58_imag;
  wire       [17:0]   twiddle_factor_table_59_real;
  wire       [17:0]   twiddle_factor_table_59_imag;
  wire       [17:0]   twiddle_factor_table_60_real;
  wire       [17:0]   twiddle_factor_table_60_imag;
  wire       [17:0]   twiddle_factor_table_61_real;
  wire       [17:0]   twiddle_factor_table_61_imag;
  wire       [17:0]   twiddle_factor_table_62_real;
  wire       [17:0]   twiddle_factor_table_62_imag;
  wire       [17:0]   data_reorder_0_real;
  wire       [17:0]   data_reorder_0_imag;
  wire       [17:0]   data_reorder_1_real;
  wire       [17:0]   data_reorder_1_imag;
  wire       [17:0]   data_reorder_2_real;
  wire       [17:0]   data_reorder_2_imag;
  wire       [17:0]   data_reorder_3_real;
  wire       [17:0]   data_reorder_3_imag;
  wire       [17:0]   data_reorder_4_real;
  wire       [17:0]   data_reorder_4_imag;
  wire       [17:0]   data_reorder_5_real;
  wire       [17:0]   data_reorder_5_imag;
  wire       [17:0]   data_reorder_6_real;
  wire       [17:0]   data_reorder_6_imag;
  wire       [17:0]   data_reorder_7_real;
  wire       [17:0]   data_reorder_7_imag;
  wire       [17:0]   data_reorder_8_real;
  wire       [17:0]   data_reorder_8_imag;
  wire       [17:0]   data_reorder_9_real;
  wire       [17:0]   data_reorder_9_imag;
  wire       [17:0]   data_reorder_10_real;
  wire       [17:0]   data_reorder_10_imag;
  wire       [17:0]   data_reorder_11_real;
  wire       [17:0]   data_reorder_11_imag;
  wire       [17:0]   data_reorder_12_real;
  wire       [17:0]   data_reorder_12_imag;
  wire       [17:0]   data_reorder_13_real;
  wire       [17:0]   data_reorder_13_imag;
  wire       [17:0]   data_reorder_14_real;
  wire       [17:0]   data_reorder_14_imag;
  wire       [17:0]   data_reorder_15_real;
  wire       [17:0]   data_reorder_15_imag;
  wire       [17:0]   data_reorder_16_real;
  wire       [17:0]   data_reorder_16_imag;
  wire       [17:0]   data_reorder_17_real;
  wire       [17:0]   data_reorder_17_imag;
  wire       [17:0]   data_reorder_18_real;
  wire       [17:0]   data_reorder_18_imag;
  wire       [17:0]   data_reorder_19_real;
  wire       [17:0]   data_reorder_19_imag;
  wire       [17:0]   data_reorder_20_real;
  wire       [17:0]   data_reorder_20_imag;
  wire       [17:0]   data_reorder_21_real;
  wire       [17:0]   data_reorder_21_imag;
  wire       [17:0]   data_reorder_22_real;
  wire       [17:0]   data_reorder_22_imag;
  wire       [17:0]   data_reorder_23_real;
  wire       [17:0]   data_reorder_23_imag;
  wire       [17:0]   data_reorder_24_real;
  wire       [17:0]   data_reorder_24_imag;
  wire       [17:0]   data_reorder_25_real;
  wire       [17:0]   data_reorder_25_imag;
  wire       [17:0]   data_reorder_26_real;
  wire       [17:0]   data_reorder_26_imag;
  wire       [17:0]   data_reorder_27_real;
  wire       [17:0]   data_reorder_27_imag;
  wire       [17:0]   data_reorder_28_real;
  wire       [17:0]   data_reorder_28_imag;
  wire       [17:0]   data_reorder_29_real;
  wire       [17:0]   data_reorder_29_imag;
  wire       [17:0]   data_reorder_30_real;
  wire       [17:0]   data_reorder_30_imag;
  wire       [17:0]   data_reorder_31_real;
  wire       [17:0]   data_reorder_31_imag;
  wire       [17:0]   data_reorder_32_real;
  wire       [17:0]   data_reorder_32_imag;
  wire       [17:0]   data_reorder_33_real;
  wire       [17:0]   data_reorder_33_imag;
  wire       [17:0]   data_reorder_34_real;
  wire       [17:0]   data_reorder_34_imag;
  wire       [17:0]   data_reorder_35_real;
  wire       [17:0]   data_reorder_35_imag;
  wire       [17:0]   data_reorder_36_real;
  wire       [17:0]   data_reorder_36_imag;
  wire       [17:0]   data_reorder_37_real;
  wire       [17:0]   data_reorder_37_imag;
  wire       [17:0]   data_reorder_38_real;
  wire       [17:0]   data_reorder_38_imag;
  wire       [17:0]   data_reorder_39_real;
  wire       [17:0]   data_reorder_39_imag;
  wire       [17:0]   data_reorder_40_real;
  wire       [17:0]   data_reorder_40_imag;
  wire       [17:0]   data_reorder_41_real;
  wire       [17:0]   data_reorder_41_imag;
  wire       [17:0]   data_reorder_42_real;
  wire       [17:0]   data_reorder_42_imag;
  wire       [17:0]   data_reorder_43_real;
  wire       [17:0]   data_reorder_43_imag;
  wire       [17:0]   data_reorder_44_real;
  wire       [17:0]   data_reorder_44_imag;
  wire       [17:0]   data_reorder_45_real;
  wire       [17:0]   data_reorder_45_imag;
  wire       [17:0]   data_reorder_46_real;
  wire       [17:0]   data_reorder_46_imag;
  wire       [17:0]   data_reorder_47_real;
  wire       [17:0]   data_reorder_47_imag;
  wire       [17:0]   data_reorder_48_real;
  wire       [17:0]   data_reorder_48_imag;
  wire       [17:0]   data_reorder_49_real;
  wire       [17:0]   data_reorder_49_imag;
  wire       [17:0]   data_reorder_50_real;
  wire       [17:0]   data_reorder_50_imag;
  wire       [17:0]   data_reorder_51_real;
  wire       [17:0]   data_reorder_51_imag;
  wire       [17:0]   data_reorder_52_real;
  wire       [17:0]   data_reorder_52_imag;
  wire       [17:0]   data_reorder_53_real;
  wire       [17:0]   data_reorder_53_imag;
  wire       [17:0]   data_reorder_54_real;
  wire       [17:0]   data_reorder_54_imag;
  wire       [17:0]   data_reorder_55_real;
  wire       [17:0]   data_reorder_55_imag;
  wire       [17:0]   data_reorder_56_real;
  wire       [17:0]   data_reorder_56_imag;
  wire       [17:0]   data_reorder_57_real;
  wire       [17:0]   data_reorder_57_imag;
  wire       [17:0]   data_reorder_58_real;
  wire       [17:0]   data_reorder_58_imag;
  wire       [17:0]   data_reorder_59_real;
  wire       [17:0]   data_reorder_59_imag;
  wire       [17:0]   data_reorder_60_real;
  wire       [17:0]   data_reorder_60_imag;
  wire       [17:0]   data_reorder_61_real;
  wire       [17:0]   data_reorder_61_imag;
  wire       [17:0]   data_reorder_62_real;
  wire       [17:0]   data_reorder_62_imag;
  wire       [17:0]   data_reorder_63_real;
  wire       [17:0]   data_reorder_63_imag;
  reg        [17:0]   data_mid_0_0_real;
  reg        [17:0]   data_mid_0_0_imag;
  reg        [17:0]   data_mid_0_1_real;
  reg        [17:0]   data_mid_0_1_imag;
  reg        [17:0]   data_mid_0_2_real;
  reg        [17:0]   data_mid_0_2_imag;
  reg        [17:0]   data_mid_0_3_real;
  reg        [17:0]   data_mid_0_3_imag;
  reg        [17:0]   data_mid_0_4_real;
  reg        [17:0]   data_mid_0_4_imag;
  reg        [17:0]   data_mid_0_5_real;
  reg        [17:0]   data_mid_0_5_imag;
  reg        [17:0]   data_mid_0_6_real;
  reg        [17:0]   data_mid_0_6_imag;
  reg        [17:0]   data_mid_0_7_real;
  reg        [17:0]   data_mid_0_7_imag;
  reg        [17:0]   data_mid_0_8_real;
  reg        [17:0]   data_mid_0_8_imag;
  reg        [17:0]   data_mid_0_9_real;
  reg        [17:0]   data_mid_0_9_imag;
  reg        [17:0]   data_mid_0_10_real;
  reg        [17:0]   data_mid_0_10_imag;
  reg        [17:0]   data_mid_0_11_real;
  reg        [17:0]   data_mid_0_11_imag;
  reg        [17:0]   data_mid_0_12_real;
  reg        [17:0]   data_mid_0_12_imag;
  reg        [17:0]   data_mid_0_13_real;
  reg        [17:0]   data_mid_0_13_imag;
  reg        [17:0]   data_mid_0_14_real;
  reg        [17:0]   data_mid_0_14_imag;
  reg        [17:0]   data_mid_0_15_real;
  reg        [17:0]   data_mid_0_15_imag;
  reg        [17:0]   data_mid_0_16_real;
  reg        [17:0]   data_mid_0_16_imag;
  reg        [17:0]   data_mid_0_17_real;
  reg        [17:0]   data_mid_0_17_imag;
  reg        [17:0]   data_mid_0_18_real;
  reg        [17:0]   data_mid_0_18_imag;
  reg        [17:0]   data_mid_0_19_real;
  reg        [17:0]   data_mid_0_19_imag;
  reg        [17:0]   data_mid_0_20_real;
  reg        [17:0]   data_mid_0_20_imag;
  reg        [17:0]   data_mid_0_21_real;
  reg        [17:0]   data_mid_0_21_imag;
  reg        [17:0]   data_mid_0_22_real;
  reg        [17:0]   data_mid_0_22_imag;
  reg        [17:0]   data_mid_0_23_real;
  reg        [17:0]   data_mid_0_23_imag;
  reg        [17:0]   data_mid_0_24_real;
  reg        [17:0]   data_mid_0_24_imag;
  reg        [17:0]   data_mid_0_25_real;
  reg        [17:0]   data_mid_0_25_imag;
  reg        [17:0]   data_mid_0_26_real;
  reg        [17:0]   data_mid_0_26_imag;
  reg        [17:0]   data_mid_0_27_real;
  reg        [17:0]   data_mid_0_27_imag;
  reg        [17:0]   data_mid_0_28_real;
  reg        [17:0]   data_mid_0_28_imag;
  reg        [17:0]   data_mid_0_29_real;
  reg        [17:0]   data_mid_0_29_imag;
  reg        [17:0]   data_mid_0_30_real;
  reg        [17:0]   data_mid_0_30_imag;
  reg        [17:0]   data_mid_0_31_real;
  reg        [17:0]   data_mid_0_31_imag;
  reg        [17:0]   data_mid_0_32_real;
  reg        [17:0]   data_mid_0_32_imag;
  reg        [17:0]   data_mid_0_33_real;
  reg        [17:0]   data_mid_0_33_imag;
  reg        [17:0]   data_mid_0_34_real;
  reg        [17:0]   data_mid_0_34_imag;
  reg        [17:0]   data_mid_0_35_real;
  reg        [17:0]   data_mid_0_35_imag;
  reg        [17:0]   data_mid_0_36_real;
  reg        [17:0]   data_mid_0_36_imag;
  reg        [17:0]   data_mid_0_37_real;
  reg        [17:0]   data_mid_0_37_imag;
  reg        [17:0]   data_mid_0_38_real;
  reg        [17:0]   data_mid_0_38_imag;
  reg        [17:0]   data_mid_0_39_real;
  reg        [17:0]   data_mid_0_39_imag;
  reg        [17:0]   data_mid_0_40_real;
  reg        [17:0]   data_mid_0_40_imag;
  reg        [17:0]   data_mid_0_41_real;
  reg        [17:0]   data_mid_0_41_imag;
  reg        [17:0]   data_mid_0_42_real;
  reg        [17:0]   data_mid_0_42_imag;
  reg        [17:0]   data_mid_0_43_real;
  reg        [17:0]   data_mid_0_43_imag;
  reg        [17:0]   data_mid_0_44_real;
  reg        [17:0]   data_mid_0_44_imag;
  reg        [17:0]   data_mid_0_45_real;
  reg        [17:0]   data_mid_0_45_imag;
  reg        [17:0]   data_mid_0_46_real;
  reg        [17:0]   data_mid_0_46_imag;
  reg        [17:0]   data_mid_0_47_real;
  reg        [17:0]   data_mid_0_47_imag;
  reg        [17:0]   data_mid_0_48_real;
  reg        [17:0]   data_mid_0_48_imag;
  reg        [17:0]   data_mid_0_49_real;
  reg        [17:0]   data_mid_0_49_imag;
  reg        [17:0]   data_mid_0_50_real;
  reg        [17:0]   data_mid_0_50_imag;
  reg        [17:0]   data_mid_0_51_real;
  reg        [17:0]   data_mid_0_51_imag;
  reg        [17:0]   data_mid_0_52_real;
  reg        [17:0]   data_mid_0_52_imag;
  reg        [17:0]   data_mid_0_53_real;
  reg        [17:0]   data_mid_0_53_imag;
  reg        [17:0]   data_mid_0_54_real;
  reg        [17:0]   data_mid_0_54_imag;
  reg        [17:0]   data_mid_0_55_real;
  reg        [17:0]   data_mid_0_55_imag;
  reg        [17:0]   data_mid_0_56_real;
  reg        [17:0]   data_mid_0_56_imag;
  reg        [17:0]   data_mid_0_57_real;
  reg        [17:0]   data_mid_0_57_imag;
  reg        [17:0]   data_mid_0_58_real;
  reg        [17:0]   data_mid_0_58_imag;
  reg        [17:0]   data_mid_0_59_real;
  reg        [17:0]   data_mid_0_59_imag;
  reg        [17:0]   data_mid_0_60_real;
  reg        [17:0]   data_mid_0_60_imag;
  reg        [17:0]   data_mid_0_61_real;
  reg        [17:0]   data_mid_0_61_imag;
  reg        [17:0]   data_mid_0_62_real;
  reg        [17:0]   data_mid_0_62_imag;
  reg        [17:0]   data_mid_0_63_real;
  reg        [17:0]   data_mid_0_63_imag;
  reg        [17:0]   data_mid_1_0_real;
  reg        [17:0]   data_mid_1_0_imag;
  reg        [17:0]   data_mid_1_1_real;
  reg        [17:0]   data_mid_1_1_imag;
  reg        [17:0]   data_mid_1_2_real;
  reg        [17:0]   data_mid_1_2_imag;
  reg        [17:0]   data_mid_1_3_real;
  reg        [17:0]   data_mid_1_3_imag;
  reg        [17:0]   data_mid_1_4_real;
  reg        [17:0]   data_mid_1_4_imag;
  reg        [17:0]   data_mid_1_5_real;
  reg        [17:0]   data_mid_1_5_imag;
  reg        [17:0]   data_mid_1_6_real;
  reg        [17:0]   data_mid_1_6_imag;
  reg        [17:0]   data_mid_1_7_real;
  reg        [17:0]   data_mid_1_7_imag;
  reg        [17:0]   data_mid_1_8_real;
  reg        [17:0]   data_mid_1_8_imag;
  reg        [17:0]   data_mid_1_9_real;
  reg        [17:0]   data_mid_1_9_imag;
  reg        [17:0]   data_mid_1_10_real;
  reg        [17:0]   data_mid_1_10_imag;
  reg        [17:0]   data_mid_1_11_real;
  reg        [17:0]   data_mid_1_11_imag;
  reg        [17:0]   data_mid_1_12_real;
  reg        [17:0]   data_mid_1_12_imag;
  reg        [17:0]   data_mid_1_13_real;
  reg        [17:0]   data_mid_1_13_imag;
  reg        [17:0]   data_mid_1_14_real;
  reg        [17:0]   data_mid_1_14_imag;
  reg        [17:0]   data_mid_1_15_real;
  reg        [17:0]   data_mid_1_15_imag;
  reg        [17:0]   data_mid_1_16_real;
  reg        [17:0]   data_mid_1_16_imag;
  reg        [17:0]   data_mid_1_17_real;
  reg        [17:0]   data_mid_1_17_imag;
  reg        [17:0]   data_mid_1_18_real;
  reg        [17:0]   data_mid_1_18_imag;
  reg        [17:0]   data_mid_1_19_real;
  reg        [17:0]   data_mid_1_19_imag;
  reg        [17:0]   data_mid_1_20_real;
  reg        [17:0]   data_mid_1_20_imag;
  reg        [17:0]   data_mid_1_21_real;
  reg        [17:0]   data_mid_1_21_imag;
  reg        [17:0]   data_mid_1_22_real;
  reg        [17:0]   data_mid_1_22_imag;
  reg        [17:0]   data_mid_1_23_real;
  reg        [17:0]   data_mid_1_23_imag;
  reg        [17:0]   data_mid_1_24_real;
  reg        [17:0]   data_mid_1_24_imag;
  reg        [17:0]   data_mid_1_25_real;
  reg        [17:0]   data_mid_1_25_imag;
  reg        [17:0]   data_mid_1_26_real;
  reg        [17:0]   data_mid_1_26_imag;
  reg        [17:0]   data_mid_1_27_real;
  reg        [17:0]   data_mid_1_27_imag;
  reg        [17:0]   data_mid_1_28_real;
  reg        [17:0]   data_mid_1_28_imag;
  reg        [17:0]   data_mid_1_29_real;
  reg        [17:0]   data_mid_1_29_imag;
  reg        [17:0]   data_mid_1_30_real;
  reg        [17:0]   data_mid_1_30_imag;
  reg        [17:0]   data_mid_1_31_real;
  reg        [17:0]   data_mid_1_31_imag;
  reg        [17:0]   data_mid_1_32_real;
  reg        [17:0]   data_mid_1_32_imag;
  reg        [17:0]   data_mid_1_33_real;
  reg        [17:0]   data_mid_1_33_imag;
  reg        [17:0]   data_mid_1_34_real;
  reg        [17:0]   data_mid_1_34_imag;
  reg        [17:0]   data_mid_1_35_real;
  reg        [17:0]   data_mid_1_35_imag;
  reg        [17:0]   data_mid_1_36_real;
  reg        [17:0]   data_mid_1_36_imag;
  reg        [17:0]   data_mid_1_37_real;
  reg        [17:0]   data_mid_1_37_imag;
  reg        [17:0]   data_mid_1_38_real;
  reg        [17:0]   data_mid_1_38_imag;
  reg        [17:0]   data_mid_1_39_real;
  reg        [17:0]   data_mid_1_39_imag;
  reg        [17:0]   data_mid_1_40_real;
  reg        [17:0]   data_mid_1_40_imag;
  reg        [17:0]   data_mid_1_41_real;
  reg        [17:0]   data_mid_1_41_imag;
  reg        [17:0]   data_mid_1_42_real;
  reg        [17:0]   data_mid_1_42_imag;
  reg        [17:0]   data_mid_1_43_real;
  reg        [17:0]   data_mid_1_43_imag;
  reg        [17:0]   data_mid_1_44_real;
  reg        [17:0]   data_mid_1_44_imag;
  reg        [17:0]   data_mid_1_45_real;
  reg        [17:0]   data_mid_1_45_imag;
  reg        [17:0]   data_mid_1_46_real;
  reg        [17:0]   data_mid_1_46_imag;
  reg        [17:0]   data_mid_1_47_real;
  reg        [17:0]   data_mid_1_47_imag;
  reg        [17:0]   data_mid_1_48_real;
  reg        [17:0]   data_mid_1_48_imag;
  reg        [17:0]   data_mid_1_49_real;
  reg        [17:0]   data_mid_1_49_imag;
  reg        [17:0]   data_mid_1_50_real;
  reg        [17:0]   data_mid_1_50_imag;
  reg        [17:0]   data_mid_1_51_real;
  reg        [17:0]   data_mid_1_51_imag;
  reg        [17:0]   data_mid_1_52_real;
  reg        [17:0]   data_mid_1_52_imag;
  reg        [17:0]   data_mid_1_53_real;
  reg        [17:0]   data_mid_1_53_imag;
  reg        [17:0]   data_mid_1_54_real;
  reg        [17:0]   data_mid_1_54_imag;
  reg        [17:0]   data_mid_1_55_real;
  reg        [17:0]   data_mid_1_55_imag;
  reg        [17:0]   data_mid_1_56_real;
  reg        [17:0]   data_mid_1_56_imag;
  reg        [17:0]   data_mid_1_57_real;
  reg        [17:0]   data_mid_1_57_imag;
  reg        [17:0]   data_mid_1_58_real;
  reg        [17:0]   data_mid_1_58_imag;
  reg        [17:0]   data_mid_1_59_real;
  reg        [17:0]   data_mid_1_59_imag;
  reg        [17:0]   data_mid_1_60_real;
  reg        [17:0]   data_mid_1_60_imag;
  reg        [17:0]   data_mid_1_61_real;
  reg        [17:0]   data_mid_1_61_imag;
  reg        [17:0]   data_mid_1_62_real;
  reg        [17:0]   data_mid_1_62_imag;
  reg        [17:0]   data_mid_1_63_real;
  reg        [17:0]   data_mid_1_63_imag;
  reg        [17:0]   data_mid_2_0_real;
  reg        [17:0]   data_mid_2_0_imag;
  reg        [17:0]   data_mid_2_1_real;
  reg        [17:0]   data_mid_2_1_imag;
  reg        [17:0]   data_mid_2_2_real;
  reg        [17:0]   data_mid_2_2_imag;
  reg        [17:0]   data_mid_2_3_real;
  reg        [17:0]   data_mid_2_3_imag;
  reg        [17:0]   data_mid_2_4_real;
  reg        [17:0]   data_mid_2_4_imag;
  reg        [17:0]   data_mid_2_5_real;
  reg        [17:0]   data_mid_2_5_imag;
  reg        [17:0]   data_mid_2_6_real;
  reg        [17:0]   data_mid_2_6_imag;
  reg        [17:0]   data_mid_2_7_real;
  reg        [17:0]   data_mid_2_7_imag;
  reg        [17:0]   data_mid_2_8_real;
  reg        [17:0]   data_mid_2_8_imag;
  reg        [17:0]   data_mid_2_9_real;
  reg        [17:0]   data_mid_2_9_imag;
  reg        [17:0]   data_mid_2_10_real;
  reg        [17:0]   data_mid_2_10_imag;
  reg        [17:0]   data_mid_2_11_real;
  reg        [17:0]   data_mid_2_11_imag;
  reg        [17:0]   data_mid_2_12_real;
  reg        [17:0]   data_mid_2_12_imag;
  reg        [17:0]   data_mid_2_13_real;
  reg        [17:0]   data_mid_2_13_imag;
  reg        [17:0]   data_mid_2_14_real;
  reg        [17:0]   data_mid_2_14_imag;
  reg        [17:0]   data_mid_2_15_real;
  reg        [17:0]   data_mid_2_15_imag;
  reg        [17:0]   data_mid_2_16_real;
  reg        [17:0]   data_mid_2_16_imag;
  reg        [17:0]   data_mid_2_17_real;
  reg        [17:0]   data_mid_2_17_imag;
  reg        [17:0]   data_mid_2_18_real;
  reg        [17:0]   data_mid_2_18_imag;
  reg        [17:0]   data_mid_2_19_real;
  reg        [17:0]   data_mid_2_19_imag;
  reg        [17:0]   data_mid_2_20_real;
  reg        [17:0]   data_mid_2_20_imag;
  reg        [17:0]   data_mid_2_21_real;
  reg        [17:0]   data_mid_2_21_imag;
  reg        [17:0]   data_mid_2_22_real;
  reg        [17:0]   data_mid_2_22_imag;
  reg        [17:0]   data_mid_2_23_real;
  reg        [17:0]   data_mid_2_23_imag;
  reg        [17:0]   data_mid_2_24_real;
  reg        [17:0]   data_mid_2_24_imag;
  reg        [17:0]   data_mid_2_25_real;
  reg        [17:0]   data_mid_2_25_imag;
  reg        [17:0]   data_mid_2_26_real;
  reg        [17:0]   data_mid_2_26_imag;
  reg        [17:0]   data_mid_2_27_real;
  reg        [17:0]   data_mid_2_27_imag;
  reg        [17:0]   data_mid_2_28_real;
  reg        [17:0]   data_mid_2_28_imag;
  reg        [17:0]   data_mid_2_29_real;
  reg        [17:0]   data_mid_2_29_imag;
  reg        [17:0]   data_mid_2_30_real;
  reg        [17:0]   data_mid_2_30_imag;
  reg        [17:0]   data_mid_2_31_real;
  reg        [17:0]   data_mid_2_31_imag;
  reg        [17:0]   data_mid_2_32_real;
  reg        [17:0]   data_mid_2_32_imag;
  reg        [17:0]   data_mid_2_33_real;
  reg        [17:0]   data_mid_2_33_imag;
  reg        [17:0]   data_mid_2_34_real;
  reg        [17:0]   data_mid_2_34_imag;
  reg        [17:0]   data_mid_2_35_real;
  reg        [17:0]   data_mid_2_35_imag;
  reg        [17:0]   data_mid_2_36_real;
  reg        [17:0]   data_mid_2_36_imag;
  reg        [17:0]   data_mid_2_37_real;
  reg        [17:0]   data_mid_2_37_imag;
  reg        [17:0]   data_mid_2_38_real;
  reg        [17:0]   data_mid_2_38_imag;
  reg        [17:0]   data_mid_2_39_real;
  reg        [17:0]   data_mid_2_39_imag;
  reg        [17:0]   data_mid_2_40_real;
  reg        [17:0]   data_mid_2_40_imag;
  reg        [17:0]   data_mid_2_41_real;
  reg        [17:0]   data_mid_2_41_imag;
  reg        [17:0]   data_mid_2_42_real;
  reg        [17:0]   data_mid_2_42_imag;
  reg        [17:0]   data_mid_2_43_real;
  reg        [17:0]   data_mid_2_43_imag;
  reg        [17:0]   data_mid_2_44_real;
  reg        [17:0]   data_mid_2_44_imag;
  reg        [17:0]   data_mid_2_45_real;
  reg        [17:0]   data_mid_2_45_imag;
  reg        [17:0]   data_mid_2_46_real;
  reg        [17:0]   data_mid_2_46_imag;
  reg        [17:0]   data_mid_2_47_real;
  reg        [17:0]   data_mid_2_47_imag;
  reg        [17:0]   data_mid_2_48_real;
  reg        [17:0]   data_mid_2_48_imag;
  reg        [17:0]   data_mid_2_49_real;
  reg        [17:0]   data_mid_2_49_imag;
  reg        [17:0]   data_mid_2_50_real;
  reg        [17:0]   data_mid_2_50_imag;
  reg        [17:0]   data_mid_2_51_real;
  reg        [17:0]   data_mid_2_51_imag;
  reg        [17:0]   data_mid_2_52_real;
  reg        [17:0]   data_mid_2_52_imag;
  reg        [17:0]   data_mid_2_53_real;
  reg        [17:0]   data_mid_2_53_imag;
  reg        [17:0]   data_mid_2_54_real;
  reg        [17:0]   data_mid_2_54_imag;
  reg        [17:0]   data_mid_2_55_real;
  reg        [17:0]   data_mid_2_55_imag;
  reg        [17:0]   data_mid_2_56_real;
  reg        [17:0]   data_mid_2_56_imag;
  reg        [17:0]   data_mid_2_57_real;
  reg        [17:0]   data_mid_2_57_imag;
  reg        [17:0]   data_mid_2_58_real;
  reg        [17:0]   data_mid_2_58_imag;
  reg        [17:0]   data_mid_2_59_real;
  reg        [17:0]   data_mid_2_59_imag;
  reg        [17:0]   data_mid_2_60_real;
  reg        [17:0]   data_mid_2_60_imag;
  reg        [17:0]   data_mid_2_61_real;
  reg        [17:0]   data_mid_2_61_imag;
  reg        [17:0]   data_mid_2_62_real;
  reg        [17:0]   data_mid_2_62_imag;
  reg        [17:0]   data_mid_2_63_real;
  reg        [17:0]   data_mid_2_63_imag;
  reg        [17:0]   data_mid_3_0_real;
  reg        [17:0]   data_mid_3_0_imag;
  reg        [17:0]   data_mid_3_1_real;
  reg        [17:0]   data_mid_3_1_imag;
  reg        [17:0]   data_mid_3_2_real;
  reg        [17:0]   data_mid_3_2_imag;
  reg        [17:0]   data_mid_3_3_real;
  reg        [17:0]   data_mid_3_3_imag;
  reg        [17:0]   data_mid_3_4_real;
  reg        [17:0]   data_mid_3_4_imag;
  reg        [17:0]   data_mid_3_5_real;
  reg        [17:0]   data_mid_3_5_imag;
  reg        [17:0]   data_mid_3_6_real;
  reg        [17:0]   data_mid_3_6_imag;
  reg        [17:0]   data_mid_3_7_real;
  reg        [17:0]   data_mid_3_7_imag;
  reg        [17:0]   data_mid_3_8_real;
  reg        [17:0]   data_mid_3_8_imag;
  reg        [17:0]   data_mid_3_9_real;
  reg        [17:0]   data_mid_3_9_imag;
  reg        [17:0]   data_mid_3_10_real;
  reg        [17:0]   data_mid_3_10_imag;
  reg        [17:0]   data_mid_3_11_real;
  reg        [17:0]   data_mid_3_11_imag;
  reg        [17:0]   data_mid_3_12_real;
  reg        [17:0]   data_mid_3_12_imag;
  reg        [17:0]   data_mid_3_13_real;
  reg        [17:0]   data_mid_3_13_imag;
  reg        [17:0]   data_mid_3_14_real;
  reg        [17:0]   data_mid_3_14_imag;
  reg        [17:0]   data_mid_3_15_real;
  reg        [17:0]   data_mid_3_15_imag;
  reg        [17:0]   data_mid_3_16_real;
  reg        [17:0]   data_mid_3_16_imag;
  reg        [17:0]   data_mid_3_17_real;
  reg        [17:0]   data_mid_3_17_imag;
  reg        [17:0]   data_mid_3_18_real;
  reg        [17:0]   data_mid_3_18_imag;
  reg        [17:0]   data_mid_3_19_real;
  reg        [17:0]   data_mid_3_19_imag;
  reg        [17:0]   data_mid_3_20_real;
  reg        [17:0]   data_mid_3_20_imag;
  reg        [17:0]   data_mid_3_21_real;
  reg        [17:0]   data_mid_3_21_imag;
  reg        [17:0]   data_mid_3_22_real;
  reg        [17:0]   data_mid_3_22_imag;
  reg        [17:0]   data_mid_3_23_real;
  reg        [17:0]   data_mid_3_23_imag;
  reg        [17:0]   data_mid_3_24_real;
  reg        [17:0]   data_mid_3_24_imag;
  reg        [17:0]   data_mid_3_25_real;
  reg        [17:0]   data_mid_3_25_imag;
  reg        [17:0]   data_mid_3_26_real;
  reg        [17:0]   data_mid_3_26_imag;
  reg        [17:0]   data_mid_3_27_real;
  reg        [17:0]   data_mid_3_27_imag;
  reg        [17:0]   data_mid_3_28_real;
  reg        [17:0]   data_mid_3_28_imag;
  reg        [17:0]   data_mid_3_29_real;
  reg        [17:0]   data_mid_3_29_imag;
  reg        [17:0]   data_mid_3_30_real;
  reg        [17:0]   data_mid_3_30_imag;
  reg        [17:0]   data_mid_3_31_real;
  reg        [17:0]   data_mid_3_31_imag;
  reg        [17:0]   data_mid_3_32_real;
  reg        [17:0]   data_mid_3_32_imag;
  reg        [17:0]   data_mid_3_33_real;
  reg        [17:0]   data_mid_3_33_imag;
  reg        [17:0]   data_mid_3_34_real;
  reg        [17:0]   data_mid_3_34_imag;
  reg        [17:0]   data_mid_3_35_real;
  reg        [17:0]   data_mid_3_35_imag;
  reg        [17:0]   data_mid_3_36_real;
  reg        [17:0]   data_mid_3_36_imag;
  reg        [17:0]   data_mid_3_37_real;
  reg        [17:0]   data_mid_3_37_imag;
  reg        [17:0]   data_mid_3_38_real;
  reg        [17:0]   data_mid_3_38_imag;
  reg        [17:0]   data_mid_3_39_real;
  reg        [17:0]   data_mid_3_39_imag;
  reg        [17:0]   data_mid_3_40_real;
  reg        [17:0]   data_mid_3_40_imag;
  reg        [17:0]   data_mid_3_41_real;
  reg        [17:0]   data_mid_3_41_imag;
  reg        [17:0]   data_mid_3_42_real;
  reg        [17:0]   data_mid_3_42_imag;
  reg        [17:0]   data_mid_3_43_real;
  reg        [17:0]   data_mid_3_43_imag;
  reg        [17:0]   data_mid_3_44_real;
  reg        [17:0]   data_mid_3_44_imag;
  reg        [17:0]   data_mid_3_45_real;
  reg        [17:0]   data_mid_3_45_imag;
  reg        [17:0]   data_mid_3_46_real;
  reg        [17:0]   data_mid_3_46_imag;
  reg        [17:0]   data_mid_3_47_real;
  reg        [17:0]   data_mid_3_47_imag;
  reg        [17:0]   data_mid_3_48_real;
  reg        [17:0]   data_mid_3_48_imag;
  reg        [17:0]   data_mid_3_49_real;
  reg        [17:0]   data_mid_3_49_imag;
  reg        [17:0]   data_mid_3_50_real;
  reg        [17:0]   data_mid_3_50_imag;
  reg        [17:0]   data_mid_3_51_real;
  reg        [17:0]   data_mid_3_51_imag;
  reg        [17:0]   data_mid_3_52_real;
  reg        [17:0]   data_mid_3_52_imag;
  reg        [17:0]   data_mid_3_53_real;
  reg        [17:0]   data_mid_3_53_imag;
  reg        [17:0]   data_mid_3_54_real;
  reg        [17:0]   data_mid_3_54_imag;
  reg        [17:0]   data_mid_3_55_real;
  reg        [17:0]   data_mid_3_55_imag;
  reg        [17:0]   data_mid_3_56_real;
  reg        [17:0]   data_mid_3_56_imag;
  reg        [17:0]   data_mid_3_57_real;
  reg        [17:0]   data_mid_3_57_imag;
  reg        [17:0]   data_mid_3_58_real;
  reg        [17:0]   data_mid_3_58_imag;
  reg        [17:0]   data_mid_3_59_real;
  reg        [17:0]   data_mid_3_59_imag;
  reg        [17:0]   data_mid_3_60_real;
  reg        [17:0]   data_mid_3_60_imag;
  reg        [17:0]   data_mid_3_61_real;
  reg        [17:0]   data_mid_3_61_imag;
  reg        [17:0]   data_mid_3_62_real;
  reg        [17:0]   data_mid_3_62_imag;
  reg        [17:0]   data_mid_3_63_real;
  reg        [17:0]   data_mid_3_63_imag;
  reg        [17:0]   data_mid_4_0_real;
  reg        [17:0]   data_mid_4_0_imag;
  reg        [17:0]   data_mid_4_1_real;
  reg        [17:0]   data_mid_4_1_imag;
  reg        [17:0]   data_mid_4_2_real;
  reg        [17:0]   data_mid_4_2_imag;
  reg        [17:0]   data_mid_4_3_real;
  reg        [17:0]   data_mid_4_3_imag;
  reg        [17:0]   data_mid_4_4_real;
  reg        [17:0]   data_mid_4_4_imag;
  reg        [17:0]   data_mid_4_5_real;
  reg        [17:0]   data_mid_4_5_imag;
  reg        [17:0]   data_mid_4_6_real;
  reg        [17:0]   data_mid_4_6_imag;
  reg        [17:0]   data_mid_4_7_real;
  reg        [17:0]   data_mid_4_7_imag;
  reg        [17:0]   data_mid_4_8_real;
  reg        [17:0]   data_mid_4_8_imag;
  reg        [17:0]   data_mid_4_9_real;
  reg        [17:0]   data_mid_4_9_imag;
  reg        [17:0]   data_mid_4_10_real;
  reg        [17:0]   data_mid_4_10_imag;
  reg        [17:0]   data_mid_4_11_real;
  reg        [17:0]   data_mid_4_11_imag;
  reg        [17:0]   data_mid_4_12_real;
  reg        [17:0]   data_mid_4_12_imag;
  reg        [17:0]   data_mid_4_13_real;
  reg        [17:0]   data_mid_4_13_imag;
  reg        [17:0]   data_mid_4_14_real;
  reg        [17:0]   data_mid_4_14_imag;
  reg        [17:0]   data_mid_4_15_real;
  reg        [17:0]   data_mid_4_15_imag;
  reg        [17:0]   data_mid_4_16_real;
  reg        [17:0]   data_mid_4_16_imag;
  reg        [17:0]   data_mid_4_17_real;
  reg        [17:0]   data_mid_4_17_imag;
  reg        [17:0]   data_mid_4_18_real;
  reg        [17:0]   data_mid_4_18_imag;
  reg        [17:0]   data_mid_4_19_real;
  reg        [17:0]   data_mid_4_19_imag;
  reg        [17:0]   data_mid_4_20_real;
  reg        [17:0]   data_mid_4_20_imag;
  reg        [17:0]   data_mid_4_21_real;
  reg        [17:0]   data_mid_4_21_imag;
  reg        [17:0]   data_mid_4_22_real;
  reg        [17:0]   data_mid_4_22_imag;
  reg        [17:0]   data_mid_4_23_real;
  reg        [17:0]   data_mid_4_23_imag;
  reg        [17:0]   data_mid_4_24_real;
  reg        [17:0]   data_mid_4_24_imag;
  reg        [17:0]   data_mid_4_25_real;
  reg        [17:0]   data_mid_4_25_imag;
  reg        [17:0]   data_mid_4_26_real;
  reg        [17:0]   data_mid_4_26_imag;
  reg        [17:0]   data_mid_4_27_real;
  reg        [17:0]   data_mid_4_27_imag;
  reg        [17:0]   data_mid_4_28_real;
  reg        [17:0]   data_mid_4_28_imag;
  reg        [17:0]   data_mid_4_29_real;
  reg        [17:0]   data_mid_4_29_imag;
  reg        [17:0]   data_mid_4_30_real;
  reg        [17:0]   data_mid_4_30_imag;
  reg        [17:0]   data_mid_4_31_real;
  reg        [17:0]   data_mid_4_31_imag;
  reg        [17:0]   data_mid_4_32_real;
  reg        [17:0]   data_mid_4_32_imag;
  reg        [17:0]   data_mid_4_33_real;
  reg        [17:0]   data_mid_4_33_imag;
  reg        [17:0]   data_mid_4_34_real;
  reg        [17:0]   data_mid_4_34_imag;
  reg        [17:0]   data_mid_4_35_real;
  reg        [17:0]   data_mid_4_35_imag;
  reg        [17:0]   data_mid_4_36_real;
  reg        [17:0]   data_mid_4_36_imag;
  reg        [17:0]   data_mid_4_37_real;
  reg        [17:0]   data_mid_4_37_imag;
  reg        [17:0]   data_mid_4_38_real;
  reg        [17:0]   data_mid_4_38_imag;
  reg        [17:0]   data_mid_4_39_real;
  reg        [17:0]   data_mid_4_39_imag;
  reg        [17:0]   data_mid_4_40_real;
  reg        [17:0]   data_mid_4_40_imag;
  reg        [17:0]   data_mid_4_41_real;
  reg        [17:0]   data_mid_4_41_imag;
  reg        [17:0]   data_mid_4_42_real;
  reg        [17:0]   data_mid_4_42_imag;
  reg        [17:0]   data_mid_4_43_real;
  reg        [17:0]   data_mid_4_43_imag;
  reg        [17:0]   data_mid_4_44_real;
  reg        [17:0]   data_mid_4_44_imag;
  reg        [17:0]   data_mid_4_45_real;
  reg        [17:0]   data_mid_4_45_imag;
  reg        [17:0]   data_mid_4_46_real;
  reg        [17:0]   data_mid_4_46_imag;
  reg        [17:0]   data_mid_4_47_real;
  reg        [17:0]   data_mid_4_47_imag;
  reg        [17:0]   data_mid_4_48_real;
  reg        [17:0]   data_mid_4_48_imag;
  reg        [17:0]   data_mid_4_49_real;
  reg        [17:0]   data_mid_4_49_imag;
  reg        [17:0]   data_mid_4_50_real;
  reg        [17:0]   data_mid_4_50_imag;
  reg        [17:0]   data_mid_4_51_real;
  reg        [17:0]   data_mid_4_51_imag;
  reg        [17:0]   data_mid_4_52_real;
  reg        [17:0]   data_mid_4_52_imag;
  reg        [17:0]   data_mid_4_53_real;
  reg        [17:0]   data_mid_4_53_imag;
  reg        [17:0]   data_mid_4_54_real;
  reg        [17:0]   data_mid_4_54_imag;
  reg        [17:0]   data_mid_4_55_real;
  reg        [17:0]   data_mid_4_55_imag;
  reg        [17:0]   data_mid_4_56_real;
  reg        [17:0]   data_mid_4_56_imag;
  reg        [17:0]   data_mid_4_57_real;
  reg        [17:0]   data_mid_4_57_imag;
  reg        [17:0]   data_mid_4_58_real;
  reg        [17:0]   data_mid_4_58_imag;
  reg        [17:0]   data_mid_4_59_real;
  reg        [17:0]   data_mid_4_59_imag;
  reg        [17:0]   data_mid_4_60_real;
  reg        [17:0]   data_mid_4_60_imag;
  reg        [17:0]   data_mid_4_61_real;
  reg        [17:0]   data_mid_4_61_imag;
  reg        [17:0]   data_mid_4_62_real;
  reg        [17:0]   data_mid_4_62_imag;
  reg        [17:0]   data_mid_4_63_real;
  reg        [17:0]   data_mid_4_63_imag;
  reg        [17:0]   data_mid_5_0_real;
  reg        [17:0]   data_mid_5_0_imag;
  reg        [17:0]   data_mid_5_1_real;
  reg        [17:0]   data_mid_5_1_imag;
  reg        [17:0]   data_mid_5_2_real;
  reg        [17:0]   data_mid_5_2_imag;
  reg        [17:0]   data_mid_5_3_real;
  reg        [17:0]   data_mid_5_3_imag;
  reg        [17:0]   data_mid_5_4_real;
  reg        [17:0]   data_mid_5_4_imag;
  reg        [17:0]   data_mid_5_5_real;
  reg        [17:0]   data_mid_5_5_imag;
  reg        [17:0]   data_mid_5_6_real;
  reg        [17:0]   data_mid_5_6_imag;
  reg        [17:0]   data_mid_5_7_real;
  reg        [17:0]   data_mid_5_7_imag;
  reg        [17:0]   data_mid_5_8_real;
  reg        [17:0]   data_mid_5_8_imag;
  reg        [17:0]   data_mid_5_9_real;
  reg        [17:0]   data_mid_5_9_imag;
  reg        [17:0]   data_mid_5_10_real;
  reg        [17:0]   data_mid_5_10_imag;
  reg        [17:0]   data_mid_5_11_real;
  reg        [17:0]   data_mid_5_11_imag;
  reg        [17:0]   data_mid_5_12_real;
  reg        [17:0]   data_mid_5_12_imag;
  reg        [17:0]   data_mid_5_13_real;
  reg        [17:0]   data_mid_5_13_imag;
  reg        [17:0]   data_mid_5_14_real;
  reg        [17:0]   data_mid_5_14_imag;
  reg        [17:0]   data_mid_5_15_real;
  reg        [17:0]   data_mid_5_15_imag;
  reg        [17:0]   data_mid_5_16_real;
  reg        [17:0]   data_mid_5_16_imag;
  reg        [17:0]   data_mid_5_17_real;
  reg        [17:0]   data_mid_5_17_imag;
  reg        [17:0]   data_mid_5_18_real;
  reg        [17:0]   data_mid_5_18_imag;
  reg        [17:0]   data_mid_5_19_real;
  reg        [17:0]   data_mid_5_19_imag;
  reg        [17:0]   data_mid_5_20_real;
  reg        [17:0]   data_mid_5_20_imag;
  reg        [17:0]   data_mid_5_21_real;
  reg        [17:0]   data_mid_5_21_imag;
  reg        [17:0]   data_mid_5_22_real;
  reg        [17:0]   data_mid_5_22_imag;
  reg        [17:0]   data_mid_5_23_real;
  reg        [17:0]   data_mid_5_23_imag;
  reg        [17:0]   data_mid_5_24_real;
  reg        [17:0]   data_mid_5_24_imag;
  reg        [17:0]   data_mid_5_25_real;
  reg        [17:0]   data_mid_5_25_imag;
  reg        [17:0]   data_mid_5_26_real;
  reg        [17:0]   data_mid_5_26_imag;
  reg        [17:0]   data_mid_5_27_real;
  reg        [17:0]   data_mid_5_27_imag;
  reg        [17:0]   data_mid_5_28_real;
  reg        [17:0]   data_mid_5_28_imag;
  reg        [17:0]   data_mid_5_29_real;
  reg        [17:0]   data_mid_5_29_imag;
  reg        [17:0]   data_mid_5_30_real;
  reg        [17:0]   data_mid_5_30_imag;
  reg        [17:0]   data_mid_5_31_real;
  reg        [17:0]   data_mid_5_31_imag;
  reg        [17:0]   data_mid_5_32_real;
  reg        [17:0]   data_mid_5_32_imag;
  reg        [17:0]   data_mid_5_33_real;
  reg        [17:0]   data_mid_5_33_imag;
  reg        [17:0]   data_mid_5_34_real;
  reg        [17:0]   data_mid_5_34_imag;
  reg        [17:0]   data_mid_5_35_real;
  reg        [17:0]   data_mid_5_35_imag;
  reg        [17:0]   data_mid_5_36_real;
  reg        [17:0]   data_mid_5_36_imag;
  reg        [17:0]   data_mid_5_37_real;
  reg        [17:0]   data_mid_5_37_imag;
  reg        [17:0]   data_mid_5_38_real;
  reg        [17:0]   data_mid_5_38_imag;
  reg        [17:0]   data_mid_5_39_real;
  reg        [17:0]   data_mid_5_39_imag;
  reg        [17:0]   data_mid_5_40_real;
  reg        [17:0]   data_mid_5_40_imag;
  reg        [17:0]   data_mid_5_41_real;
  reg        [17:0]   data_mid_5_41_imag;
  reg        [17:0]   data_mid_5_42_real;
  reg        [17:0]   data_mid_5_42_imag;
  reg        [17:0]   data_mid_5_43_real;
  reg        [17:0]   data_mid_5_43_imag;
  reg        [17:0]   data_mid_5_44_real;
  reg        [17:0]   data_mid_5_44_imag;
  reg        [17:0]   data_mid_5_45_real;
  reg        [17:0]   data_mid_5_45_imag;
  reg        [17:0]   data_mid_5_46_real;
  reg        [17:0]   data_mid_5_46_imag;
  reg        [17:0]   data_mid_5_47_real;
  reg        [17:0]   data_mid_5_47_imag;
  reg        [17:0]   data_mid_5_48_real;
  reg        [17:0]   data_mid_5_48_imag;
  reg        [17:0]   data_mid_5_49_real;
  reg        [17:0]   data_mid_5_49_imag;
  reg        [17:0]   data_mid_5_50_real;
  reg        [17:0]   data_mid_5_50_imag;
  reg        [17:0]   data_mid_5_51_real;
  reg        [17:0]   data_mid_5_51_imag;
  reg        [17:0]   data_mid_5_52_real;
  reg        [17:0]   data_mid_5_52_imag;
  reg        [17:0]   data_mid_5_53_real;
  reg        [17:0]   data_mid_5_53_imag;
  reg        [17:0]   data_mid_5_54_real;
  reg        [17:0]   data_mid_5_54_imag;
  reg        [17:0]   data_mid_5_55_real;
  reg        [17:0]   data_mid_5_55_imag;
  reg        [17:0]   data_mid_5_56_real;
  reg        [17:0]   data_mid_5_56_imag;
  reg        [17:0]   data_mid_5_57_real;
  reg        [17:0]   data_mid_5_57_imag;
  reg        [17:0]   data_mid_5_58_real;
  reg        [17:0]   data_mid_5_58_imag;
  reg        [17:0]   data_mid_5_59_real;
  reg        [17:0]   data_mid_5_59_imag;
  reg        [17:0]   data_mid_5_60_real;
  reg        [17:0]   data_mid_5_60_imag;
  reg        [17:0]   data_mid_5_61_real;
  reg        [17:0]   data_mid_5_61_imag;
  reg        [17:0]   data_mid_5_62_real;
  reg        [17:0]   data_mid_5_62_imag;
  reg        [17:0]   data_mid_5_63_real;
  reg        [17:0]   data_mid_5_63_imag;
  reg        [17:0]   data_mid_6_0_real;
  reg        [17:0]   data_mid_6_0_imag;
  reg        [17:0]   data_mid_6_1_real;
  reg        [17:0]   data_mid_6_1_imag;
  reg        [17:0]   data_mid_6_2_real;
  reg        [17:0]   data_mid_6_2_imag;
  reg        [17:0]   data_mid_6_3_real;
  reg        [17:0]   data_mid_6_3_imag;
  reg        [17:0]   data_mid_6_4_real;
  reg        [17:0]   data_mid_6_4_imag;
  reg        [17:0]   data_mid_6_5_real;
  reg        [17:0]   data_mid_6_5_imag;
  reg        [17:0]   data_mid_6_6_real;
  reg        [17:0]   data_mid_6_6_imag;
  reg        [17:0]   data_mid_6_7_real;
  reg        [17:0]   data_mid_6_7_imag;
  reg        [17:0]   data_mid_6_8_real;
  reg        [17:0]   data_mid_6_8_imag;
  reg        [17:0]   data_mid_6_9_real;
  reg        [17:0]   data_mid_6_9_imag;
  reg        [17:0]   data_mid_6_10_real;
  reg        [17:0]   data_mid_6_10_imag;
  reg        [17:0]   data_mid_6_11_real;
  reg        [17:0]   data_mid_6_11_imag;
  reg        [17:0]   data_mid_6_12_real;
  reg        [17:0]   data_mid_6_12_imag;
  reg        [17:0]   data_mid_6_13_real;
  reg        [17:0]   data_mid_6_13_imag;
  reg        [17:0]   data_mid_6_14_real;
  reg        [17:0]   data_mid_6_14_imag;
  reg        [17:0]   data_mid_6_15_real;
  reg        [17:0]   data_mid_6_15_imag;
  reg        [17:0]   data_mid_6_16_real;
  reg        [17:0]   data_mid_6_16_imag;
  reg        [17:0]   data_mid_6_17_real;
  reg        [17:0]   data_mid_6_17_imag;
  reg        [17:0]   data_mid_6_18_real;
  reg        [17:0]   data_mid_6_18_imag;
  reg        [17:0]   data_mid_6_19_real;
  reg        [17:0]   data_mid_6_19_imag;
  reg        [17:0]   data_mid_6_20_real;
  reg        [17:0]   data_mid_6_20_imag;
  reg        [17:0]   data_mid_6_21_real;
  reg        [17:0]   data_mid_6_21_imag;
  reg        [17:0]   data_mid_6_22_real;
  reg        [17:0]   data_mid_6_22_imag;
  reg        [17:0]   data_mid_6_23_real;
  reg        [17:0]   data_mid_6_23_imag;
  reg        [17:0]   data_mid_6_24_real;
  reg        [17:0]   data_mid_6_24_imag;
  reg        [17:0]   data_mid_6_25_real;
  reg        [17:0]   data_mid_6_25_imag;
  reg        [17:0]   data_mid_6_26_real;
  reg        [17:0]   data_mid_6_26_imag;
  reg        [17:0]   data_mid_6_27_real;
  reg        [17:0]   data_mid_6_27_imag;
  reg        [17:0]   data_mid_6_28_real;
  reg        [17:0]   data_mid_6_28_imag;
  reg        [17:0]   data_mid_6_29_real;
  reg        [17:0]   data_mid_6_29_imag;
  reg        [17:0]   data_mid_6_30_real;
  reg        [17:0]   data_mid_6_30_imag;
  reg        [17:0]   data_mid_6_31_real;
  reg        [17:0]   data_mid_6_31_imag;
  reg        [17:0]   data_mid_6_32_real;
  reg        [17:0]   data_mid_6_32_imag;
  reg        [17:0]   data_mid_6_33_real;
  reg        [17:0]   data_mid_6_33_imag;
  reg        [17:0]   data_mid_6_34_real;
  reg        [17:0]   data_mid_6_34_imag;
  reg        [17:0]   data_mid_6_35_real;
  reg        [17:0]   data_mid_6_35_imag;
  reg        [17:0]   data_mid_6_36_real;
  reg        [17:0]   data_mid_6_36_imag;
  reg        [17:0]   data_mid_6_37_real;
  reg        [17:0]   data_mid_6_37_imag;
  reg        [17:0]   data_mid_6_38_real;
  reg        [17:0]   data_mid_6_38_imag;
  reg        [17:0]   data_mid_6_39_real;
  reg        [17:0]   data_mid_6_39_imag;
  reg        [17:0]   data_mid_6_40_real;
  reg        [17:0]   data_mid_6_40_imag;
  reg        [17:0]   data_mid_6_41_real;
  reg        [17:0]   data_mid_6_41_imag;
  reg        [17:0]   data_mid_6_42_real;
  reg        [17:0]   data_mid_6_42_imag;
  reg        [17:0]   data_mid_6_43_real;
  reg        [17:0]   data_mid_6_43_imag;
  reg        [17:0]   data_mid_6_44_real;
  reg        [17:0]   data_mid_6_44_imag;
  reg        [17:0]   data_mid_6_45_real;
  reg        [17:0]   data_mid_6_45_imag;
  reg        [17:0]   data_mid_6_46_real;
  reg        [17:0]   data_mid_6_46_imag;
  reg        [17:0]   data_mid_6_47_real;
  reg        [17:0]   data_mid_6_47_imag;
  reg        [17:0]   data_mid_6_48_real;
  reg        [17:0]   data_mid_6_48_imag;
  reg        [17:0]   data_mid_6_49_real;
  reg        [17:0]   data_mid_6_49_imag;
  reg        [17:0]   data_mid_6_50_real;
  reg        [17:0]   data_mid_6_50_imag;
  reg        [17:0]   data_mid_6_51_real;
  reg        [17:0]   data_mid_6_51_imag;
  reg        [17:0]   data_mid_6_52_real;
  reg        [17:0]   data_mid_6_52_imag;
  reg        [17:0]   data_mid_6_53_real;
  reg        [17:0]   data_mid_6_53_imag;
  reg        [17:0]   data_mid_6_54_real;
  reg        [17:0]   data_mid_6_54_imag;
  reg        [17:0]   data_mid_6_55_real;
  reg        [17:0]   data_mid_6_55_imag;
  reg        [17:0]   data_mid_6_56_real;
  reg        [17:0]   data_mid_6_56_imag;
  reg        [17:0]   data_mid_6_57_real;
  reg        [17:0]   data_mid_6_57_imag;
  reg        [17:0]   data_mid_6_58_real;
  reg        [17:0]   data_mid_6_58_imag;
  reg        [17:0]   data_mid_6_59_real;
  reg        [17:0]   data_mid_6_59_imag;
  reg        [17:0]   data_mid_6_60_real;
  reg        [17:0]   data_mid_6_60_imag;
  reg        [17:0]   data_mid_6_61_real;
  reg        [17:0]   data_mid_6_61_imag;
  reg        [17:0]   data_mid_6_62_real;
  reg        [17:0]   data_mid_6_62_imag;
  reg        [17:0]   data_mid_6_63_real;
  reg        [17:0]   data_mid_6_63_imag;
  wire       [35:0]   _zz_1;
  wire       [35:0]   _zz_2;
  wire       [35:0]   _zz_3;
  wire       [0:0]    _zz_4;
  wire       [0:0]    _zz_5;
  wire       [35:0]   _zz_6;
  wire       [35:0]   _zz_7;
  wire       [35:0]   _zz_8;
  wire       [0:0]    _zz_9;
  wire       [0:0]    _zz_10;
  wire       [35:0]   _zz_11;
  wire       [35:0]   _zz_12;
  wire       [35:0]   _zz_13;
  wire       [0:0]    _zz_14;
  wire       [0:0]    _zz_15;
  wire       [35:0]   _zz_16;
  wire       [35:0]   _zz_17;
  wire       [35:0]   _zz_18;
  wire       [0:0]    _zz_19;
  wire       [0:0]    _zz_20;
  wire       [35:0]   _zz_21;
  wire       [35:0]   _zz_22;
  wire       [35:0]   _zz_23;
  wire       [0:0]    _zz_24;
  wire       [0:0]    _zz_25;
  wire       [35:0]   _zz_26;
  wire       [35:0]   _zz_27;
  wire       [35:0]   _zz_28;
  wire       [0:0]    _zz_29;
  wire       [0:0]    _zz_30;
  wire       [35:0]   _zz_31;
  wire       [35:0]   _zz_32;
  wire       [35:0]   _zz_33;
  wire       [0:0]    _zz_34;
  wire       [0:0]    _zz_35;
  wire       [35:0]   _zz_36;
  wire       [35:0]   _zz_37;
  wire       [35:0]   _zz_38;
  wire       [0:0]    _zz_39;
  wire       [0:0]    _zz_40;
  wire       [35:0]   _zz_41;
  wire       [35:0]   _zz_42;
  wire       [35:0]   _zz_43;
  wire       [0:0]    _zz_44;
  wire       [0:0]    _zz_45;
  wire       [35:0]   _zz_46;
  wire       [35:0]   _zz_47;
  wire       [35:0]   _zz_48;
  wire       [0:0]    _zz_49;
  wire       [0:0]    _zz_50;
  wire       [35:0]   _zz_51;
  wire       [35:0]   _zz_52;
  wire       [35:0]   _zz_53;
  wire       [0:0]    _zz_54;
  wire       [0:0]    _zz_55;
  wire       [35:0]   _zz_56;
  wire       [35:0]   _zz_57;
  wire       [35:0]   _zz_58;
  wire       [0:0]    _zz_59;
  wire       [0:0]    _zz_60;
  wire       [35:0]   _zz_61;
  wire       [35:0]   _zz_62;
  wire       [35:0]   _zz_63;
  wire       [0:0]    _zz_64;
  wire       [0:0]    _zz_65;
  wire       [35:0]   _zz_66;
  wire       [35:0]   _zz_67;
  wire       [35:0]   _zz_68;
  wire       [0:0]    _zz_69;
  wire       [0:0]    _zz_70;
  wire       [35:0]   _zz_71;
  wire       [35:0]   _zz_72;
  wire       [35:0]   _zz_73;
  wire       [0:0]    _zz_74;
  wire       [0:0]    _zz_75;
  wire       [35:0]   _zz_76;
  wire       [35:0]   _zz_77;
  wire       [35:0]   _zz_78;
  wire       [0:0]    _zz_79;
  wire       [0:0]    _zz_80;
  wire       [35:0]   _zz_81;
  wire       [35:0]   _zz_82;
  wire       [35:0]   _zz_83;
  wire       [0:0]    _zz_84;
  wire       [0:0]    _zz_85;
  wire       [35:0]   _zz_86;
  wire       [35:0]   _zz_87;
  wire       [35:0]   _zz_88;
  wire       [0:0]    _zz_89;
  wire       [0:0]    _zz_90;
  wire       [35:0]   _zz_91;
  wire       [35:0]   _zz_92;
  wire       [35:0]   _zz_93;
  wire       [0:0]    _zz_94;
  wire       [0:0]    _zz_95;
  wire       [35:0]   _zz_96;
  wire       [35:0]   _zz_97;
  wire       [35:0]   _zz_98;
  wire       [0:0]    _zz_99;
  wire       [0:0]    _zz_100;
  wire       [35:0]   _zz_101;
  wire       [35:0]   _zz_102;
  wire       [35:0]   _zz_103;
  wire       [0:0]    _zz_104;
  wire       [0:0]    _zz_105;
  wire       [35:0]   _zz_106;
  wire       [35:0]   _zz_107;
  wire       [35:0]   _zz_108;
  wire       [0:0]    _zz_109;
  wire       [0:0]    _zz_110;
  wire       [35:0]   _zz_111;
  wire       [35:0]   _zz_112;
  wire       [35:0]   _zz_113;
  wire       [0:0]    _zz_114;
  wire       [0:0]    _zz_115;
  wire       [35:0]   _zz_116;
  wire       [35:0]   _zz_117;
  wire       [35:0]   _zz_118;
  wire       [0:0]    _zz_119;
  wire       [0:0]    _zz_120;
  wire       [35:0]   _zz_121;
  wire       [35:0]   _zz_122;
  wire       [35:0]   _zz_123;
  wire       [0:0]    _zz_124;
  wire       [0:0]    _zz_125;
  wire       [35:0]   _zz_126;
  wire       [35:0]   _zz_127;
  wire       [35:0]   _zz_128;
  wire       [0:0]    _zz_129;
  wire       [0:0]    _zz_130;
  wire       [35:0]   _zz_131;
  wire       [35:0]   _zz_132;
  wire       [35:0]   _zz_133;
  wire       [0:0]    _zz_134;
  wire       [0:0]    _zz_135;
  wire       [35:0]   _zz_136;
  wire       [35:0]   _zz_137;
  wire       [35:0]   _zz_138;
  wire       [0:0]    _zz_139;
  wire       [0:0]    _zz_140;
  wire       [35:0]   _zz_141;
  wire       [35:0]   _zz_142;
  wire       [35:0]   _zz_143;
  wire       [0:0]    _zz_144;
  wire       [0:0]    _zz_145;
  wire       [35:0]   _zz_146;
  wire       [35:0]   _zz_147;
  wire       [35:0]   _zz_148;
  wire       [0:0]    _zz_149;
  wire       [0:0]    _zz_150;
  wire       [35:0]   _zz_151;
  wire       [35:0]   _zz_152;
  wire       [35:0]   _zz_153;
  wire       [0:0]    _zz_154;
  wire       [0:0]    _zz_155;
  wire       [35:0]   _zz_156;
  wire       [35:0]   _zz_157;
  wire       [35:0]   _zz_158;
  wire       [0:0]    _zz_159;
  wire       [0:0]    _zz_160;
  wire       [35:0]   _zz_161;
  wire       [35:0]   _zz_162;
  wire       [35:0]   _zz_163;
  wire       [0:0]    _zz_164;
  wire       [0:0]    _zz_165;
  wire       [35:0]   _zz_166;
  wire       [35:0]   _zz_167;
  wire       [35:0]   _zz_168;
  wire       [0:0]    _zz_169;
  wire       [0:0]    _zz_170;
  wire       [35:0]   _zz_171;
  wire       [35:0]   _zz_172;
  wire       [35:0]   _zz_173;
  wire       [0:0]    _zz_174;
  wire       [0:0]    _zz_175;
  wire       [35:0]   _zz_176;
  wire       [35:0]   _zz_177;
  wire       [35:0]   _zz_178;
  wire       [0:0]    _zz_179;
  wire       [0:0]    _zz_180;
  wire       [35:0]   _zz_181;
  wire       [35:0]   _zz_182;
  wire       [35:0]   _zz_183;
  wire       [0:0]    _zz_184;
  wire       [0:0]    _zz_185;
  wire       [35:0]   _zz_186;
  wire       [35:0]   _zz_187;
  wire       [35:0]   _zz_188;
  wire       [0:0]    _zz_189;
  wire       [0:0]    _zz_190;
  wire       [35:0]   _zz_191;
  wire       [35:0]   _zz_192;
  wire       [35:0]   _zz_193;
  wire       [0:0]    _zz_194;
  wire       [0:0]    _zz_195;
  wire       [35:0]   _zz_196;
  wire       [35:0]   _zz_197;
  wire       [35:0]   _zz_198;
  wire       [0:0]    _zz_199;
  wire       [0:0]    _zz_200;
  wire       [35:0]   _zz_201;
  wire       [35:0]   _zz_202;
  wire       [35:0]   _zz_203;
  wire       [0:0]    _zz_204;
  wire       [0:0]    _zz_205;
  wire       [35:0]   _zz_206;
  wire       [35:0]   _zz_207;
  wire       [35:0]   _zz_208;
  wire       [0:0]    _zz_209;
  wire       [0:0]    _zz_210;
  wire       [35:0]   _zz_211;
  wire       [35:0]   _zz_212;
  wire       [35:0]   _zz_213;
  wire       [0:0]    _zz_214;
  wire       [0:0]    _zz_215;
  wire       [35:0]   _zz_216;
  wire       [35:0]   _zz_217;
  wire       [35:0]   _zz_218;
  wire       [0:0]    _zz_219;
  wire       [0:0]    _zz_220;
  wire       [35:0]   _zz_221;
  wire       [35:0]   _zz_222;
  wire       [35:0]   _zz_223;
  wire       [0:0]    _zz_224;
  wire       [0:0]    _zz_225;
  wire       [35:0]   _zz_226;
  wire       [35:0]   _zz_227;
  wire       [35:0]   _zz_228;
  wire       [0:0]    _zz_229;
  wire       [0:0]    _zz_230;
  wire       [35:0]   _zz_231;
  wire       [35:0]   _zz_232;
  wire       [35:0]   _zz_233;
  wire       [0:0]    _zz_234;
  wire       [0:0]    _zz_235;
  wire       [35:0]   _zz_236;
  wire       [35:0]   _zz_237;
  wire       [35:0]   _zz_238;
  wire       [0:0]    _zz_239;
  wire       [0:0]    _zz_240;
  wire       [35:0]   _zz_241;
  wire       [35:0]   _zz_242;
  wire       [35:0]   _zz_243;
  wire       [0:0]    _zz_244;
  wire       [0:0]    _zz_245;
  wire       [35:0]   _zz_246;
  wire       [35:0]   _zz_247;
  wire       [35:0]   _zz_248;
  wire       [0:0]    _zz_249;
  wire       [0:0]    _zz_250;
  wire       [35:0]   _zz_251;
  wire       [35:0]   _zz_252;
  wire       [35:0]   _zz_253;
  wire       [0:0]    _zz_254;
  wire       [0:0]    _zz_255;
  wire       [35:0]   _zz_256;
  wire       [35:0]   _zz_257;
  wire       [35:0]   _zz_258;
  wire       [0:0]    _zz_259;
  wire       [0:0]    _zz_260;
  wire       [35:0]   _zz_261;
  wire       [35:0]   _zz_262;
  wire       [35:0]   _zz_263;
  wire       [0:0]    _zz_264;
  wire       [0:0]    _zz_265;
  wire       [35:0]   _zz_266;
  wire       [35:0]   _zz_267;
  wire       [35:0]   _zz_268;
  wire       [0:0]    _zz_269;
  wire       [0:0]    _zz_270;
  wire       [35:0]   _zz_271;
  wire       [35:0]   _zz_272;
  wire       [35:0]   _zz_273;
  wire       [0:0]    _zz_274;
  wire       [0:0]    _zz_275;
  wire       [35:0]   _zz_276;
  wire       [35:0]   _zz_277;
  wire       [35:0]   _zz_278;
  wire       [0:0]    _zz_279;
  wire       [0:0]    _zz_280;
  wire       [35:0]   _zz_281;
  wire       [35:0]   _zz_282;
  wire       [35:0]   _zz_283;
  wire       [0:0]    _zz_284;
  wire       [0:0]    _zz_285;
  wire       [35:0]   _zz_286;
  wire       [35:0]   _zz_287;
  wire       [35:0]   _zz_288;
  wire       [0:0]    _zz_289;
  wire       [0:0]    _zz_290;
  wire       [35:0]   _zz_291;
  wire       [35:0]   _zz_292;
  wire       [35:0]   _zz_293;
  wire       [0:0]    _zz_294;
  wire       [0:0]    _zz_295;
  wire       [35:0]   _zz_296;
  wire       [35:0]   _zz_297;
  wire       [35:0]   _zz_298;
  wire       [0:0]    _zz_299;
  wire       [0:0]    _zz_300;
  wire       [35:0]   _zz_301;
  wire       [35:0]   _zz_302;
  wire       [35:0]   _zz_303;
  wire       [0:0]    _zz_304;
  wire       [0:0]    _zz_305;
  wire       [35:0]   _zz_306;
  wire       [35:0]   _zz_307;
  wire       [35:0]   _zz_308;
  wire       [0:0]    _zz_309;
  wire       [0:0]    _zz_310;
  wire       [35:0]   _zz_311;
  wire       [35:0]   _zz_312;
  wire       [35:0]   _zz_313;
  wire       [0:0]    _zz_314;
  wire       [0:0]    _zz_315;
  wire       [35:0]   _zz_316;
  wire       [35:0]   _zz_317;
  wire       [35:0]   _zz_318;
  wire       [0:0]    _zz_319;
  wire       [0:0]    _zz_320;
  wire       [35:0]   _zz_321;
  wire       [35:0]   _zz_322;
  wire       [35:0]   _zz_323;
  wire       [0:0]    _zz_324;
  wire       [0:0]    _zz_325;
  wire       [35:0]   _zz_326;
  wire       [35:0]   _zz_327;
  wire       [35:0]   _zz_328;
  wire       [0:0]    _zz_329;
  wire       [0:0]    _zz_330;
  wire       [35:0]   _zz_331;
  wire       [35:0]   _zz_332;
  wire       [35:0]   _zz_333;
  wire       [0:0]    _zz_334;
  wire       [0:0]    _zz_335;
  wire       [35:0]   _zz_336;
  wire       [35:0]   _zz_337;
  wire       [35:0]   _zz_338;
  wire       [0:0]    _zz_339;
  wire       [0:0]    _zz_340;
  wire       [35:0]   _zz_341;
  wire       [35:0]   _zz_342;
  wire       [35:0]   _zz_343;
  wire       [0:0]    _zz_344;
  wire       [0:0]    _zz_345;
  wire       [35:0]   _zz_346;
  wire       [35:0]   _zz_347;
  wire       [35:0]   _zz_348;
  wire       [0:0]    _zz_349;
  wire       [0:0]    _zz_350;
  wire       [35:0]   _zz_351;
  wire       [35:0]   _zz_352;
  wire       [35:0]   _zz_353;
  wire       [0:0]    _zz_354;
  wire       [0:0]    _zz_355;
  wire       [35:0]   _zz_356;
  wire       [35:0]   _zz_357;
  wire       [35:0]   _zz_358;
  wire       [0:0]    _zz_359;
  wire       [0:0]    _zz_360;
  wire       [35:0]   _zz_361;
  wire       [35:0]   _zz_362;
  wire       [35:0]   _zz_363;
  wire       [0:0]    _zz_364;
  wire       [0:0]    _zz_365;
  wire       [35:0]   _zz_366;
  wire       [35:0]   _zz_367;
  wire       [35:0]   _zz_368;
  wire       [0:0]    _zz_369;
  wire       [0:0]    _zz_370;
  wire       [35:0]   _zz_371;
  wire       [35:0]   _zz_372;
  wire       [35:0]   _zz_373;
  wire       [0:0]    _zz_374;
  wire       [0:0]    _zz_375;
  wire       [35:0]   _zz_376;
  wire       [35:0]   _zz_377;
  wire       [35:0]   _zz_378;
  wire       [0:0]    _zz_379;
  wire       [0:0]    _zz_380;
  wire       [35:0]   _zz_381;
  wire       [35:0]   _zz_382;
  wire       [35:0]   _zz_383;
  wire       [0:0]    _zz_384;
  wire       [0:0]    _zz_385;
  wire       [35:0]   _zz_386;
  wire       [35:0]   _zz_387;
  wire       [35:0]   _zz_388;
  wire       [0:0]    _zz_389;
  wire       [0:0]    _zz_390;
  wire       [35:0]   _zz_391;
  wire       [35:0]   _zz_392;
  wire       [35:0]   _zz_393;
  wire       [0:0]    _zz_394;
  wire       [0:0]    _zz_395;
  wire       [35:0]   _zz_396;
  wire       [35:0]   _zz_397;
  wire       [35:0]   _zz_398;
  wire       [0:0]    _zz_399;
  wire       [0:0]    _zz_400;
  wire       [35:0]   _zz_401;
  wire       [35:0]   _zz_402;
  wire       [35:0]   _zz_403;
  wire       [0:0]    _zz_404;
  wire       [0:0]    _zz_405;
  wire       [35:0]   _zz_406;
  wire       [35:0]   _zz_407;
  wire       [35:0]   _zz_408;
  wire       [0:0]    _zz_409;
  wire       [0:0]    _zz_410;
  wire       [35:0]   _zz_411;
  wire       [35:0]   _zz_412;
  wire       [35:0]   _zz_413;
  wire       [0:0]    _zz_414;
  wire       [0:0]    _zz_415;
  wire       [35:0]   _zz_416;
  wire       [35:0]   _zz_417;
  wire       [35:0]   _zz_418;
  wire       [0:0]    _zz_419;
  wire       [0:0]    _zz_420;
  wire       [35:0]   _zz_421;
  wire       [35:0]   _zz_422;
  wire       [35:0]   _zz_423;
  wire       [0:0]    _zz_424;
  wire       [0:0]    _zz_425;
  wire       [35:0]   _zz_426;
  wire       [35:0]   _zz_427;
  wire       [35:0]   _zz_428;
  wire       [0:0]    _zz_429;
  wire       [0:0]    _zz_430;
  wire       [35:0]   _zz_431;
  wire       [35:0]   _zz_432;
  wire       [35:0]   _zz_433;
  wire       [0:0]    _zz_434;
  wire       [0:0]    _zz_435;
  wire       [35:0]   _zz_436;
  wire       [35:0]   _zz_437;
  wire       [35:0]   _zz_438;
  wire       [0:0]    _zz_439;
  wire       [0:0]    _zz_440;
  wire       [35:0]   _zz_441;
  wire       [35:0]   _zz_442;
  wire       [35:0]   _zz_443;
  wire       [0:0]    _zz_444;
  wire       [0:0]    _zz_445;
  wire       [35:0]   _zz_446;
  wire       [35:0]   _zz_447;
  wire       [35:0]   _zz_448;
  wire       [0:0]    _zz_449;
  wire       [0:0]    _zz_450;
  wire       [35:0]   _zz_451;
  wire       [35:0]   _zz_452;
  wire       [35:0]   _zz_453;
  wire       [0:0]    _zz_454;
  wire       [0:0]    _zz_455;
  wire       [35:0]   _zz_456;
  wire       [35:0]   _zz_457;
  wire       [35:0]   _zz_458;
  wire       [0:0]    _zz_459;
  wire       [0:0]    _zz_460;
  wire       [35:0]   _zz_461;
  wire       [35:0]   _zz_462;
  wire       [35:0]   _zz_463;
  wire       [0:0]    _zz_464;
  wire       [0:0]    _zz_465;
  wire       [35:0]   _zz_466;
  wire       [35:0]   _zz_467;
  wire       [35:0]   _zz_468;
  wire       [0:0]    _zz_469;
  wire       [0:0]    _zz_470;
  wire       [35:0]   _zz_471;
  wire       [35:0]   _zz_472;
  wire       [35:0]   _zz_473;
  wire       [0:0]    _zz_474;
  wire       [0:0]    _zz_475;
  wire       [35:0]   _zz_476;
  wire       [35:0]   _zz_477;
  wire       [35:0]   _zz_478;
  wire       [0:0]    _zz_479;
  wire       [0:0]    _zz_480;
  wire       [35:0]   _zz_481;
  wire       [35:0]   _zz_482;
  wire       [35:0]   _zz_483;
  wire       [0:0]    _zz_484;
  wire       [0:0]    _zz_485;
  wire       [35:0]   _zz_486;
  wire       [35:0]   _zz_487;
  wire       [35:0]   _zz_488;
  wire       [0:0]    _zz_489;
  wire       [0:0]    _zz_490;
  wire       [35:0]   _zz_491;
  wire       [35:0]   _zz_492;
  wire       [35:0]   _zz_493;
  wire       [0:0]    _zz_494;
  wire       [0:0]    _zz_495;
  wire       [35:0]   _zz_496;
  wire       [35:0]   _zz_497;
  wire       [35:0]   _zz_498;
  wire       [0:0]    _zz_499;
  wire       [0:0]    _zz_500;
  wire       [35:0]   _zz_501;
  wire       [35:0]   _zz_502;
  wire       [35:0]   _zz_503;
  wire       [0:0]    _zz_504;
  wire       [0:0]    _zz_505;
  wire       [35:0]   _zz_506;
  wire       [35:0]   _zz_507;
  wire       [35:0]   _zz_508;
  wire       [0:0]    _zz_509;
  wire       [0:0]    _zz_510;
  wire       [35:0]   _zz_511;
  wire       [35:0]   _zz_512;
  wire       [35:0]   _zz_513;
  wire       [0:0]    _zz_514;
  wire       [0:0]    _zz_515;
  wire       [35:0]   _zz_516;
  wire       [35:0]   _zz_517;
  wire       [35:0]   _zz_518;
  wire       [0:0]    _zz_519;
  wire       [0:0]    _zz_520;
  wire       [35:0]   _zz_521;
  wire       [35:0]   _zz_522;
  wire       [35:0]   _zz_523;
  wire       [0:0]    _zz_524;
  wire       [0:0]    _zz_525;
  wire       [35:0]   _zz_526;
  wire       [35:0]   _zz_527;
  wire       [35:0]   _zz_528;
  wire       [0:0]    _zz_529;
  wire       [0:0]    _zz_530;
  wire       [35:0]   _zz_531;
  wire       [35:0]   _zz_532;
  wire       [35:0]   _zz_533;
  wire       [0:0]    _zz_534;
  wire       [0:0]    _zz_535;
  wire       [35:0]   _zz_536;
  wire       [35:0]   _zz_537;
  wire       [35:0]   _zz_538;
  wire       [0:0]    _zz_539;
  wire       [0:0]    _zz_540;
  wire       [35:0]   _zz_541;
  wire       [35:0]   _zz_542;
  wire       [35:0]   _zz_543;
  wire       [0:0]    _zz_544;
  wire       [0:0]    _zz_545;
  wire       [35:0]   _zz_546;
  wire       [35:0]   _zz_547;
  wire       [35:0]   _zz_548;
  wire       [0:0]    _zz_549;
  wire       [0:0]    _zz_550;
  wire       [35:0]   _zz_551;
  wire       [35:0]   _zz_552;
  wire       [35:0]   _zz_553;
  wire       [0:0]    _zz_554;
  wire       [0:0]    _zz_555;
  wire       [35:0]   _zz_556;
  wire       [35:0]   _zz_557;
  wire       [35:0]   _zz_558;
  wire       [0:0]    _zz_559;
  wire       [0:0]    _zz_560;
  wire       [35:0]   _zz_561;
  wire       [35:0]   _zz_562;
  wire       [35:0]   _zz_563;
  wire       [0:0]    _zz_564;
  wire       [0:0]    _zz_565;
  wire       [35:0]   _zz_566;
  wire       [35:0]   _zz_567;
  wire       [35:0]   _zz_568;
  wire       [0:0]    _zz_569;
  wire       [0:0]    _zz_570;
  wire       [35:0]   _zz_571;
  wire       [35:0]   _zz_572;
  wire       [35:0]   _zz_573;
  wire       [0:0]    _zz_574;
  wire       [0:0]    _zz_575;
  wire       [35:0]   _zz_576;
  wire       [35:0]   _zz_577;
  wire       [35:0]   _zz_578;
  wire       [0:0]    _zz_579;
  wire       [0:0]    _zz_580;
  wire       [35:0]   _zz_581;
  wire       [35:0]   _zz_582;
  wire       [35:0]   _zz_583;
  wire       [0:0]    _zz_584;
  wire       [0:0]    _zz_585;
  wire       [35:0]   _zz_586;
  wire       [35:0]   _zz_587;
  wire       [35:0]   _zz_588;
  wire       [0:0]    _zz_589;
  wire       [0:0]    _zz_590;
  wire       [35:0]   _zz_591;
  wire       [35:0]   _zz_592;
  wire       [35:0]   _zz_593;
  wire       [0:0]    _zz_594;
  wire       [0:0]    _zz_595;
  wire       [35:0]   _zz_596;
  wire       [35:0]   _zz_597;
  wire       [35:0]   _zz_598;
  wire       [0:0]    _zz_599;
  wire       [0:0]    _zz_600;
  wire       [35:0]   _zz_601;
  wire       [35:0]   _zz_602;
  wire       [35:0]   _zz_603;
  wire       [0:0]    _zz_604;
  wire       [0:0]    _zz_605;
  wire       [35:0]   _zz_606;
  wire       [35:0]   _zz_607;
  wire       [35:0]   _zz_608;
  wire       [0:0]    _zz_609;
  wire       [0:0]    _zz_610;
  wire       [35:0]   _zz_611;
  wire       [35:0]   _zz_612;
  wire       [35:0]   _zz_613;
  wire       [0:0]    _zz_614;
  wire       [0:0]    _zz_615;
  wire       [35:0]   _zz_616;
  wire       [35:0]   _zz_617;
  wire       [35:0]   _zz_618;
  wire       [0:0]    _zz_619;
  wire       [0:0]    _zz_620;
  wire       [35:0]   _zz_621;
  wire       [35:0]   _zz_622;
  wire       [35:0]   _zz_623;
  wire       [0:0]    _zz_624;
  wire       [0:0]    _zz_625;
  wire       [35:0]   _zz_626;
  wire       [35:0]   _zz_627;
  wire       [35:0]   _zz_628;
  wire       [0:0]    _zz_629;
  wire       [0:0]    _zz_630;
  wire       [35:0]   _zz_631;
  wire       [35:0]   _zz_632;
  wire       [35:0]   _zz_633;
  wire       [0:0]    _zz_634;
  wire       [0:0]    _zz_635;
  wire       [35:0]   _zz_636;
  wire       [35:0]   _zz_637;
  wire       [35:0]   _zz_638;
  wire       [0:0]    _zz_639;
  wire       [0:0]    _zz_640;
  wire       [35:0]   _zz_641;
  wire       [35:0]   _zz_642;
  wire       [35:0]   _zz_643;
  wire       [0:0]    _zz_644;
  wire       [0:0]    _zz_645;
  wire       [35:0]   _zz_646;
  wire       [35:0]   _zz_647;
  wire       [35:0]   _zz_648;
  wire       [0:0]    _zz_649;
  wire       [0:0]    _zz_650;
  wire       [35:0]   _zz_651;
  wire       [35:0]   _zz_652;
  wire       [35:0]   _zz_653;
  wire       [0:0]    _zz_654;
  wire       [0:0]    _zz_655;
  wire       [35:0]   _zz_656;
  wire       [35:0]   _zz_657;
  wire       [35:0]   _zz_658;
  wire       [0:0]    _zz_659;
  wire       [0:0]    _zz_660;
  wire       [35:0]   _zz_661;
  wire       [35:0]   _zz_662;
  wire       [35:0]   _zz_663;
  wire       [0:0]    _zz_664;
  wire       [0:0]    _zz_665;
  wire       [35:0]   _zz_666;
  wire       [35:0]   _zz_667;
  wire       [35:0]   _zz_668;
  wire       [0:0]    _zz_669;
  wire       [0:0]    _zz_670;
  wire       [35:0]   _zz_671;
  wire       [35:0]   _zz_672;
  wire       [35:0]   _zz_673;
  wire       [0:0]    _zz_674;
  wire       [0:0]    _zz_675;
  wire       [35:0]   _zz_676;
  wire       [35:0]   _zz_677;
  wire       [35:0]   _zz_678;
  wire       [0:0]    _zz_679;
  wire       [0:0]    _zz_680;
  wire       [35:0]   _zz_681;
  wire       [35:0]   _zz_682;
  wire       [35:0]   _zz_683;
  wire       [0:0]    _zz_684;
  wire       [0:0]    _zz_685;
  wire       [35:0]   _zz_686;
  wire       [35:0]   _zz_687;
  wire       [35:0]   _zz_688;
  wire       [0:0]    _zz_689;
  wire       [0:0]    _zz_690;
  wire       [35:0]   _zz_691;
  wire       [35:0]   _zz_692;
  wire       [35:0]   _zz_693;
  wire       [0:0]    _zz_694;
  wire       [0:0]    _zz_695;
  wire       [35:0]   _zz_696;
  wire       [35:0]   _zz_697;
  wire       [35:0]   _zz_698;
  wire       [0:0]    _zz_699;
  wire       [0:0]    _zz_700;
  wire       [35:0]   _zz_701;
  wire       [35:0]   _zz_702;
  wire       [35:0]   _zz_703;
  wire       [0:0]    _zz_704;
  wire       [0:0]    _zz_705;
  wire       [35:0]   _zz_706;
  wire       [35:0]   _zz_707;
  wire       [35:0]   _zz_708;
  wire       [0:0]    _zz_709;
  wire       [0:0]    _zz_710;
  wire       [35:0]   _zz_711;
  wire       [35:0]   _zz_712;
  wire       [35:0]   _zz_713;
  wire       [0:0]    _zz_714;
  wire       [0:0]    _zz_715;
  wire       [35:0]   _zz_716;
  wire       [35:0]   _zz_717;
  wire       [35:0]   _zz_718;
  wire       [0:0]    _zz_719;
  wire       [0:0]    _zz_720;
  wire       [35:0]   _zz_721;
  wire       [35:0]   _zz_722;
  wire       [35:0]   _zz_723;
  wire       [0:0]    _zz_724;
  wire       [0:0]    _zz_725;
  wire       [35:0]   _zz_726;
  wire       [35:0]   _zz_727;
  wire       [35:0]   _zz_728;
  wire       [0:0]    _zz_729;
  wire       [0:0]    _zz_730;
  wire       [35:0]   _zz_731;
  wire       [35:0]   _zz_732;
  wire       [35:0]   _zz_733;
  wire       [0:0]    _zz_734;
  wire       [0:0]    _zz_735;
  wire       [35:0]   _zz_736;
  wire       [35:0]   _zz_737;
  wire       [35:0]   _zz_738;
  wire       [0:0]    _zz_739;
  wire       [0:0]    _zz_740;
  wire       [35:0]   _zz_741;
  wire       [35:0]   _zz_742;
  wire       [35:0]   _zz_743;
  wire       [0:0]    _zz_744;
  wire       [0:0]    _zz_745;
  wire       [35:0]   _zz_746;
  wire       [35:0]   _zz_747;
  wire       [35:0]   _zz_748;
  wire       [0:0]    _zz_749;
  wire       [0:0]    _zz_750;
  wire       [35:0]   _zz_751;
  wire       [35:0]   _zz_752;
  wire       [35:0]   _zz_753;
  wire       [0:0]    _zz_754;
  wire       [0:0]    _zz_755;
  wire       [35:0]   _zz_756;
  wire       [35:0]   _zz_757;
  wire       [35:0]   _zz_758;
  wire       [0:0]    _zz_759;
  wire       [0:0]    _zz_760;
  wire       [35:0]   _zz_761;
  wire       [35:0]   _zz_762;
  wire       [35:0]   _zz_763;
  wire       [0:0]    _zz_764;
  wire       [0:0]    _zz_765;
  wire       [35:0]   _zz_766;
  wire       [35:0]   _zz_767;
  wire       [35:0]   _zz_768;
  wire       [0:0]    _zz_769;
  wire       [0:0]    _zz_770;
  wire       [35:0]   _zz_771;
  wire       [35:0]   _zz_772;
  wire       [35:0]   _zz_773;
  wire       [0:0]    _zz_774;
  wire       [0:0]    _zz_775;
  wire       [35:0]   _zz_776;
  wire       [35:0]   _zz_777;
  wire       [35:0]   _zz_778;
  wire       [0:0]    _zz_779;
  wire       [0:0]    _zz_780;
  wire       [35:0]   _zz_781;
  wire       [35:0]   _zz_782;
  wire       [35:0]   _zz_783;
  wire       [0:0]    _zz_784;
  wire       [0:0]    _zz_785;
  wire       [35:0]   _zz_786;
  wire       [35:0]   _zz_787;
  wire       [35:0]   _zz_788;
  wire       [0:0]    _zz_789;
  wire       [0:0]    _zz_790;
  wire       [35:0]   _zz_791;
  wire       [35:0]   _zz_792;
  wire       [35:0]   _zz_793;
  wire       [0:0]    _zz_794;
  wire       [0:0]    _zz_795;
  wire       [35:0]   _zz_796;
  wire       [35:0]   _zz_797;
  wire       [35:0]   _zz_798;
  wire       [0:0]    _zz_799;
  wire       [0:0]    _zz_800;
  wire       [35:0]   _zz_801;
  wire       [35:0]   _zz_802;
  wire       [35:0]   _zz_803;
  wire       [0:0]    _zz_804;
  wire       [0:0]    _zz_805;
  wire       [35:0]   _zz_806;
  wire       [35:0]   _zz_807;
  wire       [35:0]   _zz_808;
  wire       [0:0]    _zz_809;
  wire       [0:0]    _zz_810;
  wire       [35:0]   _zz_811;
  wire       [35:0]   _zz_812;
  wire       [35:0]   _zz_813;
  wire       [0:0]    _zz_814;
  wire       [0:0]    _zz_815;
  wire       [35:0]   _zz_816;
  wire       [35:0]   _zz_817;
  wire       [35:0]   _zz_818;
  wire       [0:0]    _zz_819;
  wire       [0:0]    _zz_820;
  wire       [35:0]   _zz_821;
  wire       [35:0]   _zz_822;
  wire       [35:0]   _zz_823;
  wire       [0:0]    _zz_824;
  wire       [0:0]    _zz_825;
  wire       [35:0]   _zz_826;
  wire       [35:0]   _zz_827;
  wire       [35:0]   _zz_828;
  wire       [0:0]    _zz_829;
  wire       [0:0]    _zz_830;
  wire       [35:0]   _zz_831;
  wire       [35:0]   _zz_832;
  wire       [35:0]   _zz_833;
  wire       [0:0]    _zz_834;
  wire       [0:0]    _zz_835;
  wire       [35:0]   _zz_836;
  wire       [35:0]   _zz_837;
  wire       [35:0]   _zz_838;
  wire       [0:0]    _zz_839;
  wire       [0:0]    _zz_840;
  wire       [35:0]   _zz_841;
  wire       [35:0]   _zz_842;
  wire       [35:0]   _zz_843;
  wire       [0:0]    _zz_844;
  wire       [0:0]    _zz_845;
  wire       [35:0]   _zz_846;
  wire       [35:0]   _zz_847;
  wire       [35:0]   _zz_848;
  wire       [0:0]    _zz_849;
  wire       [0:0]    _zz_850;
  wire       [35:0]   _zz_851;
  wire       [35:0]   _zz_852;
  wire       [35:0]   _zz_853;
  wire       [0:0]    _zz_854;
  wire       [0:0]    _zz_855;
  wire       [35:0]   _zz_856;
  wire       [35:0]   _zz_857;
  wire       [35:0]   _zz_858;
  wire       [0:0]    _zz_859;
  wire       [0:0]    _zz_860;
  wire       [35:0]   _zz_861;
  wire       [35:0]   _zz_862;
  wire       [35:0]   _zz_863;
  wire       [0:0]    _zz_864;
  wire       [0:0]    _zz_865;
  wire       [35:0]   _zz_866;
  wire       [35:0]   _zz_867;
  wire       [35:0]   _zz_868;
  wire       [0:0]    _zz_869;
  wire       [0:0]    _zz_870;
  wire       [35:0]   _zz_871;
  wire       [35:0]   _zz_872;
  wire       [35:0]   _zz_873;
  wire       [0:0]    _zz_874;
  wire       [0:0]    _zz_875;
  wire       [35:0]   _zz_876;
  wire       [35:0]   _zz_877;
  wire       [35:0]   _zz_878;
  wire       [0:0]    _zz_879;
  wire       [0:0]    _zz_880;
  wire       [35:0]   _zz_881;
  wire       [35:0]   _zz_882;
  wire       [35:0]   _zz_883;
  wire       [0:0]    _zz_884;
  wire       [0:0]    _zz_885;
  wire       [35:0]   _zz_886;
  wire       [35:0]   _zz_887;
  wire       [35:0]   _zz_888;
  wire       [0:0]    _zz_889;
  wire       [0:0]    _zz_890;
  wire       [35:0]   _zz_891;
  wire       [35:0]   _zz_892;
  wire       [35:0]   _zz_893;
  wire       [0:0]    _zz_894;
  wire       [0:0]    _zz_895;
  wire       [35:0]   _zz_896;
  wire       [35:0]   _zz_897;
  wire       [35:0]   _zz_898;
  wire       [0:0]    _zz_899;
  wire       [0:0]    _zz_900;
  wire       [35:0]   _zz_901;
  wire       [35:0]   _zz_902;
  wire       [35:0]   _zz_903;
  wire       [0:0]    _zz_904;
  wire       [0:0]    _zz_905;
  wire       [35:0]   _zz_906;
  wire       [35:0]   _zz_907;
  wire       [35:0]   _zz_908;
  wire       [0:0]    _zz_909;
  wire       [0:0]    _zz_910;
  wire       [35:0]   _zz_911;
  wire       [35:0]   _zz_912;
  wire       [35:0]   _zz_913;
  wire       [0:0]    _zz_914;
  wire       [0:0]    _zz_915;
  wire       [35:0]   _zz_916;
  wire       [35:0]   _zz_917;
  wire       [35:0]   _zz_918;
  wire       [0:0]    _zz_919;
  wire       [0:0]    _zz_920;
  wire       [35:0]   _zz_921;
  wire       [35:0]   _zz_922;
  wire       [35:0]   _zz_923;
  wire       [0:0]    _zz_924;
  wire       [0:0]    _zz_925;
  wire       [35:0]   _zz_926;
  wire       [35:0]   _zz_927;
  wire       [35:0]   _zz_928;
  wire       [0:0]    _zz_929;
  wire       [0:0]    _zz_930;
  wire       [35:0]   _zz_931;
  wire       [35:0]   _zz_932;
  wire       [35:0]   _zz_933;
  wire       [0:0]    _zz_934;
  wire       [0:0]    _zz_935;
  wire       [35:0]   _zz_936;
  wire       [35:0]   _zz_937;
  wire       [35:0]   _zz_938;
  wire       [0:0]    _zz_939;
  wire       [0:0]    _zz_940;
  wire       [35:0]   _zz_941;
  wire       [35:0]   _zz_942;
  wire       [35:0]   _zz_943;
  wire       [0:0]    _zz_944;
  wire       [0:0]    _zz_945;
  wire       [35:0]   _zz_946;
  wire       [35:0]   _zz_947;
  wire       [35:0]   _zz_948;
  wire       [0:0]    _zz_949;
  wire       [0:0]    _zz_950;
  wire       [35:0]   _zz_951;
  wire       [35:0]   _zz_952;
  wire       [35:0]   _zz_953;
  wire       [0:0]    _zz_954;
  wire       [0:0]    _zz_955;
  wire       [35:0]   _zz_956;
  wire       [35:0]   _zz_957;
  wire       [35:0]   _zz_958;
  wire       [0:0]    _zz_959;
  wire       [0:0]    _zz_960;
  reg                 io_data_in_valid_delay_1;
  reg                 io_data_in_valid_delay_2;
  reg                 io_data_in_valid_delay_3;
  reg                 io_data_in_valid_delay_4;
  reg                 io_data_in_valid_delay_5;
  reg                 io_data_in_valid_delay_6;
  reg                 io_data_in_valid_delay_7;
  reg                 io_data_in_valid_delay_8;

  assign _zz_2113 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2114 = ($signed(_zz_3) - $signed(_zz_2115));
  assign _zz_2115 = ($signed(_zz_2116) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2116 = ($signed(data_mid_0_1_real) + $signed(data_mid_0_1_imag));
  assign _zz_2117 = fixTo_dout;
  assign _zz_2118 = ($signed(_zz_3) + $signed(_zz_2119));
  assign _zz_2119 = ($signed(_zz_2120) * $signed(twiddle_factor_table_0_real));
  assign _zz_2120 = ($signed(data_mid_0_1_imag) - $signed(data_mid_0_1_real));
  assign _zz_2121 = fixTo_1_dout;
  assign _zz_2122 = _zz_2123[35 : 0];
  assign _zz_2123 = _zz_2124;
  assign _zz_2124 = ($signed(_zz_2125) >>> _zz_4);
  assign _zz_2125 = _zz_2126;
  assign _zz_2126 = ($signed(_zz_2128) - $signed(_zz_1));
  assign _zz_2127 = ({9'd0,data_mid_0_0_real} <<< 9);
  assign _zz_2128 = {{9{_zz_2127[26]}}, _zz_2127};
  assign _zz_2129 = fixTo_2_dout;
  assign _zz_2130 = _zz_2131[35 : 0];
  assign _zz_2131 = _zz_2132;
  assign _zz_2132 = ($signed(_zz_2133) >>> _zz_4);
  assign _zz_2133 = _zz_2134;
  assign _zz_2134 = ($signed(_zz_2136) - $signed(_zz_2));
  assign _zz_2135 = ({9'd0,data_mid_0_0_imag} <<< 9);
  assign _zz_2136 = {{9{_zz_2135[26]}}, _zz_2135};
  assign _zz_2137 = fixTo_3_dout;
  assign _zz_2138 = _zz_2139[35 : 0];
  assign _zz_2139 = _zz_2140;
  assign _zz_2140 = ($signed(_zz_2141) >>> _zz_5);
  assign _zz_2141 = _zz_2142;
  assign _zz_2142 = ($signed(_zz_2144) + $signed(_zz_1));
  assign _zz_2143 = ({9'd0,data_mid_0_0_real} <<< 9);
  assign _zz_2144 = {{9{_zz_2143[26]}}, _zz_2143};
  assign _zz_2145 = fixTo_4_dout;
  assign _zz_2146 = _zz_2147[35 : 0];
  assign _zz_2147 = _zz_2148;
  assign _zz_2148 = ($signed(_zz_2149) >>> _zz_5);
  assign _zz_2149 = _zz_2150;
  assign _zz_2150 = ($signed(_zz_2152) + $signed(_zz_2));
  assign _zz_2151 = ({9'd0,data_mid_0_0_imag} <<< 9);
  assign _zz_2152 = {{9{_zz_2151[26]}}, _zz_2151};
  assign _zz_2153 = fixTo_5_dout;
  assign _zz_2154 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2155 = ($signed(_zz_8) - $signed(_zz_2156));
  assign _zz_2156 = ($signed(_zz_2157) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2157 = ($signed(data_mid_0_3_real) + $signed(data_mid_0_3_imag));
  assign _zz_2158 = fixTo_6_dout;
  assign _zz_2159 = ($signed(_zz_8) + $signed(_zz_2160));
  assign _zz_2160 = ($signed(_zz_2161) * $signed(twiddle_factor_table_0_real));
  assign _zz_2161 = ($signed(data_mid_0_3_imag) - $signed(data_mid_0_3_real));
  assign _zz_2162 = fixTo_7_dout;
  assign _zz_2163 = _zz_2164[35 : 0];
  assign _zz_2164 = _zz_2165;
  assign _zz_2165 = ($signed(_zz_2166) >>> _zz_9);
  assign _zz_2166 = _zz_2167;
  assign _zz_2167 = ($signed(_zz_2169) - $signed(_zz_6));
  assign _zz_2168 = ({9'd0,data_mid_0_2_real} <<< 9);
  assign _zz_2169 = {{9{_zz_2168[26]}}, _zz_2168};
  assign _zz_2170 = fixTo_8_dout;
  assign _zz_2171 = _zz_2172[35 : 0];
  assign _zz_2172 = _zz_2173;
  assign _zz_2173 = ($signed(_zz_2174) >>> _zz_9);
  assign _zz_2174 = _zz_2175;
  assign _zz_2175 = ($signed(_zz_2177) - $signed(_zz_7));
  assign _zz_2176 = ({9'd0,data_mid_0_2_imag} <<< 9);
  assign _zz_2177 = {{9{_zz_2176[26]}}, _zz_2176};
  assign _zz_2178 = fixTo_9_dout;
  assign _zz_2179 = _zz_2180[35 : 0];
  assign _zz_2180 = _zz_2181;
  assign _zz_2181 = ($signed(_zz_2182) >>> _zz_10);
  assign _zz_2182 = _zz_2183;
  assign _zz_2183 = ($signed(_zz_2185) + $signed(_zz_6));
  assign _zz_2184 = ({9'd0,data_mid_0_2_real} <<< 9);
  assign _zz_2185 = {{9{_zz_2184[26]}}, _zz_2184};
  assign _zz_2186 = fixTo_10_dout;
  assign _zz_2187 = _zz_2188[35 : 0];
  assign _zz_2188 = _zz_2189;
  assign _zz_2189 = ($signed(_zz_2190) >>> _zz_10);
  assign _zz_2190 = _zz_2191;
  assign _zz_2191 = ($signed(_zz_2193) + $signed(_zz_7));
  assign _zz_2192 = ({9'd0,data_mid_0_2_imag} <<< 9);
  assign _zz_2193 = {{9{_zz_2192[26]}}, _zz_2192};
  assign _zz_2194 = fixTo_11_dout;
  assign _zz_2195 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2196 = ($signed(_zz_13) - $signed(_zz_2197));
  assign _zz_2197 = ($signed(_zz_2198) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2198 = ($signed(data_mid_0_5_real) + $signed(data_mid_0_5_imag));
  assign _zz_2199 = fixTo_12_dout;
  assign _zz_2200 = ($signed(_zz_13) + $signed(_zz_2201));
  assign _zz_2201 = ($signed(_zz_2202) * $signed(twiddle_factor_table_0_real));
  assign _zz_2202 = ($signed(data_mid_0_5_imag) - $signed(data_mid_0_5_real));
  assign _zz_2203 = fixTo_13_dout;
  assign _zz_2204 = _zz_2205[35 : 0];
  assign _zz_2205 = _zz_2206;
  assign _zz_2206 = ($signed(_zz_2207) >>> _zz_14);
  assign _zz_2207 = _zz_2208;
  assign _zz_2208 = ($signed(_zz_2210) - $signed(_zz_11));
  assign _zz_2209 = ({9'd0,data_mid_0_4_real} <<< 9);
  assign _zz_2210 = {{9{_zz_2209[26]}}, _zz_2209};
  assign _zz_2211 = fixTo_14_dout;
  assign _zz_2212 = _zz_2213[35 : 0];
  assign _zz_2213 = _zz_2214;
  assign _zz_2214 = ($signed(_zz_2215) >>> _zz_14);
  assign _zz_2215 = _zz_2216;
  assign _zz_2216 = ($signed(_zz_2218) - $signed(_zz_12));
  assign _zz_2217 = ({9'd0,data_mid_0_4_imag} <<< 9);
  assign _zz_2218 = {{9{_zz_2217[26]}}, _zz_2217};
  assign _zz_2219 = fixTo_15_dout;
  assign _zz_2220 = _zz_2221[35 : 0];
  assign _zz_2221 = _zz_2222;
  assign _zz_2222 = ($signed(_zz_2223) >>> _zz_15);
  assign _zz_2223 = _zz_2224;
  assign _zz_2224 = ($signed(_zz_2226) + $signed(_zz_11));
  assign _zz_2225 = ({9'd0,data_mid_0_4_real} <<< 9);
  assign _zz_2226 = {{9{_zz_2225[26]}}, _zz_2225};
  assign _zz_2227 = fixTo_16_dout;
  assign _zz_2228 = _zz_2229[35 : 0];
  assign _zz_2229 = _zz_2230;
  assign _zz_2230 = ($signed(_zz_2231) >>> _zz_15);
  assign _zz_2231 = _zz_2232;
  assign _zz_2232 = ($signed(_zz_2234) + $signed(_zz_12));
  assign _zz_2233 = ({9'd0,data_mid_0_4_imag} <<< 9);
  assign _zz_2234 = {{9{_zz_2233[26]}}, _zz_2233};
  assign _zz_2235 = fixTo_17_dout;
  assign _zz_2236 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2237 = ($signed(_zz_18) - $signed(_zz_2238));
  assign _zz_2238 = ($signed(_zz_2239) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2239 = ($signed(data_mid_0_7_real) + $signed(data_mid_0_7_imag));
  assign _zz_2240 = fixTo_18_dout;
  assign _zz_2241 = ($signed(_zz_18) + $signed(_zz_2242));
  assign _zz_2242 = ($signed(_zz_2243) * $signed(twiddle_factor_table_0_real));
  assign _zz_2243 = ($signed(data_mid_0_7_imag) - $signed(data_mid_0_7_real));
  assign _zz_2244 = fixTo_19_dout;
  assign _zz_2245 = _zz_2246[35 : 0];
  assign _zz_2246 = _zz_2247;
  assign _zz_2247 = ($signed(_zz_2248) >>> _zz_19);
  assign _zz_2248 = _zz_2249;
  assign _zz_2249 = ($signed(_zz_2251) - $signed(_zz_16));
  assign _zz_2250 = ({9'd0,data_mid_0_6_real} <<< 9);
  assign _zz_2251 = {{9{_zz_2250[26]}}, _zz_2250};
  assign _zz_2252 = fixTo_20_dout;
  assign _zz_2253 = _zz_2254[35 : 0];
  assign _zz_2254 = _zz_2255;
  assign _zz_2255 = ($signed(_zz_2256) >>> _zz_19);
  assign _zz_2256 = _zz_2257;
  assign _zz_2257 = ($signed(_zz_2259) - $signed(_zz_17));
  assign _zz_2258 = ({9'd0,data_mid_0_6_imag} <<< 9);
  assign _zz_2259 = {{9{_zz_2258[26]}}, _zz_2258};
  assign _zz_2260 = fixTo_21_dout;
  assign _zz_2261 = _zz_2262[35 : 0];
  assign _zz_2262 = _zz_2263;
  assign _zz_2263 = ($signed(_zz_2264) >>> _zz_20);
  assign _zz_2264 = _zz_2265;
  assign _zz_2265 = ($signed(_zz_2267) + $signed(_zz_16));
  assign _zz_2266 = ({9'd0,data_mid_0_6_real} <<< 9);
  assign _zz_2267 = {{9{_zz_2266[26]}}, _zz_2266};
  assign _zz_2268 = fixTo_22_dout;
  assign _zz_2269 = _zz_2270[35 : 0];
  assign _zz_2270 = _zz_2271;
  assign _zz_2271 = ($signed(_zz_2272) >>> _zz_20);
  assign _zz_2272 = _zz_2273;
  assign _zz_2273 = ($signed(_zz_2275) + $signed(_zz_17));
  assign _zz_2274 = ({9'd0,data_mid_0_6_imag} <<< 9);
  assign _zz_2275 = {{9{_zz_2274[26]}}, _zz_2274};
  assign _zz_2276 = fixTo_23_dout;
  assign _zz_2277 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2278 = ($signed(_zz_23) - $signed(_zz_2279));
  assign _zz_2279 = ($signed(_zz_2280) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2280 = ($signed(data_mid_0_9_real) + $signed(data_mid_0_9_imag));
  assign _zz_2281 = fixTo_24_dout;
  assign _zz_2282 = ($signed(_zz_23) + $signed(_zz_2283));
  assign _zz_2283 = ($signed(_zz_2284) * $signed(twiddle_factor_table_0_real));
  assign _zz_2284 = ($signed(data_mid_0_9_imag) - $signed(data_mid_0_9_real));
  assign _zz_2285 = fixTo_25_dout;
  assign _zz_2286 = _zz_2287[35 : 0];
  assign _zz_2287 = _zz_2288;
  assign _zz_2288 = ($signed(_zz_2289) >>> _zz_24);
  assign _zz_2289 = _zz_2290;
  assign _zz_2290 = ($signed(_zz_2292) - $signed(_zz_21));
  assign _zz_2291 = ({9'd0,data_mid_0_8_real} <<< 9);
  assign _zz_2292 = {{9{_zz_2291[26]}}, _zz_2291};
  assign _zz_2293 = fixTo_26_dout;
  assign _zz_2294 = _zz_2295[35 : 0];
  assign _zz_2295 = _zz_2296;
  assign _zz_2296 = ($signed(_zz_2297) >>> _zz_24);
  assign _zz_2297 = _zz_2298;
  assign _zz_2298 = ($signed(_zz_2300) - $signed(_zz_22));
  assign _zz_2299 = ({9'd0,data_mid_0_8_imag} <<< 9);
  assign _zz_2300 = {{9{_zz_2299[26]}}, _zz_2299};
  assign _zz_2301 = fixTo_27_dout;
  assign _zz_2302 = _zz_2303[35 : 0];
  assign _zz_2303 = _zz_2304;
  assign _zz_2304 = ($signed(_zz_2305) >>> _zz_25);
  assign _zz_2305 = _zz_2306;
  assign _zz_2306 = ($signed(_zz_2308) + $signed(_zz_21));
  assign _zz_2307 = ({9'd0,data_mid_0_8_real} <<< 9);
  assign _zz_2308 = {{9{_zz_2307[26]}}, _zz_2307};
  assign _zz_2309 = fixTo_28_dout;
  assign _zz_2310 = _zz_2311[35 : 0];
  assign _zz_2311 = _zz_2312;
  assign _zz_2312 = ($signed(_zz_2313) >>> _zz_25);
  assign _zz_2313 = _zz_2314;
  assign _zz_2314 = ($signed(_zz_2316) + $signed(_zz_22));
  assign _zz_2315 = ({9'd0,data_mid_0_8_imag} <<< 9);
  assign _zz_2316 = {{9{_zz_2315[26]}}, _zz_2315};
  assign _zz_2317 = fixTo_29_dout;
  assign _zz_2318 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2319 = ($signed(_zz_28) - $signed(_zz_2320));
  assign _zz_2320 = ($signed(_zz_2321) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2321 = ($signed(data_mid_0_11_real) + $signed(data_mid_0_11_imag));
  assign _zz_2322 = fixTo_30_dout;
  assign _zz_2323 = ($signed(_zz_28) + $signed(_zz_2324));
  assign _zz_2324 = ($signed(_zz_2325) * $signed(twiddle_factor_table_0_real));
  assign _zz_2325 = ($signed(data_mid_0_11_imag) - $signed(data_mid_0_11_real));
  assign _zz_2326 = fixTo_31_dout;
  assign _zz_2327 = _zz_2328[35 : 0];
  assign _zz_2328 = _zz_2329;
  assign _zz_2329 = ($signed(_zz_2330) >>> _zz_29);
  assign _zz_2330 = _zz_2331;
  assign _zz_2331 = ($signed(_zz_2333) - $signed(_zz_26));
  assign _zz_2332 = ({9'd0,data_mid_0_10_real} <<< 9);
  assign _zz_2333 = {{9{_zz_2332[26]}}, _zz_2332};
  assign _zz_2334 = fixTo_32_dout;
  assign _zz_2335 = _zz_2336[35 : 0];
  assign _zz_2336 = _zz_2337;
  assign _zz_2337 = ($signed(_zz_2338) >>> _zz_29);
  assign _zz_2338 = _zz_2339;
  assign _zz_2339 = ($signed(_zz_2341) - $signed(_zz_27));
  assign _zz_2340 = ({9'd0,data_mid_0_10_imag} <<< 9);
  assign _zz_2341 = {{9{_zz_2340[26]}}, _zz_2340};
  assign _zz_2342 = fixTo_33_dout;
  assign _zz_2343 = _zz_2344[35 : 0];
  assign _zz_2344 = _zz_2345;
  assign _zz_2345 = ($signed(_zz_2346) >>> _zz_30);
  assign _zz_2346 = _zz_2347;
  assign _zz_2347 = ($signed(_zz_2349) + $signed(_zz_26));
  assign _zz_2348 = ({9'd0,data_mid_0_10_real} <<< 9);
  assign _zz_2349 = {{9{_zz_2348[26]}}, _zz_2348};
  assign _zz_2350 = fixTo_34_dout;
  assign _zz_2351 = _zz_2352[35 : 0];
  assign _zz_2352 = _zz_2353;
  assign _zz_2353 = ($signed(_zz_2354) >>> _zz_30);
  assign _zz_2354 = _zz_2355;
  assign _zz_2355 = ($signed(_zz_2357) + $signed(_zz_27));
  assign _zz_2356 = ({9'd0,data_mid_0_10_imag} <<< 9);
  assign _zz_2357 = {{9{_zz_2356[26]}}, _zz_2356};
  assign _zz_2358 = fixTo_35_dout;
  assign _zz_2359 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2360 = ($signed(_zz_33) - $signed(_zz_2361));
  assign _zz_2361 = ($signed(_zz_2362) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2362 = ($signed(data_mid_0_13_real) + $signed(data_mid_0_13_imag));
  assign _zz_2363 = fixTo_36_dout;
  assign _zz_2364 = ($signed(_zz_33) + $signed(_zz_2365));
  assign _zz_2365 = ($signed(_zz_2366) * $signed(twiddle_factor_table_0_real));
  assign _zz_2366 = ($signed(data_mid_0_13_imag) - $signed(data_mid_0_13_real));
  assign _zz_2367 = fixTo_37_dout;
  assign _zz_2368 = _zz_2369[35 : 0];
  assign _zz_2369 = _zz_2370;
  assign _zz_2370 = ($signed(_zz_2371) >>> _zz_34);
  assign _zz_2371 = _zz_2372;
  assign _zz_2372 = ($signed(_zz_2374) - $signed(_zz_31));
  assign _zz_2373 = ({9'd0,data_mid_0_12_real} <<< 9);
  assign _zz_2374 = {{9{_zz_2373[26]}}, _zz_2373};
  assign _zz_2375 = fixTo_38_dout;
  assign _zz_2376 = _zz_2377[35 : 0];
  assign _zz_2377 = _zz_2378;
  assign _zz_2378 = ($signed(_zz_2379) >>> _zz_34);
  assign _zz_2379 = _zz_2380;
  assign _zz_2380 = ($signed(_zz_2382) - $signed(_zz_32));
  assign _zz_2381 = ({9'd0,data_mid_0_12_imag} <<< 9);
  assign _zz_2382 = {{9{_zz_2381[26]}}, _zz_2381};
  assign _zz_2383 = fixTo_39_dout;
  assign _zz_2384 = _zz_2385[35 : 0];
  assign _zz_2385 = _zz_2386;
  assign _zz_2386 = ($signed(_zz_2387) >>> _zz_35);
  assign _zz_2387 = _zz_2388;
  assign _zz_2388 = ($signed(_zz_2390) + $signed(_zz_31));
  assign _zz_2389 = ({9'd0,data_mid_0_12_real} <<< 9);
  assign _zz_2390 = {{9{_zz_2389[26]}}, _zz_2389};
  assign _zz_2391 = fixTo_40_dout;
  assign _zz_2392 = _zz_2393[35 : 0];
  assign _zz_2393 = _zz_2394;
  assign _zz_2394 = ($signed(_zz_2395) >>> _zz_35);
  assign _zz_2395 = _zz_2396;
  assign _zz_2396 = ($signed(_zz_2398) + $signed(_zz_32));
  assign _zz_2397 = ({9'd0,data_mid_0_12_imag} <<< 9);
  assign _zz_2398 = {{9{_zz_2397[26]}}, _zz_2397};
  assign _zz_2399 = fixTo_41_dout;
  assign _zz_2400 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2401 = ($signed(_zz_38) - $signed(_zz_2402));
  assign _zz_2402 = ($signed(_zz_2403) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2403 = ($signed(data_mid_0_15_real) + $signed(data_mid_0_15_imag));
  assign _zz_2404 = fixTo_42_dout;
  assign _zz_2405 = ($signed(_zz_38) + $signed(_zz_2406));
  assign _zz_2406 = ($signed(_zz_2407) * $signed(twiddle_factor_table_0_real));
  assign _zz_2407 = ($signed(data_mid_0_15_imag) - $signed(data_mid_0_15_real));
  assign _zz_2408 = fixTo_43_dout;
  assign _zz_2409 = _zz_2410[35 : 0];
  assign _zz_2410 = _zz_2411;
  assign _zz_2411 = ($signed(_zz_2412) >>> _zz_39);
  assign _zz_2412 = _zz_2413;
  assign _zz_2413 = ($signed(_zz_2415) - $signed(_zz_36));
  assign _zz_2414 = ({9'd0,data_mid_0_14_real} <<< 9);
  assign _zz_2415 = {{9{_zz_2414[26]}}, _zz_2414};
  assign _zz_2416 = fixTo_44_dout;
  assign _zz_2417 = _zz_2418[35 : 0];
  assign _zz_2418 = _zz_2419;
  assign _zz_2419 = ($signed(_zz_2420) >>> _zz_39);
  assign _zz_2420 = _zz_2421;
  assign _zz_2421 = ($signed(_zz_2423) - $signed(_zz_37));
  assign _zz_2422 = ({9'd0,data_mid_0_14_imag} <<< 9);
  assign _zz_2423 = {{9{_zz_2422[26]}}, _zz_2422};
  assign _zz_2424 = fixTo_45_dout;
  assign _zz_2425 = _zz_2426[35 : 0];
  assign _zz_2426 = _zz_2427;
  assign _zz_2427 = ($signed(_zz_2428) >>> _zz_40);
  assign _zz_2428 = _zz_2429;
  assign _zz_2429 = ($signed(_zz_2431) + $signed(_zz_36));
  assign _zz_2430 = ({9'd0,data_mid_0_14_real} <<< 9);
  assign _zz_2431 = {{9{_zz_2430[26]}}, _zz_2430};
  assign _zz_2432 = fixTo_46_dout;
  assign _zz_2433 = _zz_2434[35 : 0];
  assign _zz_2434 = _zz_2435;
  assign _zz_2435 = ($signed(_zz_2436) >>> _zz_40);
  assign _zz_2436 = _zz_2437;
  assign _zz_2437 = ($signed(_zz_2439) + $signed(_zz_37));
  assign _zz_2438 = ({9'd0,data_mid_0_14_imag} <<< 9);
  assign _zz_2439 = {{9{_zz_2438[26]}}, _zz_2438};
  assign _zz_2440 = fixTo_47_dout;
  assign _zz_2441 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2442 = ($signed(_zz_43) - $signed(_zz_2443));
  assign _zz_2443 = ($signed(_zz_2444) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2444 = ($signed(data_mid_0_17_real) + $signed(data_mid_0_17_imag));
  assign _zz_2445 = fixTo_48_dout;
  assign _zz_2446 = ($signed(_zz_43) + $signed(_zz_2447));
  assign _zz_2447 = ($signed(_zz_2448) * $signed(twiddle_factor_table_0_real));
  assign _zz_2448 = ($signed(data_mid_0_17_imag) - $signed(data_mid_0_17_real));
  assign _zz_2449 = fixTo_49_dout;
  assign _zz_2450 = _zz_2451[35 : 0];
  assign _zz_2451 = _zz_2452;
  assign _zz_2452 = ($signed(_zz_2453) >>> _zz_44);
  assign _zz_2453 = _zz_2454;
  assign _zz_2454 = ($signed(_zz_2456) - $signed(_zz_41));
  assign _zz_2455 = ({9'd0,data_mid_0_16_real} <<< 9);
  assign _zz_2456 = {{9{_zz_2455[26]}}, _zz_2455};
  assign _zz_2457 = fixTo_50_dout;
  assign _zz_2458 = _zz_2459[35 : 0];
  assign _zz_2459 = _zz_2460;
  assign _zz_2460 = ($signed(_zz_2461) >>> _zz_44);
  assign _zz_2461 = _zz_2462;
  assign _zz_2462 = ($signed(_zz_2464) - $signed(_zz_42));
  assign _zz_2463 = ({9'd0,data_mid_0_16_imag} <<< 9);
  assign _zz_2464 = {{9{_zz_2463[26]}}, _zz_2463};
  assign _zz_2465 = fixTo_51_dout;
  assign _zz_2466 = _zz_2467[35 : 0];
  assign _zz_2467 = _zz_2468;
  assign _zz_2468 = ($signed(_zz_2469) >>> _zz_45);
  assign _zz_2469 = _zz_2470;
  assign _zz_2470 = ($signed(_zz_2472) + $signed(_zz_41));
  assign _zz_2471 = ({9'd0,data_mid_0_16_real} <<< 9);
  assign _zz_2472 = {{9{_zz_2471[26]}}, _zz_2471};
  assign _zz_2473 = fixTo_52_dout;
  assign _zz_2474 = _zz_2475[35 : 0];
  assign _zz_2475 = _zz_2476;
  assign _zz_2476 = ($signed(_zz_2477) >>> _zz_45);
  assign _zz_2477 = _zz_2478;
  assign _zz_2478 = ($signed(_zz_2480) + $signed(_zz_42));
  assign _zz_2479 = ({9'd0,data_mid_0_16_imag} <<< 9);
  assign _zz_2480 = {{9{_zz_2479[26]}}, _zz_2479};
  assign _zz_2481 = fixTo_53_dout;
  assign _zz_2482 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2483 = ($signed(_zz_48) - $signed(_zz_2484));
  assign _zz_2484 = ($signed(_zz_2485) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2485 = ($signed(data_mid_0_19_real) + $signed(data_mid_0_19_imag));
  assign _zz_2486 = fixTo_54_dout;
  assign _zz_2487 = ($signed(_zz_48) + $signed(_zz_2488));
  assign _zz_2488 = ($signed(_zz_2489) * $signed(twiddle_factor_table_0_real));
  assign _zz_2489 = ($signed(data_mid_0_19_imag) - $signed(data_mid_0_19_real));
  assign _zz_2490 = fixTo_55_dout;
  assign _zz_2491 = _zz_2492[35 : 0];
  assign _zz_2492 = _zz_2493;
  assign _zz_2493 = ($signed(_zz_2494) >>> _zz_49);
  assign _zz_2494 = _zz_2495;
  assign _zz_2495 = ($signed(_zz_2497) - $signed(_zz_46));
  assign _zz_2496 = ({9'd0,data_mid_0_18_real} <<< 9);
  assign _zz_2497 = {{9{_zz_2496[26]}}, _zz_2496};
  assign _zz_2498 = fixTo_56_dout;
  assign _zz_2499 = _zz_2500[35 : 0];
  assign _zz_2500 = _zz_2501;
  assign _zz_2501 = ($signed(_zz_2502) >>> _zz_49);
  assign _zz_2502 = _zz_2503;
  assign _zz_2503 = ($signed(_zz_2505) - $signed(_zz_47));
  assign _zz_2504 = ({9'd0,data_mid_0_18_imag} <<< 9);
  assign _zz_2505 = {{9{_zz_2504[26]}}, _zz_2504};
  assign _zz_2506 = fixTo_57_dout;
  assign _zz_2507 = _zz_2508[35 : 0];
  assign _zz_2508 = _zz_2509;
  assign _zz_2509 = ($signed(_zz_2510) >>> _zz_50);
  assign _zz_2510 = _zz_2511;
  assign _zz_2511 = ($signed(_zz_2513) + $signed(_zz_46));
  assign _zz_2512 = ({9'd0,data_mid_0_18_real} <<< 9);
  assign _zz_2513 = {{9{_zz_2512[26]}}, _zz_2512};
  assign _zz_2514 = fixTo_58_dout;
  assign _zz_2515 = _zz_2516[35 : 0];
  assign _zz_2516 = _zz_2517;
  assign _zz_2517 = ($signed(_zz_2518) >>> _zz_50);
  assign _zz_2518 = _zz_2519;
  assign _zz_2519 = ($signed(_zz_2521) + $signed(_zz_47));
  assign _zz_2520 = ({9'd0,data_mid_0_18_imag} <<< 9);
  assign _zz_2521 = {{9{_zz_2520[26]}}, _zz_2520};
  assign _zz_2522 = fixTo_59_dout;
  assign _zz_2523 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2524 = ($signed(_zz_53) - $signed(_zz_2525));
  assign _zz_2525 = ($signed(_zz_2526) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2526 = ($signed(data_mid_0_21_real) + $signed(data_mid_0_21_imag));
  assign _zz_2527 = fixTo_60_dout;
  assign _zz_2528 = ($signed(_zz_53) + $signed(_zz_2529));
  assign _zz_2529 = ($signed(_zz_2530) * $signed(twiddle_factor_table_0_real));
  assign _zz_2530 = ($signed(data_mid_0_21_imag) - $signed(data_mid_0_21_real));
  assign _zz_2531 = fixTo_61_dout;
  assign _zz_2532 = _zz_2533[35 : 0];
  assign _zz_2533 = _zz_2534;
  assign _zz_2534 = ($signed(_zz_2535) >>> _zz_54);
  assign _zz_2535 = _zz_2536;
  assign _zz_2536 = ($signed(_zz_2538) - $signed(_zz_51));
  assign _zz_2537 = ({9'd0,data_mid_0_20_real} <<< 9);
  assign _zz_2538 = {{9{_zz_2537[26]}}, _zz_2537};
  assign _zz_2539 = fixTo_62_dout;
  assign _zz_2540 = _zz_2541[35 : 0];
  assign _zz_2541 = _zz_2542;
  assign _zz_2542 = ($signed(_zz_2543) >>> _zz_54);
  assign _zz_2543 = _zz_2544;
  assign _zz_2544 = ($signed(_zz_2546) - $signed(_zz_52));
  assign _zz_2545 = ({9'd0,data_mid_0_20_imag} <<< 9);
  assign _zz_2546 = {{9{_zz_2545[26]}}, _zz_2545};
  assign _zz_2547 = fixTo_63_dout;
  assign _zz_2548 = _zz_2549[35 : 0];
  assign _zz_2549 = _zz_2550;
  assign _zz_2550 = ($signed(_zz_2551) >>> _zz_55);
  assign _zz_2551 = _zz_2552;
  assign _zz_2552 = ($signed(_zz_2554) + $signed(_zz_51));
  assign _zz_2553 = ({9'd0,data_mid_0_20_real} <<< 9);
  assign _zz_2554 = {{9{_zz_2553[26]}}, _zz_2553};
  assign _zz_2555 = fixTo_64_dout;
  assign _zz_2556 = _zz_2557[35 : 0];
  assign _zz_2557 = _zz_2558;
  assign _zz_2558 = ($signed(_zz_2559) >>> _zz_55);
  assign _zz_2559 = _zz_2560;
  assign _zz_2560 = ($signed(_zz_2562) + $signed(_zz_52));
  assign _zz_2561 = ({9'd0,data_mid_0_20_imag} <<< 9);
  assign _zz_2562 = {{9{_zz_2561[26]}}, _zz_2561};
  assign _zz_2563 = fixTo_65_dout;
  assign _zz_2564 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2565 = ($signed(_zz_58) - $signed(_zz_2566));
  assign _zz_2566 = ($signed(_zz_2567) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2567 = ($signed(data_mid_0_23_real) + $signed(data_mid_0_23_imag));
  assign _zz_2568 = fixTo_66_dout;
  assign _zz_2569 = ($signed(_zz_58) + $signed(_zz_2570));
  assign _zz_2570 = ($signed(_zz_2571) * $signed(twiddle_factor_table_0_real));
  assign _zz_2571 = ($signed(data_mid_0_23_imag) - $signed(data_mid_0_23_real));
  assign _zz_2572 = fixTo_67_dout;
  assign _zz_2573 = _zz_2574[35 : 0];
  assign _zz_2574 = _zz_2575;
  assign _zz_2575 = ($signed(_zz_2576) >>> _zz_59);
  assign _zz_2576 = _zz_2577;
  assign _zz_2577 = ($signed(_zz_2579) - $signed(_zz_56));
  assign _zz_2578 = ({9'd0,data_mid_0_22_real} <<< 9);
  assign _zz_2579 = {{9{_zz_2578[26]}}, _zz_2578};
  assign _zz_2580 = fixTo_68_dout;
  assign _zz_2581 = _zz_2582[35 : 0];
  assign _zz_2582 = _zz_2583;
  assign _zz_2583 = ($signed(_zz_2584) >>> _zz_59);
  assign _zz_2584 = _zz_2585;
  assign _zz_2585 = ($signed(_zz_2587) - $signed(_zz_57));
  assign _zz_2586 = ({9'd0,data_mid_0_22_imag} <<< 9);
  assign _zz_2587 = {{9{_zz_2586[26]}}, _zz_2586};
  assign _zz_2588 = fixTo_69_dout;
  assign _zz_2589 = _zz_2590[35 : 0];
  assign _zz_2590 = _zz_2591;
  assign _zz_2591 = ($signed(_zz_2592) >>> _zz_60);
  assign _zz_2592 = _zz_2593;
  assign _zz_2593 = ($signed(_zz_2595) + $signed(_zz_56));
  assign _zz_2594 = ({9'd0,data_mid_0_22_real} <<< 9);
  assign _zz_2595 = {{9{_zz_2594[26]}}, _zz_2594};
  assign _zz_2596 = fixTo_70_dout;
  assign _zz_2597 = _zz_2598[35 : 0];
  assign _zz_2598 = _zz_2599;
  assign _zz_2599 = ($signed(_zz_2600) >>> _zz_60);
  assign _zz_2600 = _zz_2601;
  assign _zz_2601 = ($signed(_zz_2603) + $signed(_zz_57));
  assign _zz_2602 = ({9'd0,data_mid_0_22_imag} <<< 9);
  assign _zz_2603 = {{9{_zz_2602[26]}}, _zz_2602};
  assign _zz_2604 = fixTo_71_dout;
  assign _zz_2605 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2606 = ($signed(_zz_63) - $signed(_zz_2607));
  assign _zz_2607 = ($signed(_zz_2608) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2608 = ($signed(data_mid_0_25_real) + $signed(data_mid_0_25_imag));
  assign _zz_2609 = fixTo_72_dout;
  assign _zz_2610 = ($signed(_zz_63) + $signed(_zz_2611));
  assign _zz_2611 = ($signed(_zz_2612) * $signed(twiddle_factor_table_0_real));
  assign _zz_2612 = ($signed(data_mid_0_25_imag) - $signed(data_mid_0_25_real));
  assign _zz_2613 = fixTo_73_dout;
  assign _zz_2614 = _zz_2615[35 : 0];
  assign _zz_2615 = _zz_2616;
  assign _zz_2616 = ($signed(_zz_2617) >>> _zz_64);
  assign _zz_2617 = _zz_2618;
  assign _zz_2618 = ($signed(_zz_2620) - $signed(_zz_61));
  assign _zz_2619 = ({9'd0,data_mid_0_24_real} <<< 9);
  assign _zz_2620 = {{9{_zz_2619[26]}}, _zz_2619};
  assign _zz_2621 = fixTo_74_dout;
  assign _zz_2622 = _zz_2623[35 : 0];
  assign _zz_2623 = _zz_2624;
  assign _zz_2624 = ($signed(_zz_2625) >>> _zz_64);
  assign _zz_2625 = _zz_2626;
  assign _zz_2626 = ($signed(_zz_2628) - $signed(_zz_62));
  assign _zz_2627 = ({9'd0,data_mid_0_24_imag} <<< 9);
  assign _zz_2628 = {{9{_zz_2627[26]}}, _zz_2627};
  assign _zz_2629 = fixTo_75_dout;
  assign _zz_2630 = _zz_2631[35 : 0];
  assign _zz_2631 = _zz_2632;
  assign _zz_2632 = ($signed(_zz_2633) >>> _zz_65);
  assign _zz_2633 = _zz_2634;
  assign _zz_2634 = ($signed(_zz_2636) + $signed(_zz_61));
  assign _zz_2635 = ({9'd0,data_mid_0_24_real} <<< 9);
  assign _zz_2636 = {{9{_zz_2635[26]}}, _zz_2635};
  assign _zz_2637 = fixTo_76_dout;
  assign _zz_2638 = _zz_2639[35 : 0];
  assign _zz_2639 = _zz_2640;
  assign _zz_2640 = ($signed(_zz_2641) >>> _zz_65);
  assign _zz_2641 = _zz_2642;
  assign _zz_2642 = ($signed(_zz_2644) + $signed(_zz_62));
  assign _zz_2643 = ({9'd0,data_mid_0_24_imag} <<< 9);
  assign _zz_2644 = {{9{_zz_2643[26]}}, _zz_2643};
  assign _zz_2645 = fixTo_77_dout;
  assign _zz_2646 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2647 = ($signed(_zz_68) - $signed(_zz_2648));
  assign _zz_2648 = ($signed(_zz_2649) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2649 = ($signed(data_mid_0_27_real) + $signed(data_mid_0_27_imag));
  assign _zz_2650 = fixTo_78_dout;
  assign _zz_2651 = ($signed(_zz_68) + $signed(_zz_2652));
  assign _zz_2652 = ($signed(_zz_2653) * $signed(twiddle_factor_table_0_real));
  assign _zz_2653 = ($signed(data_mid_0_27_imag) - $signed(data_mid_0_27_real));
  assign _zz_2654 = fixTo_79_dout;
  assign _zz_2655 = _zz_2656[35 : 0];
  assign _zz_2656 = _zz_2657;
  assign _zz_2657 = ($signed(_zz_2658) >>> _zz_69);
  assign _zz_2658 = _zz_2659;
  assign _zz_2659 = ($signed(_zz_2661) - $signed(_zz_66));
  assign _zz_2660 = ({9'd0,data_mid_0_26_real} <<< 9);
  assign _zz_2661 = {{9{_zz_2660[26]}}, _zz_2660};
  assign _zz_2662 = fixTo_80_dout;
  assign _zz_2663 = _zz_2664[35 : 0];
  assign _zz_2664 = _zz_2665;
  assign _zz_2665 = ($signed(_zz_2666) >>> _zz_69);
  assign _zz_2666 = _zz_2667;
  assign _zz_2667 = ($signed(_zz_2669) - $signed(_zz_67));
  assign _zz_2668 = ({9'd0,data_mid_0_26_imag} <<< 9);
  assign _zz_2669 = {{9{_zz_2668[26]}}, _zz_2668};
  assign _zz_2670 = fixTo_81_dout;
  assign _zz_2671 = _zz_2672[35 : 0];
  assign _zz_2672 = _zz_2673;
  assign _zz_2673 = ($signed(_zz_2674) >>> _zz_70);
  assign _zz_2674 = _zz_2675;
  assign _zz_2675 = ($signed(_zz_2677) + $signed(_zz_66));
  assign _zz_2676 = ({9'd0,data_mid_0_26_real} <<< 9);
  assign _zz_2677 = {{9{_zz_2676[26]}}, _zz_2676};
  assign _zz_2678 = fixTo_82_dout;
  assign _zz_2679 = _zz_2680[35 : 0];
  assign _zz_2680 = _zz_2681;
  assign _zz_2681 = ($signed(_zz_2682) >>> _zz_70);
  assign _zz_2682 = _zz_2683;
  assign _zz_2683 = ($signed(_zz_2685) + $signed(_zz_67));
  assign _zz_2684 = ({9'd0,data_mid_0_26_imag} <<< 9);
  assign _zz_2685 = {{9{_zz_2684[26]}}, _zz_2684};
  assign _zz_2686 = fixTo_83_dout;
  assign _zz_2687 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2688 = ($signed(_zz_73) - $signed(_zz_2689));
  assign _zz_2689 = ($signed(_zz_2690) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2690 = ($signed(data_mid_0_29_real) + $signed(data_mid_0_29_imag));
  assign _zz_2691 = fixTo_84_dout;
  assign _zz_2692 = ($signed(_zz_73) + $signed(_zz_2693));
  assign _zz_2693 = ($signed(_zz_2694) * $signed(twiddle_factor_table_0_real));
  assign _zz_2694 = ($signed(data_mid_0_29_imag) - $signed(data_mid_0_29_real));
  assign _zz_2695 = fixTo_85_dout;
  assign _zz_2696 = _zz_2697[35 : 0];
  assign _zz_2697 = _zz_2698;
  assign _zz_2698 = ($signed(_zz_2699) >>> _zz_74);
  assign _zz_2699 = _zz_2700;
  assign _zz_2700 = ($signed(_zz_2702) - $signed(_zz_71));
  assign _zz_2701 = ({9'd0,data_mid_0_28_real} <<< 9);
  assign _zz_2702 = {{9{_zz_2701[26]}}, _zz_2701};
  assign _zz_2703 = fixTo_86_dout;
  assign _zz_2704 = _zz_2705[35 : 0];
  assign _zz_2705 = _zz_2706;
  assign _zz_2706 = ($signed(_zz_2707) >>> _zz_74);
  assign _zz_2707 = _zz_2708;
  assign _zz_2708 = ($signed(_zz_2710) - $signed(_zz_72));
  assign _zz_2709 = ({9'd0,data_mid_0_28_imag} <<< 9);
  assign _zz_2710 = {{9{_zz_2709[26]}}, _zz_2709};
  assign _zz_2711 = fixTo_87_dout;
  assign _zz_2712 = _zz_2713[35 : 0];
  assign _zz_2713 = _zz_2714;
  assign _zz_2714 = ($signed(_zz_2715) >>> _zz_75);
  assign _zz_2715 = _zz_2716;
  assign _zz_2716 = ($signed(_zz_2718) + $signed(_zz_71));
  assign _zz_2717 = ({9'd0,data_mid_0_28_real} <<< 9);
  assign _zz_2718 = {{9{_zz_2717[26]}}, _zz_2717};
  assign _zz_2719 = fixTo_88_dout;
  assign _zz_2720 = _zz_2721[35 : 0];
  assign _zz_2721 = _zz_2722;
  assign _zz_2722 = ($signed(_zz_2723) >>> _zz_75);
  assign _zz_2723 = _zz_2724;
  assign _zz_2724 = ($signed(_zz_2726) + $signed(_zz_72));
  assign _zz_2725 = ({9'd0,data_mid_0_28_imag} <<< 9);
  assign _zz_2726 = {{9{_zz_2725[26]}}, _zz_2725};
  assign _zz_2727 = fixTo_89_dout;
  assign _zz_2728 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2729 = ($signed(_zz_78) - $signed(_zz_2730));
  assign _zz_2730 = ($signed(_zz_2731) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2731 = ($signed(data_mid_0_31_real) + $signed(data_mid_0_31_imag));
  assign _zz_2732 = fixTo_90_dout;
  assign _zz_2733 = ($signed(_zz_78) + $signed(_zz_2734));
  assign _zz_2734 = ($signed(_zz_2735) * $signed(twiddle_factor_table_0_real));
  assign _zz_2735 = ($signed(data_mid_0_31_imag) - $signed(data_mid_0_31_real));
  assign _zz_2736 = fixTo_91_dout;
  assign _zz_2737 = _zz_2738[35 : 0];
  assign _zz_2738 = _zz_2739;
  assign _zz_2739 = ($signed(_zz_2740) >>> _zz_79);
  assign _zz_2740 = _zz_2741;
  assign _zz_2741 = ($signed(_zz_2743) - $signed(_zz_76));
  assign _zz_2742 = ({9'd0,data_mid_0_30_real} <<< 9);
  assign _zz_2743 = {{9{_zz_2742[26]}}, _zz_2742};
  assign _zz_2744 = fixTo_92_dout;
  assign _zz_2745 = _zz_2746[35 : 0];
  assign _zz_2746 = _zz_2747;
  assign _zz_2747 = ($signed(_zz_2748) >>> _zz_79);
  assign _zz_2748 = _zz_2749;
  assign _zz_2749 = ($signed(_zz_2751) - $signed(_zz_77));
  assign _zz_2750 = ({9'd0,data_mid_0_30_imag} <<< 9);
  assign _zz_2751 = {{9{_zz_2750[26]}}, _zz_2750};
  assign _zz_2752 = fixTo_93_dout;
  assign _zz_2753 = _zz_2754[35 : 0];
  assign _zz_2754 = _zz_2755;
  assign _zz_2755 = ($signed(_zz_2756) >>> _zz_80);
  assign _zz_2756 = _zz_2757;
  assign _zz_2757 = ($signed(_zz_2759) + $signed(_zz_76));
  assign _zz_2758 = ({9'd0,data_mid_0_30_real} <<< 9);
  assign _zz_2759 = {{9{_zz_2758[26]}}, _zz_2758};
  assign _zz_2760 = fixTo_94_dout;
  assign _zz_2761 = _zz_2762[35 : 0];
  assign _zz_2762 = _zz_2763;
  assign _zz_2763 = ($signed(_zz_2764) >>> _zz_80);
  assign _zz_2764 = _zz_2765;
  assign _zz_2765 = ($signed(_zz_2767) + $signed(_zz_77));
  assign _zz_2766 = ({9'd0,data_mid_0_30_imag} <<< 9);
  assign _zz_2767 = {{9{_zz_2766[26]}}, _zz_2766};
  assign _zz_2768 = fixTo_95_dout;
  assign _zz_2769 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2770 = ($signed(_zz_83) - $signed(_zz_2771));
  assign _zz_2771 = ($signed(_zz_2772) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2772 = ($signed(data_mid_0_33_real) + $signed(data_mid_0_33_imag));
  assign _zz_2773 = fixTo_96_dout;
  assign _zz_2774 = ($signed(_zz_83) + $signed(_zz_2775));
  assign _zz_2775 = ($signed(_zz_2776) * $signed(twiddle_factor_table_0_real));
  assign _zz_2776 = ($signed(data_mid_0_33_imag) - $signed(data_mid_0_33_real));
  assign _zz_2777 = fixTo_97_dout;
  assign _zz_2778 = _zz_2779[35 : 0];
  assign _zz_2779 = _zz_2780;
  assign _zz_2780 = ($signed(_zz_2781) >>> _zz_84);
  assign _zz_2781 = _zz_2782;
  assign _zz_2782 = ($signed(_zz_2784) - $signed(_zz_81));
  assign _zz_2783 = ({9'd0,data_mid_0_32_real} <<< 9);
  assign _zz_2784 = {{9{_zz_2783[26]}}, _zz_2783};
  assign _zz_2785 = fixTo_98_dout;
  assign _zz_2786 = _zz_2787[35 : 0];
  assign _zz_2787 = _zz_2788;
  assign _zz_2788 = ($signed(_zz_2789) >>> _zz_84);
  assign _zz_2789 = _zz_2790;
  assign _zz_2790 = ($signed(_zz_2792) - $signed(_zz_82));
  assign _zz_2791 = ({9'd0,data_mid_0_32_imag} <<< 9);
  assign _zz_2792 = {{9{_zz_2791[26]}}, _zz_2791};
  assign _zz_2793 = fixTo_99_dout;
  assign _zz_2794 = _zz_2795[35 : 0];
  assign _zz_2795 = _zz_2796;
  assign _zz_2796 = ($signed(_zz_2797) >>> _zz_85);
  assign _zz_2797 = _zz_2798;
  assign _zz_2798 = ($signed(_zz_2800) + $signed(_zz_81));
  assign _zz_2799 = ({9'd0,data_mid_0_32_real} <<< 9);
  assign _zz_2800 = {{9{_zz_2799[26]}}, _zz_2799};
  assign _zz_2801 = fixTo_100_dout;
  assign _zz_2802 = _zz_2803[35 : 0];
  assign _zz_2803 = _zz_2804;
  assign _zz_2804 = ($signed(_zz_2805) >>> _zz_85);
  assign _zz_2805 = _zz_2806;
  assign _zz_2806 = ($signed(_zz_2808) + $signed(_zz_82));
  assign _zz_2807 = ({9'd0,data_mid_0_32_imag} <<< 9);
  assign _zz_2808 = {{9{_zz_2807[26]}}, _zz_2807};
  assign _zz_2809 = fixTo_101_dout;
  assign _zz_2810 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2811 = ($signed(_zz_88) - $signed(_zz_2812));
  assign _zz_2812 = ($signed(_zz_2813) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2813 = ($signed(data_mid_0_35_real) + $signed(data_mid_0_35_imag));
  assign _zz_2814 = fixTo_102_dout;
  assign _zz_2815 = ($signed(_zz_88) + $signed(_zz_2816));
  assign _zz_2816 = ($signed(_zz_2817) * $signed(twiddle_factor_table_0_real));
  assign _zz_2817 = ($signed(data_mid_0_35_imag) - $signed(data_mid_0_35_real));
  assign _zz_2818 = fixTo_103_dout;
  assign _zz_2819 = _zz_2820[35 : 0];
  assign _zz_2820 = _zz_2821;
  assign _zz_2821 = ($signed(_zz_2822) >>> _zz_89);
  assign _zz_2822 = _zz_2823;
  assign _zz_2823 = ($signed(_zz_2825) - $signed(_zz_86));
  assign _zz_2824 = ({9'd0,data_mid_0_34_real} <<< 9);
  assign _zz_2825 = {{9{_zz_2824[26]}}, _zz_2824};
  assign _zz_2826 = fixTo_104_dout;
  assign _zz_2827 = _zz_2828[35 : 0];
  assign _zz_2828 = _zz_2829;
  assign _zz_2829 = ($signed(_zz_2830) >>> _zz_89);
  assign _zz_2830 = _zz_2831;
  assign _zz_2831 = ($signed(_zz_2833) - $signed(_zz_87));
  assign _zz_2832 = ({9'd0,data_mid_0_34_imag} <<< 9);
  assign _zz_2833 = {{9{_zz_2832[26]}}, _zz_2832};
  assign _zz_2834 = fixTo_105_dout;
  assign _zz_2835 = _zz_2836[35 : 0];
  assign _zz_2836 = _zz_2837;
  assign _zz_2837 = ($signed(_zz_2838) >>> _zz_90);
  assign _zz_2838 = _zz_2839;
  assign _zz_2839 = ($signed(_zz_2841) + $signed(_zz_86));
  assign _zz_2840 = ({9'd0,data_mid_0_34_real} <<< 9);
  assign _zz_2841 = {{9{_zz_2840[26]}}, _zz_2840};
  assign _zz_2842 = fixTo_106_dout;
  assign _zz_2843 = _zz_2844[35 : 0];
  assign _zz_2844 = _zz_2845;
  assign _zz_2845 = ($signed(_zz_2846) >>> _zz_90);
  assign _zz_2846 = _zz_2847;
  assign _zz_2847 = ($signed(_zz_2849) + $signed(_zz_87));
  assign _zz_2848 = ({9'd0,data_mid_0_34_imag} <<< 9);
  assign _zz_2849 = {{9{_zz_2848[26]}}, _zz_2848};
  assign _zz_2850 = fixTo_107_dout;
  assign _zz_2851 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2852 = ($signed(_zz_93) - $signed(_zz_2853));
  assign _zz_2853 = ($signed(_zz_2854) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2854 = ($signed(data_mid_0_37_real) + $signed(data_mid_0_37_imag));
  assign _zz_2855 = fixTo_108_dout;
  assign _zz_2856 = ($signed(_zz_93) + $signed(_zz_2857));
  assign _zz_2857 = ($signed(_zz_2858) * $signed(twiddle_factor_table_0_real));
  assign _zz_2858 = ($signed(data_mid_0_37_imag) - $signed(data_mid_0_37_real));
  assign _zz_2859 = fixTo_109_dout;
  assign _zz_2860 = _zz_2861[35 : 0];
  assign _zz_2861 = _zz_2862;
  assign _zz_2862 = ($signed(_zz_2863) >>> _zz_94);
  assign _zz_2863 = _zz_2864;
  assign _zz_2864 = ($signed(_zz_2866) - $signed(_zz_91));
  assign _zz_2865 = ({9'd0,data_mid_0_36_real} <<< 9);
  assign _zz_2866 = {{9{_zz_2865[26]}}, _zz_2865};
  assign _zz_2867 = fixTo_110_dout;
  assign _zz_2868 = _zz_2869[35 : 0];
  assign _zz_2869 = _zz_2870;
  assign _zz_2870 = ($signed(_zz_2871) >>> _zz_94);
  assign _zz_2871 = _zz_2872;
  assign _zz_2872 = ($signed(_zz_2874) - $signed(_zz_92));
  assign _zz_2873 = ({9'd0,data_mid_0_36_imag} <<< 9);
  assign _zz_2874 = {{9{_zz_2873[26]}}, _zz_2873};
  assign _zz_2875 = fixTo_111_dout;
  assign _zz_2876 = _zz_2877[35 : 0];
  assign _zz_2877 = _zz_2878;
  assign _zz_2878 = ($signed(_zz_2879) >>> _zz_95);
  assign _zz_2879 = _zz_2880;
  assign _zz_2880 = ($signed(_zz_2882) + $signed(_zz_91));
  assign _zz_2881 = ({9'd0,data_mid_0_36_real} <<< 9);
  assign _zz_2882 = {{9{_zz_2881[26]}}, _zz_2881};
  assign _zz_2883 = fixTo_112_dout;
  assign _zz_2884 = _zz_2885[35 : 0];
  assign _zz_2885 = _zz_2886;
  assign _zz_2886 = ($signed(_zz_2887) >>> _zz_95);
  assign _zz_2887 = _zz_2888;
  assign _zz_2888 = ($signed(_zz_2890) + $signed(_zz_92));
  assign _zz_2889 = ({9'd0,data_mid_0_36_imag} <<< 9);
  assign _zz_2890 = {{9{_zz_2889[26]}}, _zz_2889};
  assign _zz_2891 = fixTo_113_dout;
  assign _zz_2892 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2893 = ($signed(_zz_98) - $signed(_zz_2894));
  assign _zz_2894 = ($signed(_zz_2895) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2895 = ($signed(data_mid_0_39_real) + $signed(data_mid_0_39_imag));
  assign _zz_2896 = fixTo_114_dout;
  assign _zz_2897 = ($signed(_zz_98) + $signed(_zz_2898));
  assign _zz_2898 = ($signed(_zz_2899) * $signed(twiddle_factor_table_0_real));
  assign _zz_2899 = ($signed(data_mid_0_39_imag) - $signed(data_mid_0_39_real));
  assign _zz_2900 = fixTo_115_dout;
  assign _zz_2901 = _zz_2902[35 : 0];
  assign _zz_2902 = _zz_2903;
  assign _zz_2903 = ($signed(_zz_2904) >>> _zz_99);
  assign _zz_2904 = _zz_2905;
  assign _zz_2905 = ($signed(_zz_2907) - $signed(_zz_96));
  assign _zz_2906 = ({9'd0,data_mid_0_38_real} <<< 9);
  assign _zz_2907 = {{9{_zz_2906[26]}}, _zz_2906};
  assign _zz_2908 = fixTo_116_dout;
  assign _zz_2909 = _zz_2910[35 : 0];
  assign _zz_2910 = _zz_2911;
  assign _zz_2911 = ($signed(_zz_2912) >>> _zz_99);
  assign _zz_2912 = _zz_2913;
  assign _zz_2913 = ($signed(_zz_2915) - $signed(_zz_97));
  assign _zz_2914 = ({9'd0,data_mid_0_38_imag} <<< 9);
  assign _zz_2915 = {{9{_zz_2914[26]}}, _zz_2914};
  assign _zz_2916 = fixTo_117_dout;
  assign _zz_2917 = _zz_2918[35 : 0];
  assign _zz_2918 = _zz_2919;
  assign _zz_2919 = ($signed(_zz_2920) >>> _zz_100);
  assign _zz_2920 = _zz_2921;
  assign _zz_2921 = ($signed(_zz_2923) + $signed(_zz_96));
  assign _zz_2922 = ({9'd0,data_mid_0_38_real} <<< 9);
  assign _zz_2923 = {{9{_zz_2922[26]}}, _zz_2922};
  assign _zz_2924 = fixTo_118_dout;
  assign _zz_2925 = _zz_2926[35 : 0];
  assign _zz_2926 = _zz_2927;
  assign _zz_2927 = ($signed(_zz_2928) >>> _zz_100);
  assign _zz_2928 = _zz_2929;
  assign _zz_2929 = ($signed(_zz_2931) + $signed(_zz_97));
  assign _zz_2930 = ({9'd0,data_mid_0_38_imag} <<< 9);
  assign _zz_2931 = {{9{_zz_2930[26]}}, _zz_2930};
  assign _zz_2932 = fixTo_119_dout;
  assign _zz_2933 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2934 = ($signed(_zz_103) - $signed(_zz_2935));
  assign _zz_2935 = ($signed(_zz_2936) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2936 = ($signed(data_mid_0_41_real) + $signed(data_mid_0_41_imag));
  assign _zz_2937 = fixTo_120_dout;
  assign _zz_2938 = ($signed(_zz_103) + $signed(_zz_2939));
  assign _zz_2939 = ($signed(_zz_2940) * $signed(twiddle_factor_table_0_real));
  assign _zz_2940 = ($signed(data_mid_0_41_imag) - $signed(data_mid_0_41_real));
  assign _zz_2941 = fixTo_121_dout;
  assign _zz_2942 = _zz_2943[35 : 0];
  assign _zz_2943 = _zz_2944;
  assign _zz_2944 = ($signed(_zz_2945) >>> _zz_104);
  assign _zz_2945 = _zz_2946;
  assign _zz_2946 = ($signed(_zz_2948) - $signed(_zz_101));
  assign _zz_2947 = ({9'd0,data_mid_0_40_real} <<< 9);
  assign _zz_2948 = {{9{_zz_2947[26]}}, _zz_2947};
  assign _zz_2949 = fixTo_122_dout;
  assign _zz_2950 = _zz_2951[35 : 0];
  assign _zz_2951 = _zz_2952;
  assign _zz_2952 = ($signed(_zz_2953) >>> _zz_104);
  assign _zz_2953 = _zz_2954;
  assign _zz_2954 = ($signed(_zz_2956) - $signed(_zz_102));
  assign _zz_2955 = ({9'd0,data_mid_0_40_imag} <<< 9);
  assign _zz_2956 = {{9{_zz_2955[26]}}, _zz_2955};
  assign _zz_2957 = fixTo_123_dout;
  assign _zz_2958 = _zz_2959[35 : 0];
  assign _zz_2959 = _zz_2960;
  assign _zz_2960 = ($signed(_zz_2961) >>> _zz_105);
  assign _zz_2961 = _zz_2962;
  assign _zz_2962 = ($signed(_zz_2964) + $signed(_zz_101));
  assign _zz_2963 = ({9'd0,data_mid_0_40_real} <<< 9);
  assign _zz_2964 = {{9{_zz_2963[26]}}, _zz_2963};
  assign _zz_2965 = fixTo_124_dout;
  assign _zz_2966 = _zz_2967[35 : 0];
  assign _zz_2967 = _zz_2968;
  assign _zz_2968 = ($signed(_zz_2969) >>> _zz_105);
  assign _zz_2969 = _zz_2970;
  assign _zz_2970 = ($signed(_zz_2972) + $signed(_zz_102));
  assign _zz_2971 = ({9'd0,data_mid_0_40_imag} <<< 9);
  assign _zz_2972 = {{9{_zz_2971[26]}}, _zz_2971};
  assign _zz_2973 = fixTo_125_dout;
  assign _zz_2974 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2975 = ($signed(_zz_108) - $signed(_zz_2976));
  assign _zz_2976 = ($signed(_zz_2977) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2977 = ($signed(data_mid_0_43_real) + $signed(data_mid_0_43_imag));
  assign _zz_2978 = fixTo_126_dout;
  assign _zz_2979 = ($signed(_zz_108) + $signed(_zz_2980));
  assign _zz_2980 = ($signed(_zz_2981) * $signed(twiddle_factor_table_0_real));
  assign _zz_2981 = ($signed(data_mid_0_43_imag) - $signed(data_mid_0_43_real));
  assign _zz_2982 = fixTo_127_dout;
  assign _zz_2983 = _zz_2984[35 : 0];
  assign _zz_2984 = _zz_2985;
  assign _zz_2985 = ($signed(_zz_2986) >>> _zz_109);
  assign _zz_2986 = _zz_2987;
  assign _zz_2987 = ($signed(_zz_2989) - $signed(_zz_106));
  assign _zz_2988 = ({9'd0,data_mid_0_42_real} <<< 9);
  assign _zz_2989 = {{9{_zz_2988[26]}}, _zz_2988};
  assign _zz_2990 = fixTo_128_dout;
  assign _zz_2991 = _zz_2992[35 : 0];
  assign _zz_2992 = _zz_2993;
  assign _zz_2993 = ($signed(_zz_2994) >>> _zz_109);
  assign _zz_2994 = _zz_2995;
  assign _zz_2995 = ($signed(_zz_2997) - $signed(_zz_107));
  assign _zz_2996 = ({9'd0,data_mid_0_42_imag} <<< 9);
  assign _zz_2997 = {{9{_zz_2996[26]}}, _zz_2996};
  assign _zz_2998 = fixTo_129_dout;
  assign _zz_2999 = _zz_3000[35 : 0];
  assign _zz_3000 = _zz_3001;
  assign _zz_3001 = ($signed(_zz_3002) >>> _zz_110);
  assign _zz_3002 = _zz_3003;
  assign _zz_3003 = ($signed(_zz_3005) + $signed(_zz_106));
  assign _zz_3004 = ({9'd0,data_mid_0_42_real} <<< 9);
  assign _zz_3005 = {{9{_zz_3004[26]}}, _zz_3004};
  assign _zz_3006 = fixTo_130_dout;
  assign _zz_3007 = _zz_3008[35 : 0];
  assign _zz_3008 = _zz_3009;
  assign _zz_3009 = ($signed(_zz_3010) >>> _zz_110);
  assign _zz_3010 = _zz_3011;
  assign _zz_3011 = ($signed(_zz_3013) + $signed(_zz_107));
  assign _zz_3012 = ({9'd0,data_mid_0_42_imag} <<< 9);
  assign _zz_3013 = {{9{_zz_3012[26]}}, _zz_3012};
  assign _zz_3014 = fixTo_131_dout;
  assign _zz_3015 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_3016 = ($signed(_zz_113) - $signed(_zz_3017));
  assign _zz_3017 = ($signed(_zz_3018) * $signed(twiddle_factor_table_0_imag));
  assign _zz_3018 = ($signed(data_mid_0_45_real) + $signed(data_mid_0_45_imag));
  assign _zz_3019 = fixTo_132_dout;
  assign _zz_3020 = ($signed(_zz_113) + $signed(_zz_3021));
  assign _zz_3021 = ($signed(_zz_3022) * $signed(twiddle_factor_table_0_real));
  assign _zz_3022 = ($signed(data_mid_0_45_imag) - $signed(data_mid_0_45_real));
  assign _zz_3023 = fixTo_133_dout;
  assign _zz_3024 = _zz_3025[35 : 0];
  assign _zz_3025 = _zz_3026;
  assign _zz_3026 = ($signed(_zz_3027) >>> _zz_114);
  assign _zz_3027 = _zz_3028;
  assign _zz_3028 = ($signed(_zz_3030) - $signed(_zz_111));
  assign _zz_3029 = ({9'd0,data_mid_0_44_real} <<< 9);
  assign _zz_3030 = {{9{_zz_3029[26]}}, _zz_3029};
  assign _zz_3031 = fixTo_134_dout;
  assign _zz_3032 = _zz_3033[35 : 0];
  assign _zz_3033 = _zz_3034;
  assign _zz_3034 = ($signed(_zz_3035) >>> _zz_114);
  assign _zz_3035 = _zz_3036;
  assign _zz_3036 = ($signed(_zz_3038) - $signed(_zz_112));
  assign _zz_3037 = ({9'd0,data_mid_0_44_imag} <<< 9);
  assign _zz_3038 = {{9{_zz_3037[26]}}, _zz_3037};
  assign _zz_3039 = fixTo_135_dout;
  assign _zz_3040 = _zz_3041[35 : 0];
  assign _zz_3041 = _zz_3042;
  assign _zz_3042 = ($signed(_zz_3043) >>> _zz_115);
  assign _zz_3043 = _zz_3044;
  assign _zz_3044 = ($signed(_zz_3046) + $signed(_zz_111));
  assign _zz_3045 = ({9'd0,data_mid_0_44_real} <<< 9);
  assign _zz_3046 = {{9{_zz_3045[26]}}, _zz_3045};
  assign _zz_3047 = fixTo_136_dout;
  assign _zz_3048 = _zz_3049[35 : 0];
  assign _zz_3049 = _zz_3050;
  assign _zz_3050 = ($signed(_zz_3051) >>> _zz_115);
  assign _zz_3051 = _zz_3052;
  assign _zz_3052 = ($signed(_zz_3054) + $signed(_zz_112));
  assign _zz_3053 = ({9'd0,data_mid_0_44_imag} <<< 9);
  assign _zz_3054 = {{9{_zz_3053[26]}}, _zz_3053};
  assign _zz_3055 = fixTo_137_dout;
  assign _zz_3056 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_3057 = ($signed(_zz_118) - $signed(_zz_3058));
  assign _zz_3058 = ($signed(_zz_3059) * $signed(twiddle_factor_table_0_imag));
  assign _zz_3059 = ($signed(data_mid_0_47_real) + $signed(data_mid_0_47_imag));
  assign _zz_3060 = fixTo_138_dout;
  assign _zz_3061 = ($signed(_zz_118) + $signed(_zz_3062));
  assign _zz_3062 = ($signed(_zz_3063) * $signed(twiddle_factor_table_0_real));
  assign _zz_3063 = ($signed(data_mid_0_47_imag) - $signed(data_mid_0_47_real));
  assign _zz_3064 = fixTo_139_dout;
  assign _zz_3065 = _zz_3066[35 : 0];
  assign _zz_3066 = _zz_3067;
  assign _zz_3067 = ($signed(_zz_3068) >>> _zz_119);
  assign _zz_3068 = _zz_3069;
  assign _zz_3069 = ($signed(_zz_3071) - $signed(_zz_116));
  assign _zz_3070 = ({9'd0,data_mid_0_46_real} <<< 9);
  assign _zz_3071 = {{9{_zz_3070[26]}}, _zz_3070};
  assign _zz_3072 = fixTo_140_dout;
  assign _zz_3073 = _zz_3074[35 : 0];
  assign _zz_3074 = _zz_3075;
  assign _zz_3075 = ($signed(_zz_3076) >>> _zz_119);
  assign _zz_3076 = _zz_3077;
  assign _zz_3077 = ($signed(_zz_3079) - $signed(_zz_117));
  assign _zz_3078 = ({9'd0,data_mid_0_46_imag} <<< 9);
  assign _zz_3079 = {{9{_zz_3078[26]}}, _zz_3078};
  assign _zz_3080 = fixTo_141_dout;
  assign _zz_3081 = _zz_3082[35 : 0];
  assign _zz_3082 = _zz_3083;
  assign _zz_3083 = ($signed(_zz_3084) >>> _zz_120);
  assign _zz_3084 = _zz_3085;
  assign _zz_3085 = ($signed(_zz_3087) + $signed(_zz_116));
  assign _zz_3086 = ({9'd0,data_mid_0_46_real} <<< 9);
  assign _zz_3087 = {{9{_zz_3086[26]}}, _zz_3086};
  assign _zz_3088 = fixTo_142_dout;
  assign _zz_3089 = _zz_3090[35 : 0];
  assign _zz_3090 = _zz_3091;
  assign _zz_3091 = ($signed(_zz_3092) >>> _zz_120);
  assign _zz_3092 = _zz_3093;
  assign _zz_3093 = ($signed(_zz_3095) + $signed(_zz_117));
  assign _zz_3094 = ({9'd0,data_mid_0_46_imag} <<< 9);
  assign _zz_3095 = {{9{_zz_3094[26]}}, _zz_3094};
  assign _zz_3096 = fixTo_143_dout;
  assign _zz_3097 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_3098 = ($signed(_zz_123) - $signed(_zz_3099));
  assign _zz_3099 = ($signed(_zz_3100) * $signed(twiddle_factor_table_0_imag));
  assign _zz_3100 = ($signed(data_mid_0_49_real) + $signed(data_mid_0_49_imag));
  assign _zz_3101 = fixTo_144_dout;
  assign _zz_3102 = ($signed(_zz_123) + $signed(_zz_3103));
  assign _zz_3103 = ($signed(_zz_3104) * $signed(twiddle_factor_table_0_real));
  assign _zz_3104 = ($signed(data_mid_0_49_imag) - $signed(data_mid_0_49_real));
  assign _zz_3105 = fixTo_145_dout;
  assign _zz_3106 = _zz_3107[35 : 0];
  assign _zz_3107 = _zz_3108;
  assign _zz_3108 = ($signed(_zz_3109) >>> _zz_124);
  assign _zz_3109 = _zz_3110;
  assign _zz_3110 = ($signed(_zz_3112) - $signed(_zz_121));
  assign _zz_3111 = ({9'd0,data_mid_0_48_real} <<< 9);
  assign _zz_3112 = {{9{_zz_3111[26]}}, _zz_3111};
  assign _zz_3113 = fixTo_146_dout;
  assign _zz_3114 = _zz_3115[35 : 0];
  assign _zz_3115 = _zz_3116;
  assign _zz_3116 = ($signed(_zz_3117) >>> _zz_124);
  assign _zz_3117 = _zz_3118;
  assign _zz_3118 = ($signed(_zz_3120) - $signed(_zz_122));
  assign _zz_3119 = ({9'd0,data_mid_0_48_imag} <<< 9);
  assign _zz_3120 = {{9{_zz_3119[26]}}, _zz_3119};
  assign _zz_3121 = fixTo_147_dout;
  assign _zz_3122 = _zz_3123[35 : 0];
  assign _zz_3123 = _zz_3124;
  assign _zz_3124 = ($signed(_zz_3125) >>> _zz_125);
  assign _zz_3125 = _zz_3126;
  assign _zz_3126 = ($signed(_zz_3128) + $signed(_zz_121));
  assign _zz_3127 = ({9'd0,data_mid_0_48_real} <<< 9);
  assign _zz_3128 = {{9{_zz_3127[26]}}, _zz_3127};
  assign _zz_3129 = fixTo_148_dout;
  assign _zz_3130 = _zz_3131[35 : 0];
  assign _zz_3131 = _zz_3132;
  assign _zz_3132 = ($signed(_zz_3133) >>> _zz_125);
  assign _zz_3133 = _zz_3134;
  assign _zz_3134 = ($signed(_zz_3136) + $signed(_zz_122));
  assign _zz_3135 = ({9'd0,data_mid_0_48_imag} <<< 9);
  assign _zz_3136 = {{9{_zz_3135[26]}}, _zz_3135};
  assign _zz_3137 = fixTo_149_dout;
  assign _zz_3138 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_3139 = ($signed(_zz_128) - $signed(_zz_3140));
  assign _zz_3140 = ($signed(_zz_3141) * $signed(twiddle_factor_table_0_imag));
  assign _zz_3141 = ($signed(data_mid_0_51_real) + $signed(data_mid_0_51_imag));
  assign _zz_3142 = fixTo_150_dout;
  assign _zz_3143 = ($signed(_zz_128) + $signed(_zz_3144));
  assign _zz_3144 = ($signed(_zz_3145) * $signed(twiddle_factor_table_0_real));
  assign _zz_3145 = ($signed(data_mid_0_51_imag) - $signed(data_mid_0_51_real));
  assign _zz_3146 = fixTo_151_dout;
  assign _zz_3147 = _zz_3148[35 : 0];
  assign _zz_3148 = _zz_3149;
  assign _zz_3149 = ($signed(_zz_3150) >>> _zz_129);
  assign _zz_3150 = _zz_3151;
  assign _zz_3151 = ($signed(_zz_3153) - $signed(_zz_126));
  assign _zz_3152 = ({9'd0,data_mid_0_50_real} <<< 9);
  assign _zz_3153 = {{9{_zz_3152[26]}}, _zz_3152};
  assign _zz_3154 = fixTo_152_dout;
  assign _zz_3155 = _zz_3156[35 : 0];
  assign _zz_3156 = _zz_3157;
  assign _zz_3157 = ($signed(_zz_3158) >>> _zz_129);
  assign _zz_3158 = _zz_3159;
  assign _zz_3159 = ($signed(_zz_3161) - $signed(_zz_127));
  assign _zz_3160 = ({9'd0,data_mid_0_50_imag} <<< 9);
  assign _zz_3161 = {{9{_zz_3160[26]}}, _zz_3160};
  assign _zz_3162 = fixTo_153_dout;
  assign _zz_3163 = _zz_3164[35 : 0];
  assign _zz_3164 = _zz_3165;
  assign _zz_3165 = ($signed(_zz_3166) >>> _zz_130);
  assign _zz_3166 = _zz_3167;
  assign _zz_3167 = ($signed(_zz_3169) + $signed(_zz_126));
  assign _zz_3168 = ({9'd0,data_mid_0_50_real} <<< 9);
  assign _zz_3169 = {{9{_zz_3168[26]}}, _zz_3168};
  assign _zz_3170 = fixTo_154_dout;
  assign _zz_3171 = _zz_3172[35 : 0];
  assign _zz_3172 = _zz_3173;
  assign _zz_3173 = ($signed(_zz_3174) >>> _zz_130);
  assign _zz_3174 = _zz_3175;
  assign _zz_3175 = ($signed(_zz_3177) + $signed(_zz_127));
  assign _zz_3176 = ({9'd0,data_mid_0_50_imag} <<< 9);
  assign _zz_3177 = {{9{_zz_3176[26]}}, _zz_3176};
  assign _zz_3178 = fixTo_155_dout;
  assign _zz_3179 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_3180 = ($signed(_zz_133) - $signed(_zz_3181));
  assign _zz_3181 = ($signed(_zz_3182) * $signed(twiddle_factor_table_0_imag));
  assign _zz_3182 = ($signed(data_mid_0_53_real) + $signed(data_mid_0_53_imag));
  assign _zz_3183 = fixTo_156_dout;
  assign _zz_3184 = ($signed(_zz_133) + $signed(_zz_3185));
  assign _zz_3185 = ($signed(_zz_3186) * $signed(twiddle_factor_table_0_real));
  assign _zz_3186 = ($signed(data_mid_0_53_imag) - $signed(data_mid_0_53_real));
  assign _zz_3187 = fixTo_157_dout;
  assign _zz_3188 = _zz_3189[35 : 0];
  assign _zz_3189 = _zz_3190;
  assign _zz_3190 = ($signed(_zz_3191) >>> _zz_134);
  assign _zz_3191 = _zz_3192;
  assign _zz_3192 = ($signed(_zz_3194) - $signed(_zz_131));
  assign _zz_3193 = ({9'd0,data_mid_0_52_real} <<< 9);
  assign _zz_3194 = {{9{_zz_3193[26]}}, _zz_3193};
  assign _zz_3195 = fixTo_158_dout;
  assign _zz_3196 = _zz_3197[35 : 0];
  assign _zz_3197 = _zz_3198;
  assign _zz_3198 = ($signed(_zz_3199) >>> _zz_134);
  assign _zz_3199 = _zz_3200;
  assign _zz_3200 = ($signed(_zz_3202) - $signed(_zz_132));
  assign _zz_3201 = ({9'd0,data_mid_0_52_imag} <<< 9);
  assign _zz_3202 = {{9{_zz_3201[26]}}, _zz_3201};
  assign _zz_3203 = fixTo_159_dout;
  assign _zz_3204 = _zz_3205[35 : 0];
  assign _zz_3205 = _zz_3206;
  assign _zz_3206 = ($signed(_zz_3207) >>> _zz_135);
  assign _zz_3207 = _zz_3208;
  assign _zz_3208 = ($signed(_zz_3210) + $signed(_zz_131));
  assign _zz_3209 = ({9'd0,data_mid_0_52_real} <<< 9);
  assign _zz_3210 = {{9{_zz_3209[26]}}, _zz_3209};
  assign _zz_3211 = fixTo_160_dout;
  assign _zz_3212 = _zz_3213[35 : 0];
  assign _zz_3213 = _zz_3214;
  assign _zz_3214 = ($signed(_zz_3215) >>> _zz_135);
  assign _zz_3215 = _zz_3216;
  assign _zz_3216 = ($signed(_zz_3218) + $signed(_zz_132));
  assign _zz_3217 = ({9'd0,data_mid_0_52_imag} <<< 9);
  assign _zz_3218 = {{9{_zz_3217[26]}}, _zz_3217};
  assign _zz_3219 = fixTo_161_dout;
  assign _zz_3220 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_3221 = ($signed(_zz_138) - $signed(_zz_3222));
  assign _zz_3222 = ($signed(_zz_3223) * $signed(twiddle_factor_table_0_imag));
  assign _zz_3223 = ($signed(data_mid_0_55_real) + $signed(data_mid_0_55_imag));
  assign _zz_3224 = fixTo_162_dout;
  assign _zz_3225 = ($signed(_zz_138) + $signed(_zz_3226));
  assign _zz_3226 = ($signed(_zz_3227) * $signed(twiddle_factor_table_0_real));
  assign _zz_3227 = ($signed(data_mid_0_55_imag) - $signed(data_mid_0_55_real));
  assign _zz_3228 = fixTo_163_dout;
  assign _zz_3229 = _zz_3230[35 : 0];
  assign _zz_3230 = _zz_3231;
  assign _zz_3231 = ($signed(_zz_3232) >>> _zz_139);
  assign _zz_3232 = _zz_3233;
  assign _zz_3233 = ($signed(_zz_3235) - $signed(_zz_136));
  assign _zz_3234 = ({9'd0,data_mid_0_54_real} <<< 9);
  assign _zz_3235 = {{9{_zz_3234[26]}}, _zz_3234};
  assign _zz_3236 = fixTo_164_dout;
  assign _zz_3237 = _zz_3238[35 : 0];
  assign _zz_3238 = _zz_3239;
  assign _zz_3239 = ($signed(_zz_3240) >>> _zz_139);
  assign _zz_3240 = _zz_3241;
  assign _zz_3241 = ($signed(_zz_3243) - $signed(_zz_137));
  assign _zz_3242 = ({9'd0,data_mid_0_54_imag} <<< 9);
  assign _zz_3243 = {{9{_zz_3242[26]}}, _zz_3242};
  assign _zz_3244 = fixTo_165_dout;
  assign _zz_3245 = _zz_3246[35 : 0];
  assign _zz_3246 = _zz_3247;
  assign _zz_3247 = ($signed(_zz_3248) >>> _zz_140);
  assign _zz_3248 = _zz_3249;
  assign _zz_3249 = ($signed(_zz_3251) + $signed(_zz_136));
  assign _zz_3250 = ({9'd0,data_mid_0_54_real} <<< 9);
  assign _zz_3251 = {{9{_zz_3250[26]}}, _zz_3250};
  assign _zz_3252 = fixTo_166_dout;
  assign _zz_3253 = _zz_3254[35 : 0];
  assign _zz_3254 = _zz_3255;
  assign _zz_3255 = ($signed(_zz_3256) >>> _zz_140);
  assign _zz_3256 = _zz_3257;
  assign _zz_3257 = ($signed(_zz_3259) + $signed(_zz_137));
  assign _zz_3258 = ({9'd0,data_mid_0_54_imag} <<< 9);
  assign _zz_3259 = {{9{_zz_3258[26]}}, _zz_3258};
  assign _zz_3260 = fixTo_167_dout;
  assign _zz_3261 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_3262 = ($signed(_zz_143) - $signed(_zz_3263));
  assign _zz_3263 = ($signed(_zz_3264) * $signed(twiddle_factor_table_0_imag));
  assign _zz_3264 = ($signed(data_mid_0_57_real) + $signed(data_mid_0_57_imag));
  assign _zz_3265 = fixTo_168_dout;
  assign _zz_3266 = ($signed(_zz_143) + $signed(_zz_3267));
  assign _zz_3267 = ($signed(_zz_3268) * $signed(twiddle_factor_table_0_real));
  assign _zz_3268 = ($signed(data_mid_0_57_imag) - $signed(data_mid_0_57_real));
  assign _zz_3269 = fixTo_169_dout;
  assign _zz_3270 = _zz_3271[35 : 0];
  assign _zz_3271 = _zz_3272;
  assign _zz_3272 = ($signed(_zz_3273) >>> _zz_144);
  assign _zz_3273 = _zz_3274;
  assign _zz_3274 = ($signed(_zz_3276) - $signed(_zz_141));
  assign _zz_3275 = ({9'd0,data_mid_0_56_real} <<< 9);
  assign _zz_3276 = {{9{_zz_3275[26]}}, _zz_3275};
  assign _zz_3277 = fixTo_170_dout;
  assign _zz_3278 = _zz_3279[35 : 0];
  assign _zz_3279 = _zz_3280;
  assign _zz_3280 = ($signed(_zz_3281) >>> _zz_144);
  assign _zz_3281 = _zz_3282;
  assign _zz_3282 = ($signed(_zz_3284) - $signed(_zz_142));
  assign _zz_3283 = ({9'd0,data_mid_0_56_imag} <<< 9);
  assign _zz_3284 = {{9{_zz_3283[26]}}, _zz_3283};
  assign _zz_3285 = fixTo_171_dout;
  assign _zz_3286 = _zz_3287[35 : 0];
  assign _zz_3287 = _zz_3288;
  assign _zz_3288 = ($signed(_zz_3289) >>> _zz_145);
  assign _zz_3289 = _zz_3290;
  assign _zz_3290 = ($signed(_zz_3292) + $signed(_zz_141));
  assign _zz_3291 = ({9'd0,data_mid_0_56_real} <<< 9);
  assign _zz_3292 = {{9{_zz_3291[26]}}, _zz_3291};
  assign _zz_3293 = fixTo_172_dout;
  assign _zz_3294 = _zz_3295[35 : 0];
  assign _zz_3295 = _zz_3296;
  assign _zz_3296 = ($signed(_zz_3297) >>> _zz_145);
  assign _zz_3297 = _zz_3298;
  assign _zz_3298 = ($signed(_zz_3300) + $signed(_zz_142));
  assign _zz_3299 = ({9'd0,data_mid_0_56_imag} <<< 9);
  assign _zz_3300 = {{9{_zz_3299[26]}}, _zz_3299};
  assign _zz_3301 = fixTo_173_dout;
  assign _zz_3302 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_3303 = ($signed(_zz_148) - $signed(_zz_3304));
  assign _zz_3304 = ($signed(_zz_3305) * $signed(twiddle_factor_table_0_imag));
  assign _zz_3305 = ($signed(data_mid_0_59_real) + $signed(data_mid_0_59_imag));
  assign _zz_3306 = fixTo_174_dout;
  assign _zz_3307 = ($signed(_zz_148) + $signed(_zz_3308));
  assign _zz_3308 = ($signed(_zz_3309) * $signed(twiddle_factor_table_0_real));
  assign _zz_3309 = ($signed(data_mid_0_59_imag) - $signed(data_mid_0_59_real));
  assign _zz_3310 = fixTo_175_dout;
  assign _zz_3311 = _zz_3312[35 : 0];
  assign _zz_3312 = _zz_3313;
  assign _zz_3313 = ($signed(_zz_3314) >>> _zz_149);
  assign _zz_3314 = _zz_3315;
  assign _zz_3315 = ($signed(_zz_3317) - $signed(_zz_146));
  assign _zz_3316 = ({9'd0,data_mid_0_58_real} <<< 9);
  assign _zz_3317 = {{9{_zz_3316[26]}}, _zz_3316};
  assign _zz_3318 = fixTo_176_dout;
  assign _zz_3319 = _zz_3320[35 : 0];
  assign _zz_3320 = _zz_3321;
  assign _zz_3321 = ($signed(_zz_3322) >>> _zz_149);
  assign _zz_3322 = _zz_3323;
  assign _zz_3323 = ($signed(_zz_3325) - $signed(_zz_147));
  assign _zz_3324 = ({9'd0,data_mid_0_58_imag} <<< 9);
  assign _zz_3325 = {{9{_zz_3324[26]}}, _zz_3324};
  assign _zz_3326 = fixTo_177_dout;
  assign _zz_3327 = _zz_3328[35 : 0];
  assign _zz_3328 = _zz_3329;
  assign _zz_3329 = ($signed(_zz_3330) >>> _zz_150);
  assign _zz_3330 = _zz_3331;
  assign _zz_3331 = ($signed(_zz_3333) + $signed(_zz_146));
  assign _zz_3332 = ({9'd0,data_mid_0_58_real} <<< 9);
  assign _zz_3333 = {{9{_zz_3332[26]}}, _zz_3332};
  assign _zz_3334 = fixTo_178_dout;
  assign _zz_3335 = _zz_3336[35 : 0];
  assign _zz_3336 = _zz_3337;
  assign _zz_3337 = ($signed(_zz_3338) >>> _zz_150);
  assign _zz_3338 = _zz_3339;
  assign _zz_3339 = ($signed(_zz_3341) + $signed(_zz_147));
  assign _zz_3340 = ({9'd0,data_mid_0_58_imag} <<< 9);
  assign _zz_3341 = {{9{_zz_3340[26]}}, _zz_3340};
  assign _zz_3342 = fixTo_179_dout;
  assign _zz_3343 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_3344 = ($signed(_zz_153) - $signed(_zz_3345));
  assign _zz_3345 = ($signed(_zz_3346) * $signed(twiddle_factor_table_0_imag));
  assign _zz_3346 = ($signed(data_mid_0_61_real) + $signed(data_mid_0_61_imag));
  assign _zz_3347 = fixTo_180_dout;
  assign _zz_3348 = ($signed(_zz_153) + $signed(_zz_3349));
  assign _zz_3349 = ($signed(_zz_3350) * $signed(twiddle_factor_table_0_real));
  assign _zz_3350 = ($signed(data_mid_0_61_imag) - $signed(data_mid_0_61_real));
  assign _zz_3351 = fixTo_181_dout;
  assign _zz_3352 = _zz_3353[35 : 0];
  assign _zz_3353 = _zz_3354;
  assign _zz_3354 = ($signed(_zz_3355) >>> _zz_154);
  assign _zz_3355 = _zz_3356;
  assign _zz_3356 = ($signed(_zz_3358) - $signed(_zz_151));
  assign _zz_3357 = ({9'd0,data_mid_0_60_real} <<< 9);
  assign _zz_3358 = {{9{_zz_3357[26]}}, _zz_3357};
  assign _zz_3359 = fixTo_182_dout;
  assign _zz_3360 = _zz_3361[35 : 0];
  assign _zz_3361 = _zz_3362;
  assign _zz_3362 = ($signed(_zz_3363) >>> _zz_154);
  assign _zz_3363 = _zz_3364;
  assign _zz_3364 = ($signed(_zz_3366) - $signed(_zz_152));
  assign _zz_3365 = ({9'd0,data_mid_0_60_imag} <<< 9);
  assign _zz_3366 = {{9{_zz_3365[26]}}, _zz_3365};
  assign _zz_3367 = fixTo_183_dout;
  assign _zz_3368 = _zz_3369[35 : 0];
  assign _zz_3369 = _zz_3370;
  assign _zz_3370 = ($signed(_zz_3371) >>> _zz_155);
  assign _zz_3371 = _zz_3372;
  assign _zz_3372 = ($signed(_zz_3374) + $signed(_zz_151));
  assign _zz_3373 = ({9'd0,data_mid_0_60_real} <<< 9);
  assign _zz_3374 = {{9{_zz_3373[26]}}, _zz_3373};
  assign _zz_3375 = fixTo_184_dout;
  assign _zz_3376 = _zz_3377[35 : 0];
  assign _zz_3377 = _zz_3378;
  assign _zz_3378 = ($signed(_zz_3379) >>> _zz_155);
  assign _zz_3379 = _zz_3380;
  assign _zz_3380 = ($signed(_zz_3382) + $signed(_zz_152));
  assign _zz_3381 = ({9'd0,data_mid_0_60_imag} <<< 9);
  assign _zz_3382 = {{9{_zz_3381[26]}}, _zz_3381};
  assign _zz_3383 = fixTo_185_dout;
  assign _zz_3384 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_3385 = ($signed(_zz_158) - $signed(_zz_3386));
  assign _zz_3386 = ($signed(_zz_3387) * $signed(twiddle_factor_table_0_imag));
  assign _zz_3387 = ($signed(data_mid_0_63_real) + $signed(data_mid_0_63_imag));
  assign _zz_3388 = fixTo_186_dout;
  assign _zz_3389 = ($signed(_zz_158) + $signed(_zz_3390));
  assign _zz_3390 = ($signed(_zz_3391) * $signed(twiddle_factor_table_0_real));
  assign _zz_3391 = ($signed(data_mid_0_63_imag) - $signed(data_mid_0_63_real));
  assign _zz_3392 = fixTo_187_dout;
  assign _zz_3393 = _zz_3394[35 : 0];
  assign _zz_3394 = _zz_3395;
  assign _zz_3395 = ($signed(_zz_3396) >>> _zz_159);
  assign _zz_3396 = _zz_3397;
  assign _zz_3397 = ($signed(_zz_3399) - $signed(_zz_156));
  assign _zz_3398 = ({9'd0,data_mid_0_62_real} <<< 9);
  assign _zz_3399 = {{9{_zz_3398[26]}}, _zz_3398};
  assign _zz_3400 = fixTo_188_dout;
  assign _zz_3401 = _zz_3402[35 : 0];
  assign _zz_3402 = _zz_3403;
  assign _zz_3403 = ($signed(_zz_3404) >>> _zz_159);
  assign _zz_3404 = _zz_3405;
  assign _zz_3405 = ($signed(_zz_3407) - $signed(_zz_157));
  assign _zz_3406 = ({9'd0,data_mid_0_62_imag} <<< 9);
  assign _zz_3407 = {{9{_zz_3406[26]}}, _zz_3406};
  assign _zz_3408 = fixTo_189_dout;
  assign _zz_3409 = _zz_3410[35 : 0];
  assign _zz_3410 = _zz_3411;
  assign _zz_3411 = ($signed(_zz_3412) >>> _zz_160);
  assign _zz_3412 = _zz_3413;
  assign _zz_3413 = ($signed(_zz_3415) + $signed(_zz_156));
  assign _zz_3414 = ({9'd0,data_mid_0_62_real} <<< 9);
  assign _zz_3415 = {{9{_zz_3414[26]}}, _zz_3414};
  assign _zz_3416 = fixTo_190_dout;
  assign _zz_3417 = _zz_3418[35 : 0];
  assign _zz_3418 = _zz_3419;
  assign _zz_3419 = ($signed(_zz_3420) >>> _zz_160);
  assign _zz_3420 = _zz_3421;
  assign _zz_3421 = ($signed(_zz_3423) + $signed(_zz_157));
  assign _zz_3422 = ({9'd0,data_mid_0_62_imag} <<< 9);
  assign _zz_3423 = {{9{_zz_3422[26]}}, _zz_3422};
  assign _zz_3424 = fixTo_191_dout;
  assign _zz_3425 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_3426 = ($signed(_zz_163) - $signed(_zz_3427));
  assign _zz_3427 = ($signed(_zz_3428) * $signed(twiddle_factor_table_1_imag));
  assign _zz_3428 = ($signed(data_mid_1_2_real) + $signed(data_mid_1_2_imag));
  assign _zz_3429 = fixTo_192_dout;
  assign _zz_3430 = ($signed(_zz_163) + $signed(_zz_3431));
  assign _zz_3431 = ($signed(_zz_3432) * $signed(twiddle_factor_table_1_real));
  assign _zz_3432 = ($signed(data_mid_1_2_imag) - $signed(data_mid_1_2_real));
  assign _zz_3433 = fixTo_193_dout;
  assign _zz_3434 = _zz_3435[35 : 0];
  assign _zz_3435 = _zz_3436;
  assign _zz_3436 = ($signed(_zz_3437) >>> _zz_164);
  assign _zz_3437 = _zz_3438;
  assign _zz_3438 = ($signed(_zz_3440) - $signed(_zz_161));
  assign _zz_3439 = ({9'd0,data_mid_1_0_real} <<< 9);
  assign _zz_3440 = {{9{_zz_3439[26]}}, _zz_3439};
  assign _zz_3441 = fixTo_194_dout;
  assign _zz_3442 = _zz_3443[35 : 0];
  assign _zz_3443 = _zz_3444;
  assign _zz_3444 = ($signed(_zz_3445) >>> _zz_164);
  assign _zz_3445 = _zz_3446;
  assign _zz_3446 = ($signed(_zz_3448) - $signed(_zz_162));
  assign _zz_3447 = ({9'd0,data_mid_1_0_imag} <<< 9);
  assign _zz_3448 = {{9{_zz_3447[26]}}, _zz_3447};
  assign _zz_3449 = fixTo_195_dout;
  assign _zz_3450 = _zz_3451[35 : 0];
  assign _zz_3451 = _zz_3452;
  assign _zz_3452 = ($signed(_zz_3453) >>> _zz_165);
  assign _zz_3453 = _zz_3454;
  assign _zz_3454 = ($signed(_zz_3456) + $signed(_zz_161));
  assign _zz_3455 = ({9'd0,data_mid_1_0_real} <<< 9);
  assign _zz_3456 = {{9{_zz_3455[26]}}, _zz_3455};
  assign _zz_3457 = fixTo_196_dout;
  assign _zz_3458 = _zz_3459[35 : 0];
  assign _zz_3459 = _zz_3460;
  assign _zz_3460 = ($signed(_zz_3461) >>> _zz_165);
  assign _zz_3461 = _zz_3462;
  assign _zz_3462 = ($signed(_zz_3464) + $signed(_zz_162));
  assign _zz_3463 = ({9'd0,data_mid_1_0_imag} <<< 9);
  assign _zz_3464 = {{9{_zz_3463[26]}}, _zz_3463};
  assign _zz_3465 = fixTo_197_dout;
  assign _zz_3466 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_3467 = ($signed(_zz_168) - $signed(_zz_3468));
  assign _zz_3468 = ($signed(_zz_3469) * $signed(twiddle_factor_table_2_imag));
  assign _zz_3469 = ($signed(data_mid_1_3_real) + $signed(data_mid_1_3_imag));
  assign _zz_3470 = fixTo_198_dout;
  assign _zz_3471 = ($signed(_zz_168) + $signed(_zz_3472));
  assign _zz_3472 = ($signed(_zz_3473) * $signed(twiddle_factor_table_2_real));
  assign _zz_3473 = ($signed(data_mid_1_3_imag) - $signed(data_mid_1_3_real));
  assign _zz_3474 = fixTo_199_dout;
  assign _zz_3475 = _zz_3476[35 : 0];
  assign _zz_3476 = _zz_3477;
  assign _zz_3477 = ($signed(_zz_3478) >>> _zz_169);
  assign _zz_3478 = _zz_3479;
  assign _zz_3479 = ($signed(_zz_3481) - $signed(_zz_166));
  assign _zz_3480 = ({9'd0,data_mid_1_1_real} <<< 9);
  assign _zz_3481 = {{9{_zz_3480[26]}}, _zz_3480};
  assign _zz_3482 = fixTo_200_dout;
  assign _zz_3483 = _zz_3484[35 : 0];
  assign _zz_3484 = _zz_3485;
  assign _zz_3485 = ($signed(_zz_3486) >>> _zz_169);
  assign _zz_3486 = _zz_3487;
  assign _zz_3487 = ($signed(_zz_3489) - $signed(_zz_167));
  assign _zz_3488 = ({9'd0,data_mid_1_1_imag} <<< 9);
  assign _zz_3489 = {{9{_zz_3488[26]}}, _zz_3488};
  assign _zz_3490 = fixTo_201_dout;
  assign _zz_3491 = _zz_3492[35 : 0];
  assign _zz_3492 = _zz_3493;
  assign _zz_3493 = ($signed(_zz_3494) >>> _zz_170);
  assign _zz_3494 = _zz_3495;
  assign _zz_3495 = ($signed(_zz_3497) + $signed(_zz_166));
  assign _zz_3496 = ({9'd0,data_mid_1_1_real} <<< 9);
  assign _zz_3497 = {{9{_zz_3496[26]}}, _zz_3496};
  assign _zz_3498 = fixTo_202_dout;
  assign _zz_3499 = _zz_3500[35 : 0];
  assign _zz_3500 = _zz_3501;
  assign _zz_3501 = ($signed(_zz_3502) >>> _zz_170);
  assign _zz_3502 = _zz_3503;
  assign _zz_3503 = ($signed(_zz_3505) + $signed(_zz_167));
  assign _zz_3504 = ({9'd0,data_mid_1_1_imag} <<< 9);
  assign _zz_3505 = {{9{_zz_3504[26]}}, _zz_3504};
  assign _zz_3506 = fixTo_203_dout;
  assign _zz_3507 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_3508 = ($signed(_zz_173) - $signed(_zz_3509));
  assign _zz_3509 = ($signed(_zz_3510) * $signed(twiddle_factor_table_1_imag));
  assign _zz_3510 = ($signed(data_mid_1_6_real) + $signed(data_mid_1_6_imag));
  assign _zz_3511 = fixTo_204_dout;
  assign _zz_3512 = ($signed(_zz_173) + $signed(_zz_3513));
  assign _zz_3513 = ($signed(_zz_3514) * $signed(twiddle_factor_table_1_real));
  assign _zz_3514 = ($signed(data_mid_1_6_imag) - $signed(data_mid_1_6_real));
  assign _zz_3515 = fixTo_205_dout;
  assign _zz_3516 = _zz_3517[35 : 0];
  assign _zz_3517 = _zz_3518;
  assign _zz_3518 = ($signed(_zz_3519) >>> _zz_174);
  assign _zz_3519 = _zz_3520;
  assign _zz_3520 = ($signed(_zz_3522) - $signed(_zz_171));
  assign _zz_3521 = ({9'd0,data_mid_1_4_real} <<< 9);
  assign _zz_3522 = {{9{_zz_3521[26]}}, _zz_3521};
  assign _zz_3523 = fixTo_206_dout;
  assign _zz_3524 = _zz_3525[35 : 0];
  assign _zz_3525 = _zz_3526;
  assign _zz_3526 = ($signed(_zz_3527) >>> _zz_174);
  assign _zz_3527 = _zz_3528;
  assign _zz_3528 = ($signed(_zz_3530) - $signed(_zz_172));
  assign _zz_3529 = ({9'd0,data_mid_1_4_imag} <<< 9);
  assign _zz_3530 = {{9{_zz_3529[26]}}, _zz_3529};
  assign _zz_3531 = fixTo_207_dout;
  assign _zz_3532 = _zz_3533[35 : 0];
  assign _zz_3533 = _zz_3534;
  assign _zz_3534 = ($signed(_zz_3535) >>> _zz_175);
  assign _zz_3535 = _zz_3536;
  assign _zz_3536 = ($signed(_zz_3538) + $signed(_zz_171));
  assign _zz_3537 = ({9'd0,data_mid_1_4_real} <<< 9);
  assign _zz_3538 = {{9{_zz_3537[26]}}, _zz_3537};
  assign _zz_3539 = fixTo_208_dout;
  assign _zz_3540 = _zz_3541[35 : 0];
  assign _zz_3541 = _zz_3542;
  assign _zz_3542 = ($signed(_zz_3543) >>> _zz_175);
  assign _zz_3543 = _zz_3544;
  assign _zz_3544 = ($signed(_zz_3546) + $signed(_zz_172));
  assign _zz_3545 = ({9'd0,data_mid_1_4_imag} <<< 9);
  assign _zz_3546 = {{9{_zz_3545[26]}}, _zz_3545};
  assign _zz_3547 = fixTo_209_dout;
  assign _zz_3548 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_3549 = ($signed(_zz_178) - $signed(_zz_3550));
  assign _zz_3550 = ($signed(_zz_3551) * $signed(twiddle_factor_table_2_imag));
  assign _zz_3551 = ($signed(data_mid_1_7_real) + $signed(data_mid_1_7_imag));
  assign _zz_3552 = fixTo_210_dout;
  assign _zz_3553 = ($signed(_zz_178) + $signed(_zz_3554));
  assign _zz_3554 = ($signed(_zz_3555) * $signed(twiddle_factor_table_2_real));
  assign _zz_3555 = ($signed(data_mid_1_7_imag) - $signed(data_mid_1_7_real));
  assign _zz_3556 = fixTo_211_dout;
  assign _zz_3557 = _zz_3558[35 : 0];
  assign _zz_3558 = _zz_3559;
  assign _zz_3559 = ($signed(_zz_3560) >>> _zz_179);
  assign _zz_3560 = _zz_3561;
  assign _zz_3561 = ($signed(_zz_3563) - $signed(_zz_176));
  assign _zz_3562 = ({9'd0,data_mid_1_5_real} <<< 9);
  assign _zz_3563 = {{9{_zz_3562[26]}}, _zz_3562};
  assign _zz_3564 = fixTo_212_dout;
  assign _zz_3565 = _zz_3566[35 : 0];
  assign _zz_3566 = _zz_3567;
  assign _zz_3567 = ($signed(_zz_3568) >>> _zz_179);
  assign _zz_3568 = _zz_3569;
  assign _zz_3569 = ($signed(_zz_3571) - $signed(_zz_177));
  assign _zz_3570 = ({9'd0,data_mid_1_5_imag} <<< 9);
  assign _zz_3571 = {{9{_zz_3570[26]}}, _zz_3570};
  assign _zz_3572 = fixTo_213_dout;
  assign _zz_3573 = _zz_3574[35 : 0];
  assign _zz_3574 = _zz_3575;
  assign _zz_3575 = ($signed(_zz_3576) >>> _zz_180);
  assign _zz_3576 = _zz_3577;
  assign _zz_3577 = ($signed(_zz_3579) + $signed(_zz_176));
  assign _zz_3578 = ({9'd0,data_mid_1_5_real} <<< 9);
  assign _zz_3579 = {{9{_zz_3578[26]}}, _zz_3578};
  assign _zz_3580 = fixTo_214_dout;
  assign _zz_3581 = _zz_3582[35 : 0];
  assign _zz_3582 = _zz_3583;
  assign _zz_3583 = ($signed(_zz_3584) >>> _zz_180);
  assign _zz_3584 = _zz_3585;
  assign _zz_3585 = ($signed(_zz_3587) + $signed(_zz_177));
  assign _zz_3586 = ({9'd0,data_mid_1_5_imag} <<< 9);
  assign _zz_3587 = {{9{_zz_3586[26]}}, _zz_3586};
  assign _zz_3588 = fixTo_215_dout;
  assign _zz_3589 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_3590 = ($signed(_zz_183) - $signed(_zz_3591));
  assign _zz_3591 = ($signed(_zz_3592) * $signed(twiddle_factor_table_1_imag));
  assign _zz_3592 = ($signed(data_mid_1_10_real) + $signed(data_mid_1_10_imag));
  assign _zz_3593 = fixTo_216_dout;
  assign _zz_3594 = ($signed(_zz_183) + $signed(_zz_3595));
  assign _zz_3595 = ($signed(_zz_3596) * $signed(twiddle_factor_table_1_real));
  assign _zz_3596 = ($signed(data_mid_1_10_imag) - $signed(data_mid_1_10_real));
  assign _zz_3597 = fixTo_217_dout;
  assign _zz_3598 = _zz_3599[35 : 0];
  assign _zz_3599 = _zz_3600;
  assign _zz_3600 = ($signed(_zz_3601) >>> _zz_184);
  assign _zz_3601 = _zz_3602;
  assign _zz_3602 = ($signed(_zz_3604) - $signed(_zz_181));
  assign _zz_3603 = ({9'd0,data_mid_1_8_real} <<< 9);
  assign _zz_3604 = {{9{_zz_3603[26]}}, _zz_3603};
  assign _zz_3605 = fixTo_218_dout;
  assign _zz_3606 = _zz_3607[35 : 0];
  assign _zz_3607 = _zz_3608;
  assign _zz_3608 = ($signed(_zz_3609) >>> _zz_184);
  assign _zz_3609 = _zz_3610;
  assign _zz_3610 = ($signed(_zz_3612) - $signed(_zz_182));
  assign _zz_3611 = ({9'd0,data_mid_1_8_imag} <<< 9);
  assign _zz_3612 = {{9{_zz_3611[26]}}, _zz_3611};
  assign _zz_3613 = fixTo_219_dout;
  assign _zz_3614 = _zz_3615[35 : 0];
  assign _zz_3615 = _zz_3616;
  assign _zz_3616 = ($signed(_zz_3617) >>> _zz_185);
  assign _zz_3617 = _zz_3618;
  assign _zz_3618 = ($signed(_zz_3620) + $signed(_zz_181));
  assign _zz_3619 = ({9'd0,data_mid_1_8_real} <<< 9);
  assign _zz_3620 = {{9{_zz_3619[26]}}, _zz_3619};
  assign _zz_3621 = fixTo_220_dout;
  assign _zz_3622 = _zz_3623[35 : 0];
  assign _zz_3623 = _zz_3624;
  assign _zz_3624 = ($signed(_zz_3625) >>> _zz_185);
  assign _zz_3625 = _zz_3626;
  assign _zz_3626 = ($signed(_zz_3628) + $signed(_zz_182));
  assign _zz_3627 = ({9'd0,data_mid_1_8_imag} <<< 9);
  assign _zz_3628 = {{9{_zz_3627[26]}}, _zz_3627};
  assign _zz_3629 = fixTo_221_dout;
  assign _zz_3630 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_3631 = ($signed(_zz_188) - $signed(_zz_3632));
  assign _zz_3632 = ($signed(_zz_3633) * $signed(twiddle_factor_table_2_imag));
  assign _zz_3633 = ($signed(data_mid_1_11_real) + $signed(data_mid_1_11_imag));
  assign _zz_3634 = fixTo_222_dout;
  assign _zz_3635 = ($signed(_zz_188) + $signed(_zz_3636));
  assign _zz_3636 = ($signed(_zz_3637) * $signed(twiddle_factor_table_2_real));
  assign _zz_3637 = ($signed(data_mid_1_11_imag) - $signed(data_mid_1_11_real));
  assign _zz_3638 = fixTo_223_dout;
  assign _zz_3639 = _zz_3640[35 : 0];
  assign _zz_3640 = _zz_3641;
  assign _zz_3641 = ($signed(_zz_3642) >>> _zz_189);
  assign _zz_3642 = _zz_3643;
  assign _zz_3643 = ($signed(_zz_3645) - $signed(_zz_186));
  assign _zz_3644 = ({9'd0,data_mid_1_9_real} <<< 9);
  assign _zz_3645 = {{9{_zz_3644[26]}}, _zz_3644};
  assign _zz_3646 = fixTo_224_dout;
  assign _zz_3647 = _zz_3648[35 : 0];
  assign _zz_3648 = _zz_3649;
  assign _zz_3649 = ($signed(_zz_3650) >>> _zz_189);
  assign _zz_3650 = _zz_3651;
  assign _zz_3651 = ($signed(_zz_3653) - $signed(_zz_187));
  assign _zz_3652 = ({9'd0,data_mid_1_9_imag} <<< 9);
  assign _zz_3653 = {{9{_zz_3652[26]}}, _zz_3652};
  assign _zz_3654 = fixTo_225_dout;
  assign _zz_3655 = _zz_3656[35 : 0];
  assign _zz_3656 = _zz_3657;
  assign _zz_3657 = ($signed(_zz_3658) >>> _zz_190);
  assign _zz_3658 = _zz_3659;
  assign _zz_3659 = ($signed(_zz_3661) + $signed(_zz_186));
  assign _zz_3660 = ({9'd0,data_mid_1_9_real} <<< 9);
  assign _zz_3661 = {{9{_zz_3660[26]}}, _zz_3660};
  assign _zz_3662 = fixTo_226_dout;
  assign _zz_3663 = _zz_3664[35 : 0];
  assign _zz_3664 = _zz_3665;
  assign _zz_3665 = ($signed(_zz_3666) >>> _zz_190);
  assign _zz_3666 = _zz_3667;
  assign _zz_3667 = ($signed(_zz_3669) + $signed(_zz_187));
  assign _zz_3668 = ({9'd0,data_mid_1_9_imag} <<< 9);
  assign _zz_3669 = {{9{_zz_3668[26]}}, _zz_3668};
  assign _zz_3670 = fixTo_227_dout;
  assign _zz_3671 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_3672 = ($signed(_zz_193) - $signed(_zz_3673));
  assign _zz_3673 = ($signed(_zz_3674) * $signed(twiddle_factor_table_1_imag));
  assign _zz_3674 = ($signed(data_mid_1_14_real) + $signed(data_mid_1_14_imag));
  assign _zz_3675 = fixTo_228_dout;
  assign _zz_3676 = ($signed(_zz_193) + $signed(_zz_3677));
  assign _zz_3677 = ($signed(_zz_3678) * $signed(twiddle_factor_table_1_real));
  assign _zz_3678 = ($signed(data_mid_1_14_imag) - $signed(data_mid_1_14_real));
  assign _zz_3679 = fixTo_229_dout;
  assign _zz_3680 = _zz_3681[35 : 0];
  assign _zz_3681 = _zz_3682;
  assign _zz_3682 = ($signed(_zz_3683) >>> _zz_194);
  assign _zz_3683 = _zz_3684;
  assign _zz_3684 = ($signed(_zz_3686) - $signed(_zz_191));
  assign _zz_3685 = ({9'd0,data_mid_1_12_real} <<< 9);
  assign _zz_3686 = {{9{_zz_3685[26]}}, _zz_3685};
  assign _zz_3687 = fixTo_230_dout;
  assign _zz_3688 = _zz_3689[35 : 0];
  assign _zz_3689 = _zz_3690;
  assign _zz_3690 = ($signed(_zz_3691) >>> _zz_194);
  assign _zz_3691 = _zz_3692;
  assign _zz_3692 = ($signed(_zz_3694) - $signed(_zz_192));
  assign _zz_3693 = ({9'd0,data_mid_1_12_imag} <<< 9);
  assign _zz_3694 = {{9{_zz_3693[26]}}, _zz_3693};
  assign _zz_3695 = fixTo_231_dout;
  assign _zz_3696 = _zz_3697[35 : 0];
  assign _zz_3697 = _zz_3698;
  assign _zz_3698 = ($signed(_zz_3699) >>> _zz_195);
  assign _zz_3699 = _zz_3700;
  assign _zz_3700 = ($signed(_zz_3702) + $signed(_zz_191));
  assign _zz_3701 = ({9'd0,data_mid_1_12_real} <<< 9);
  assign _zz_3702 = {{9{_zz_3701[26]}}, _zz_3701};
  assign _zz_3703 = fixTo_232_dout;
  assign _zz_3704 = _zz_3705[35 : 0];
  assign _zz_3705 = _zz_3706;
  assign _zz_3706 = ($signed(_zz_3707) >>> _zz_195);
  assign _zz_3707 = _zz_3708;
  assign _zz_3708 = ($signed(_zz_3710) + $signed(_zz_192));
  assign _zz_3709 = ({9'd0,data_mid_1_12_imag} <<< 9);
  assign _zz_3710 = {{9{_zz_3709[26]}}, _zz_3709};
  assign _zz_3711 = fixTo_233_dout;
  assign _zz_3712 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_3713 = ($signed(_zz_198) - $signed(_zz_3714));
  assign _zz_3714 = ($signed(_zz_3715) * $signed(twiddle_factor_table_2_imag));
  assign _zz_3715 = ($signed(data_mid_1_15_real) + $signed(data_mid_1_15_imag));
  assign _zz_3716 = fixTo_234_dout;
  assign _zz_3717 = ($signed(_zz_198) + $signed(_zz_3718));
  assign _zz_3718 = ($signed(_zz_3719) * $signed(twiddle_factor_table_2_real));
  assign _zz_3719 = ($signed(data_mid_1_15_imag) - $signed(data_mid_1_15_real));
  assign _zz_3720 = fixTo_235_dout;
  assign _zz_3721 = _zz_3722[35 : 0];
  assign _zz_3722 = _zz_3723;
  assign _zz_3723 = ($signed(_zz_3724) >>> _zz_199);
  assign _zz_3724 = _zz_3725;
  assign _zz_3725 = ($signed(_zz_3727) - $signed(_zz_196));
  assign _zz_3726 = ({9'd0,data_mid_1_13_real} <<< 9);
  assign _zz_3727 = {{9{_zz_3726[26]}}, _zz_3726};
  assign _zz_3728 = fixTo_236_dout;
  assign _zz_3729 = _zz_3730[35 : 0];
  assign _zz_3730 = _zz_3731;
  assign _zz_3731 = ($signed(_zz_3732) >>> _zz_199);
  assign _zz_3732 = _zz_3733;
  assign _zz_3733 = ($signed(_zz_3735) - $signed(_zz_197));
  assign _zz_3734 = ({9'd0,data_mid_1_13_imag} <<< 9);
  assign _zz_3735 = {{9{_zz_3734[26]}}, _zz_3734};
  assign _zz_3736 = fixTo_237_dout;
  assign _zz_3737 = _zz_3738[35 : 0];
  assign _zz_3738 = _zz_3739;
  assign _zz_3739 = ($signed(_zz_3740) >>> _zz_200);
  assign _zz_3740 = _zz_3741;
  assign _zz_3741 = ($signed(_zz_3743) + $signed(_zz_196));
  assign _zz_3742 = ({9'd0,data_mid_1_13_real} <<< 9);
  assign _zz_3743 = {{9{_zz_3742[26]}}, _zz_3742};
  assign _zz_3744 = fixTo_238_dout;
  assign _zz_3745 = _zz_3746[35 : 0];
  assign _zz_3746 = _zz_3747;
  assign _zz_3747 = ($signed(_zz_3748) >>> _zz_200);
  assign _zz_3748 = _zz_3749;
  assign _zz_3749 = ($signed(_zz_3751) + $signed(_zz_197));
  assign _zz_3750 = ({9'd0,data_mid_1_13_imag} <<< 9);
  assign _zz_3751 = {{9{_zz_3750[26]}}, _zz_3750};
  assign _zz_3752 = fixTo_239_dout;
  assign _zz_3753 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_3754 = ($signed(_zz_203) - $signed(_zz_3755));
  assign _zz_3755 = ($signed(_zz_3756) * $signed(twiddle_factor_table_1_imag));
  assign _zz_3756 = ($signed(data_mid_1_18_real) + $signed(data_mid_1_18_imag));
  assign _zz_3757 = fixTo_240_dout;
  assign _zz_3758 = ($signed(_zz_203) + $signed(_zz_3759));
  assign _zz_3759 = ($signed(_zz_3760) * $signed(twiddle_factor_table_1_real));
  assign _zz_3760 = ($signed(data_mid_1_18_imag) - $signed(data_mid_1_18_real));
  assign _zz_3761 = fixTo_241_dout;
  assign _zz_3762 = _zz_3763[35 : 0];
  assign _zz_3763 = _zz_3764;
  assign _zz_3764 = ($signed(_zz_3765) >>> _zz_204);
  assign _zz_3765 = _zz_3766;
  assign _zz_3766 = ($signed(_zz_3768) - $signed(_zz_201));
  assign _zz_3767 = ({9'd0,data_mid_1_16_real} <<< 9);
  assign _zz_3768 = {{9{_zz_3767[26]}}, _zz_3767};
  assign _zz_3769 = fixTo_242_dout;
  assign _zz_3770 = _zz_3771[35 : 0];
  assign _zz_3771 = _zz_3772;
  assign _zz_3772 = ($signed(_zz_3773) >>> _zz_204);
  assign _zz_3773 = _zz_3774;
  assign _zz_3774 = ($signed(_zz_3776) - $signed(_zz_202));
  assign _zz_3775 = ({9'd0,data_mid_1_16_imag} <<< 9);
  assign _zz_3776 = {{9{_zz_3775[26]}}, _zz_3775};
  assign _zz_3777 = fixTo_243_dout;
  assign _zz_3778 = _zz_3779[35 : 0];
  assign _zz_3779 = _zz_3780;
  assign _zz_3780 = ($signed(_zz_3781) >>> _zz_205);
  assign _zz_3781 = _zz_3782;
  assign _zz_3782 = ($signed(_zz_3784) + $signed(_zz_201));
  assign _zz_3783 = ({9'd0,data_mid_1_16_real} <<< 9);
  assign _zz_3784 = {{9{_zz_3783[26]}}, _zz_3783};
  assign _zz_3785 = fixTo_244_dout;
  assign _zz_3786 = _zz_3787[35 : 0];
  assign _zz_3787 = _zz_3788;
  assign _zz_3788 = ($signed(_zz_3789) >>> _zz_205);
  assign _zz_3789 = _zz_3790;
  assign _zz_3790 = ($signed(_zz_3792) + $signed(_zz_202));
  assign _zz_3791 = ({9'd0,data_mid_1_16_imag} <<< 9);
  assign _zz_3792 = {{9{_zz_3791[26]}}, _zz_3791};
  assign _zz_3793 = fixTo_245_dout;
  assign _zz_3794 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_3795 = ($signed(_zz_208) - $signed(_zz_3796));
  assign _zz_3796 = ($signed(_zz_3797) * $signed(twiddle_factor_table_2_imag));
  assign _zz_3797 = ($signed(data_mid_1_19_real) + $signed(data_mid_1_19_imag));
  assign _zz_3798 = fixTo_246_dout;
  assign _zz_3799 = ($signed(_zz_208) + $signed(_zz_3800));
  assign _zz_3800 = ($signed(_zz_3801) * $signed(twiddle_factor_table_2_real));
  assign _zz_3801 = ($signed(data_mid_1_19_imag) - $signed(data_mid_1_19_real));
  assign _zz_3802 = fixTo_247_dout;
  assign _zz_3803 = _zz_3804[35 : 0];
  assign _zz_3804 = _zz_3805;
  assign _zz_3805 = ($signed(_zz_3806) >>> _zz_209);
  assign _zz_3806 = _zz_3807;
  assign _zz_3807 = ($signed(_zz_3809) - $signed(_zz_206));
  assign _zz_3808 = ({9'd0,data_mid_1_17_real} <<< 9);
  assign _zz_3809 = {{9{_zz_3808[26]}}, _zz_3808};
  assign _zz_3810 = fixTo_248_dout;
  assign _zz_3811 = _zz_3812[35 : 0];
  assign _zz_3812 = _zz_3813;
  assign _zz_3813 = ($signed(_zz_3814) >>> _zz_209);
  assign _zz_3814 = _zz_3815;
  assign _zz_3815 = ($signed(_zz_3817) - $signed(_zz_207));
  assign _zz_3816 = ({9'd0,data_mid_1_17_imag} <<< 9);
  assign _zz_3817 = {{9{_zz_3816[26]}}, _zz_3816};
  assign _zz_3818 = fixTo_249_dout;
  assign _zz_3819 = _zz_3820[35 : 0];
  assign _zz_3820 = _zz_3821;
  assign _zz_3821 = ($signed(_zz_3822) >>> _zz_210);
  assign _zz_3822 = _zz_3823;
  assign _zz_3823 = ($signed(_zz_3825) + $signed(_zz_206));
  assign _zz_3824 = ({9'd0,data_mid_1_17_real} <<< 9);
  assign _zz_3825 = {{9{_zz_3824[26]}}, _zz_3824};
  assign _zz_3826 = fixTo_250_dout;
  assign _zz_3827 = _zz_3828[35 : 0];
  assign _zz_3828 = _zz_3829;
  assign _zz_3829 = ($signed(_zz_3830) >>> _zz_210);
  assign _zz_3830 = _zz_3831;
  assign _zz_3831 = ($signed(_zz_3833) + $signed(_zz_207));
  assign _zz_3832 = ({9'd0,data_mid_1_17_imag} <<< 9);
  assign _zz_3833 = {{9{_zz_3832[26]}}, _zz_3832};
  assign _zz_3834 = fixTo_251_dout;
  assign _zz_3835 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_3836 = ($signed(_zz_213) - $signed(_zz_3837));
  assign _zz_3837 = ($signed(_zz_3838) * $signed(twiddle_factor_table_1_imag));
  assign _zz_3838 = ($signed(data_mid_1_22_real) + $signed(data_mid_1_22_imag));
  assign _zz_3839 = fixTo_252_dout;
  assign _zz_3840 = ($signed(_zz_213) + $signed(_zz_3841));
  assign _zz_3841 = ($signed(_zz_3842) * $signed(twiddle_factor_table_1_real));
  assign _zz_3842 = ($signed(data_mid_1_22_imag) - $signed(data_mid_1_22_real));
  assign _zz_3843 = fixTo_253_dout;
  assign _zz_3844 = _zz_3845[35 : 0];
  assign _zz_3845 = _zz_3846;
  assign _zz_3846 = ($signed(_zz_3847) >>> _zz_214);
  assign _zz_3847 = _zz_3848;
  assign _zz_3848 = ($signed(_zz_3850) - $signed(_zz_211));
  assign _zz_3849 = ({9'd0,data_mid_1_20_real} <<< 9);
  assign _zz_3850 = {{9{_zz_3849[26]}}, _zz_3849};
  assign _zz_3851 = fixTo_254_dout;
  assign _zz_3852 = _zz_3853[35 : 0];
  assign _zz_3853 = _zz_3854;
  assign _zz_3854 = ($signed(_zz_3855) >>> _zz_214);
  assign _zz_3855 = _zz_3856;
  assign _zz_3856 = ($signed(_zz_3858) - $signed(_zz_212));
  assign _zz_3857 = ({9'd0,data_mid_1_20_imag} <<< 9);
  assign _zz_3858 = {{9{_zz_3857[26]}}, _zz_3857};
  assign _zz_3859 = fixTo_255_dout;
  assign _zz_3860 = _zz_3861[35 : 0];
  assign _zz_3861 = _zz_3862;
  assign _zz_3862 = ($signed(_zz_3863) >>> _zz_215);
  assign _zz_3863 = _zz_3864;
  assign _zz_3864 = ($signed(_zz_3866) + $signed(_zz_211));
  assign _zz_3865 = ({9'd0,data_mid_1_20_real} <<< 9);
  assign _zz_3866 = {{9{_zz_3865[26]}}, _zz_3865};
  assign _zz_3867 = fixTo_256_dout;
  assign _zz_3868 = _zz_3869[35 : 0];
  assign _zz_3869 = _zz_3870;
  assign _zz_3870 = ($signed(_zz_3871) >>> _zz_215);
  assign _zz_3871 = _zz_3872;
  assign _zz_3872 = ($signed(_zz_3874) + $signed(_zz_212));
  assign _zz_3873 = ({9'd0,data_mid_1_20_imag} <<< 9);
  assign _zz_3874 = {{9{_zz_3873[26]}}, _zz_3873};
  assign _zz_3875 = fixTo_257_dout;
  assign _zz_3876 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_3877 = ($signed(_zz_218) - $signed(_zz_3878));
  assign _zz_3878 = ($signed(_zz_3879) * $signed(twiddle_factor_table_2_imag));
  assign _zz_3879 = ($signed(data_mid_1_23_real) + $signed(data_mid_1_23_imag));
  assign _zz_3880 = fixTo_258_dout;
  assign _zz_3881 = ($signed(_zz_218) + $signed(_zz_3882));
  assign _zz_3882 = ($signed(_zz_3883) * $signed(twiddle_factor_table_2_real));
  assign _zz_3883 = ($signed(data_mid_1_23_imag) - $signed(data_mid_1_23_real));
  assign _zz_3884 = fixTo_259_dout;
  assign _zz_3885 = _zz_3886[35 : 0];
  assign _zz_3886 = _zz_3887;
  assign _zz_3887 = ($signed(_zz_3888) >>> _zz_219);
  assign _zz_3888 = _zz_3889;
  assign _zz_3889 = ($signed(_zz_3891) - $signed(_zz_216));
  assign _zz_3890 = ({9'd0,data_mid_1_21_real} <<< 9);
  assign _zz_3891 = {{9{_zz_3890[26]}}, _zz_3890};
  assign _zz_3892 = fixTo_260_dout;
  assign _zz_3893 = _zz_3894[35 : 0];
  assign _zz_3894 = _zz_3895;
  assign _zz_3895 = ($signed(_zz_3896) >>> _zz_219);
  assign _zz_3896 = _zz_3897;
  assign _zz_3897 = ($signed(_zz_3899) - $signed(_zz_217));
  assign _zz_3898 = ({9'd0,data_mid_1_21_imag} <<< 9);
  assign _zz_3899 = {{9{_zz_3898[26]}}, _zz_3898};
  assign _zz_3900 = fixTo_261_dout;
  assign _zz_3901 = _zz_3902[35 : 0];
  assign _zz_3902 = _zz_3903;
  assign _zz_3903 = ($signed(_zz_3904) >>> _zz_220);
  assign _zz_3904 = _zz_3905;
  assign _zz_3905 = ($signed(_zz_3907) + $signed(_zz_216));
  assign _zz_3906 = ({9'd0,data_mid_1_21_real} <<< 9);
  assign _zz_3907 = {{9{_zz_3906[26]}}, _zz_3906};
  assign _zz_3908 = fixTo_262_dout;
  assign _zz_3909 = _zz_3910[35 : 0];
  assign _zz_3910 = _zz_3911;
  assign _zz_3911 = ($signed(_zz_3912) >>> _zz_220);
  assign _zz_3912 = _zz_3913;
  assign _zz_3913 = ($signed(_zz_3915) + $signed(_zz_217));
  assign _zz_3914 = ({9'd0,data_mid_1_21_imag} <<< 9);
  assign _zz_3915 = {{9{_zz_3914[26]}}, _zz_3914};
  assign _zz_3916 = fixTo_263_dout;
  assign _zz_3917 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_3918 = ($signed(_zz_223) - $signed(_zz_3919));
  assign _zz_3919 = ($signed(_zz_3920) * $signed(twiddle_factor_table_1_imag));
  assign _zz_3920 = ($signed(data_mid_1_26_real) + $signed(data_mid_1_26_imag));
  assign _zz_3921 = fixTo_264_dout;
  assign _zz_3922 = ($signed(_zz_223) + $signed(_zz_3923));
  assign _zz_3923 = ($signed(_zz_3924) * $signed(twiddle_factor_table_1_real));
  assign _zz_3924 = ($signed(data_mid_1_26_imag) - $signed(data_mid_1_26_real));
  assign _zz_3925 = fixTo_265_dout;
  assign _zz_3926 = _zz_3927[35 : 0];
  assign _zz_3927 = _zz_3928;
  assign _zz_3928 = ($signed(_zz_3929) >>> _zz_224);
  assign _zz_3929 = _zz_3930;
  assign _zz_3930 = ($signed(_zz_3932) - $signed(_zz_221));
  assign _zz_3931 = ({9'd0,data_mid_1_24_real} <<< 9);
  assign _zz_3932 = {{9{_zz_3931[26]}}, _zz_3931};
  assign _zz_3933 = fixTo_266_dout;
  assign _zz_3934 = _zz_3935[35 : 0];
  assign _zz_3935 = _zz_3936;
  assign _zz_3936 = ($signed(_zz_3937) >>> _zz_224);
  assign _zz_3937 = _zz_3938;
  assign _zz_3938 = ($signed(_zz_3940) - $signed(_zz_222));
  assign _zz_3939 = ({9'd0,data_mid_1_24_imag} <<< 9);
  assign _zz_3940 = {{9{_zz_3939[26]}}, _zz_3939};
  assign _zz_3941 = fixTo_267_dout;
  assign _zz_3942 = _zz_3943[35 : 0];
  assign _zz_3943 = _zz_3944;
  assign _zz_3944 = ($signed(_zz_3945) >>> _zz_225);
  assign _zz_3945 = _zz_3946;
  assign _zz_3946 = ($signed(_zz_3948) + $signed(_zz_221));
  assign _zz_3947 = ({9'd0,data_mid_1_24_real} <<< 9);
  assign _zz_3948 = {{9{_zz_3947[26]}}, _zz_3947};
  assign _zz_3949 = fixTo_268_dout;
  assign _zz_3950 = _zz_3951[35 : 0];
  assign _zz_3951 = _zz_3952;
  assign _zz_3952 = ($signed(_zz_3953) >>> _zz_225);
  assign _zz_3953 = _zz_3954;
  assign _zz_3954 = ($signed(_zz_3956) + $signed(_zz_222));
  assign _zz_3955 = ({9'd0,data_mid_1_24_imag} <<< 9);
  assign _zz_3956 = {{9{_zz_3955[26]}}, _zz_3955};
  assign _zz_3957 = fixTo_269_dout;
  assign _zz_3958 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_3959 = ($signed(_zz_228) - $signed(_zz_3960));
  assign _zz_3960 = ($signed(_zz_3961) * $signed(twiddle_factor_table_2_imag));
  assign _zz_3961 = ($signed(data_mid_1_27_real) + $signed(data_mid_1_27_imag));
  assign _zz_3962 = fixTo_270_dout;
  assign _zz_3963 = ($signed(_zz_228) + $signed(_zz_3964));
  assign _zz_3964 = ($signed(_zz_3965) * $signed(twiddle_factor_table_2_real));
  assign _zz_3965 = ($signed(data_mid_1_27_imag) - $signed(data_mid_1_27_real));
  assign _zz_3966 = fixTo_271_dout;
  assign _zz_3967 = _zz_3968[35 : 0];
  assign _zz_3968 = _zz_3969;
  assign _zz_3969 = ($signed(_zz_3970) >>> _zz_229);
  assign _zz_3970 = _zz_3971;
  assign _zz_3971 = ($signed(_zz_3973) - $signed(_zz_226));
  assign _zz_3972 = ({9'd0,data_mid_1_25_real} <<< 9);
  assign _zz_3973 = {{9{_zz_3972[26]}}, _zz_3972};
  assign _zz_3974 = fixTo_272_dout;
  assign _zz_3975 = _zz_3976[35 : 0];
  assign _zz_3976 = _zz_3977;
  assign _zz_3977 = ($signed(_zz_3978) >>> _zz_229);
  assign _zz_3978 = _zz_3979;
  assign _zz_3979 = ($signed(_zz_3981) - $signed(_zz_227));
  assign _zz_3980 = ({9'd0,data_mid_1_25_imag} <<< 9);
  assign _zz_3981 = {{9{_zz_3980[26]}}, _zz_3980};
  assign _zz_3982 = fixTo_273_dout;
  assign _zz_3983 = _zz_3984[35 : 0];
  assign _zz_3984 = _zz_3985;
  assign _zz_3985 = ($signed(_zz_3986) >>> _zz_230);
  assign _zz_3986 = _zz_3987;
  assign _zz_3987 = ($signed(_zz_3989) + $signed(_zz_226));
  assign _zz_3988 = ({9'd0,data_mid_1_25_real} <<< 9);
  assign _zz_3989 = {{9{_zz_3988[26]}}, _zz_3988};
  assign _zz_3990 = fixTo_274_dout;
  assign _zz_3991 = _zz_3992[35 : 0];
  assign _zz_3992 = _zz_3993;
  assign _zz_3993 = ($signed(_zz_3994) >>> _zz_230);
  assign _zz_3994 = _zz_3995;
  assign _zz_3995 = ($signed(_zz_3997) + $signed(_zz_227));
  assign _zz_3996 = ({9'd0,data_mid_1_25_imag} <<< 9);
  assign _zz_3997 = {{9{_zz_3996[26]}}, _zz_3996};
  assign _zz_3998 = fixTo_275_dout;
  assign _zz_3999 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_4000 = ($signed(_zz_233) - $signed(_zz_4001));
  assign _zz_4001 = ($signed(_zz_4002) * $signed(twiddle_factor_table_1_imag));
  assign _zz_4002 = ($signed(data_mid_1_30_real) + $signed(data_mid_1_30_imag));
  assign _zz_4003 = fixTo_276_dout;
  assign _zz_4004 = ($signed(_zz_233) + $signed(_zz_4005));
  assign _zz_4005 = ($signed(_zz_4006) * $signed(twiddle_factor_table_1_real));
  assign _zz_4006 = ($signed(data_mid_1_30_imag) - $signed(data_mid_1_30_real));
  assign _zz_4007 = fixTo_277_dout;
  assign _zz_4008 = _zz_4009[35 : 0];
  assign _zz_4009 = _zz_4010;
  assign _zz_4010 = ($signed(_zz_4011) >>> _zz_234);
  assign _zz_4011 = _zz_4012;
  assign _zz_4012 = ($signed(_zz_4014) - $signed(_zz_231));
  assign _zz_4013 = ({9'd0,data_mid_1_28_real} <<< 9);
  assign _zz_4014 = {{9{_zz_4013[26]}}, _zz_4013};
  assign _zz_4015 = fixTo_278_dout;
  assign _zz_4016 = _zz_4017[35 : 0];
  assign _zz_4017 = _zz_4018;
  assign _zz_4018 = ($signed(_zz_4019) >>> _zz_234);
  assign _zz_4019 = _zz_4020;
  assign _zz_4020 = ($signed(_zz_4022) - $signed(_zz_232));
  assign _zz_4021 = ({9'd0,data_mid_1_28_imag} <<< 9);
  assign _zz_4022 = {{9{_zz_4021[26]}}, _zz_4021};
  assign _zz_4023 = fixTo_279_dout;
  assign _zz_4024 = _zz_4025[35 : 0];
  assign _zz_4025 = _zz_4026;
  assign _zz_4026 = ($signed(_zz_4027) >>> _zz_235);
  assign _zz_4027 = _zz_4028;
  assign _zz_4028 = ($signed(_zz_4030) + $signed(_zz_231));
  assign _zz_4029 = ({9'd0,data_mid_1_28_real} <<< 9);
  assign _zz_4030 = {{9{_zz_4029[26]}}, _zz_4029};
  assign _zz_4031 = fixTo_280_dout;
  assign _zz_4032 = _zz_4033[35 : 0];
  assign _zz_4033 = _zz_4034;
  assign _zz_4034 = ($signed(_zz_4035) >>> _zz_235);
  assign _zz_4035 = _zz_4036;
  assign _zz_4036 = ($signed(_zz_4038) + $signed(_zz_232));
  assign _zz_4037 = ({9'd0,data_mid_1_28_imag} <<< 9);
  assign _zz_4038 = {{9{_zz_4037[26]}}, _zz_4037};
  assign _zz_4039 = fixTo_281_dout;
  assign _zz_4040 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_4041 = ($signed(_zz_238) - $signed(_zz_4042));
  assign _zz_4042 = ($signed(_zz_4043) * $signed(twiddle_factor_table_2_imag));
  assign _zz_4043 = ($signed(data_mid_1_31_real) + $signed(data_mid_1_31_imag));
  assign _zz_4044 = fixTo_282_dout;
  assign _zz_4045 = ($signed(_zz_238) + $signed(_zz_4046));
  assign _zz_4046 = ($signed(_zz_4047) * $signed(twiddle_factor_table_2_real));
  assign _zz_4047 = ($signed(data_mid_1_31_imag) - $signed(data_mid_1_31_real));
  assign _zz_4048 = fixTo_283_dout;
  assign _zz_4049 = _zz_4050[35 : 0];
  assign _zz_4050 = _zz_4051;
  assign _zz_4051 = ($signed(_zz_4052) >>> _zz_239);
  assign _zz_4052 = _zz_4053;
  assign _zz_4053 = ($signed(_zz_4055) - $signed(_zz_236));
  assign _zz_4054 = ({9'd0,data_mid_1_29_real} <<< 9);
  assign _zz_4055 = {{9{_zz_4054[26]}}, _zz_4054};
  assign _zz_4056 = fixTo_284_dout;
  assign _zz_4057 = _zz_4058[35 : 0];
  assign _zz_4058 = _zz_4059;
  assign _zz_4059 = ($signed(_zz_4060) >>> _zz_239);
  assign _zz_4060 = _zz_4061;
  assign _zz_4061 = ($signed(_zz_4063) - $signed(_zz_237));
  assign _zz_4062 = ({9'd0,data_mid_1_29_imag} <<< 9);
  assign _zz_4063 = {{9{_zz_4062[26]}}, _zz_4062};
  assign _zz_4064 = fixTo_285_dout;
  assign _zz_4065 = _zz_4066[35 : 0];
  assign _zz_4066 = _zz_4067;
  assign _zz_4067 = ($signed(_zz_4068) >>> _zz_240);
  assign _zz_4068 = _zz_4069;
  assign _zz_4069 = ($signed(_zz_4071) + $signed(_zz_236));
  assign _zz_4070 = ({9'd0,data_mid_1_29_real} <<< 9);
  assign _zz_4071 = {{9{_zz_4070[26]}}, _zz_4070};
  assign _zz_4072 = fixTo_286_dout;
  assign _zz_4073 = _zz_4074[35 : 0];
  assign _zz_4074 = _zz_4075;
  assign _zz_4075 = ($signed(_zz_4076) >>> _zz_240);
  assign _zz_4076 = _zz_4077;
  assign _zz_4077 = ($signed(_zz_4079) + $signed(_zz_237));
  assign _zz_4078 = ({9'd0,data_mid_1_29_imag} <<< 9);
  assign _zz_4079 = {{9{_zz_4078[26]}}, _zz_4078};
  assign _zz_4080 = fixTo_287_dout;
  assign _zz_4081 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_4082 = ($signed(_zz_243) - $signed(_zz_4083));
  assign _zz_4083 = ($signed(_zz_4084) * $signed(twiddle_factor_table_1_imag));
  assign _zz_4084 = ($signed(data_mid_1_34_real) + $signed(data_mid_1_34_imag));
  assign _zz_4085 = fixTo_288_dout;
  assign _zz_4086 = ($signed(_zz_243) + $signed(_zz_4087));
  assign _zz_4087 = ($signed(_zz_4088) * $signed(twiddle_factor_table_1_real));
  assign _zz_4088 = ($signed(data_mid_1_34_imag) - $signed(data_mid_1_34_real));
  assign _zz_4089 = fixTo_289_dout;
  assign _zz_4090 = _zz_4091[35 : 0];
  assign _zz_4091 = _zz_4092;
  assign _zz_4092 = ($signed(_zz_4093) >>> _zz_244);
  assign _zz_4093 = _zz_4094;
  assign _zz_4094 = ($signed(_zz_4096) - $signed(_zz_241));
  assign _zz_4095 = ({9'd0,data_mid_1_32_real} <<< 9);
  assign _zz_4096 = {{9{_zz_4095[26]}}, _zz_4095};
  assign _zz_4097 = fixTo_290_dout;
  assign _zz_4098 = _zz_4099[35 : 0];
  assign _zz_4099 = _zz_4100;
  assign _zz_4100 = ($signed(_zz_4101) >>> _zz_244);
  assign _zz_4101 = _zz_4102;
  assign _zz_4102 = ($signed(_zz_4104) - $signed(_zz_242));
  assign _zz_4103 = ({9'd0,data_mid_1_32_imag} <<< 9);
  assign _zz_4104 = {{9{_zz_4103[26]}}, _zz_4103};
  assign _zz_4105 = fixTo_291_dout;
  assign _zz_4106 = _zz_4107[35 : 0];
  assign _zz_4107 = _zz_4108;
  assign _zz_4108 = ($signed(_zz_4109) >>> _zz_245);
  assign _zz_4109 = _zz_4110;
  assign _zz_4110 = ($signed(_zz_4112) + $signed(_zz_241));
  assign _zz_4111 = ({9'd0,data_mid_1_32_real} <<< 9);
  assign _zz_4112 = {{9{_zz_4111[26]}}, _zz_4111};
  assign _zz_4113 = fixTo_292_dout;
  assign _zz_4114 = _zz_4115[35 : 0];
  assign _zz_4115 = _zz_4116;
  assign _zz_4116 = ($signed(_zz_4117) >>> _zz_245);
  assign _zz_4117 = _zz_4118;
  assign _zz_4118 = ($signed(_zz_4120) + $signed(_zz_242));
  assign _zz_4119 = ({9'd0,data_mid_1_32_imag} <<< 9);
  assign _zz_4120 = {{9{_zz_4119[26]}}, _zz_4119};
  assign _zz_4121 = fixTo_293_dout;
  assign _zz_4122 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_4123 = ($signed(_zz_248) - $signed(_zz_4124));
  assign _zz_4124 = ($signed(_zz_4125) * $signed(twiddle_factor_table_2_imag));
  assign _zz_4125 = ($signed(data_mid_1_35_real) + $signed(data_mid_1_35_imag));
  assign _zz_4126 = fixTo_294_dout;
  assign _zz_4127 = ($signed(_zz_248) + $signed(_zz_4128));
  assign _zz_4128 = ($signed(_zz_4129) * $signed(twiddle_factor_table_2_real));
  assign _zz_4129 = ($signed(data_mid_1_35_imag) - $signed(data_mid_1_35_real));
  assign _zz_4130 = fixTo_295_dout;
  assign _zz_4131 = _zz_4132[35 : 0];
  assign _zz_4132 = _zz_4133;
  assign _zz_4133 = ($signed(_zz_4134) >>> _zz_249);
  assign _zz_4134 = _zz_4135;
  assign _zz_4135 = ($signed(_zz_4137) - $signed(_zz_246));
  assign _zz_4136 = ({9'd0,data_mid_1_33_real} <<< 9);
  assign _zz_4137 = {{9{_zz_4136[26]}}, _zz_4136};
  assign _zz_4138 = fixTo_296_dout;
  assign _zz_4139 = _zz_4140[35 : 0];
  assign _zz_4140 = _zz_4141;
  assign _zz_4141 = ($signed(_zz_4142) >>> _zz_249);
  assign _zz_4142 = _zz_4143;
  assign _zz_4143 = ($signed(_zz_4145) - $signed(_zz_247));
  assign _zz_4144 = ({9'd0,data_mid_1_33_imag} <<< 9);
  assign _zz_4145 = {{9{_zz_4144[26]}}, _zz_4144};
  assign _zz_4146 = fixTo_297_dout;
  assign _zz_4147 = _zz_4148[35 : 0];
  assign _zz_4148 = _zz_4149;
  assign _zz_4149 = ($signed(_zz_4150) >>> _zz_250);
  assign _zz_4150 = _zz_4151;
  assign _zz_4151 = ($signed(_zz_4153) + $signed(_zz_246));
  assign _zz_4152 = ({9'd0,data_mid_1_33_real} <<< 9);
  assign _zz_4153 = {{9{_zz_4152[26]}}, _zz_4152};
  assign _zz_4154 = fixTo_298_dout;
  assign _zz_4155 = _zz_4156[35 : 0];
  assign _zz_4156 = _zz_4157;
  assign _zz_4157 = ($signed(_zz_4158) >>> _zz_250);
  assign _zz_4158 = _zz_4159;
  assign _zz_4159 = ($signed(_zz_4161) + $signed(_zz_247));
  assign _zz_4160 = ({9'd0,data_mid_1_33_imag} <<< 9);
  assign _zz_4161 = {{9{_zz_4160[26]}}, _zz_4160};
  assign _zz_4162 = fixTo_299_dout;
  assign _zz_4163 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_4164 = ($signed(_zz_253) - $signed(_zz_4165));
  assign _zz_4165 = ($signed(_zz_4166) * $signed(twiddle_factor_table_1_imag));
  assign _zz_4166 = ($signed(data_mid_1_38_real) + $signed(data_mid_1_38_imag));
  assign _zz_4167 = fixTo_300_dout;
  assign _zz_4168 = ($signed(_zz_253) + $signed(_zz_4169));
  assign _zz_4169 = ($signed(_zz_4170) * $signed(twiddle_factor_table_1_real));
  assign _zz_4170 = ($signed(data_mid_1_38_imag) - $signed(data_mid_1_38_real));
  assign _zz_4171 = fixTo_301_dout;
  assign _zz_4172 = _zz_4173[35 : 0];
  assign _zz_4173 = _zz_4174;
  assign _zz_4174 = ($signed(_zz_4175) >>> _zz_254);
  assign _zz_4175 = _zz_4176;
  assign _zz_4176 = ($signed(_zz_4178) - $signed(_zz_251));
  assign _zz_4177 = ({9'd0,data_mid_1_36_real} <<< 9);
  assign _zz_4178 = {{9{_zz_4177[26]}}, _zz_4177};
  assign _zz_4179 = fixTo_302_dout;
  assign _zz_4180 = _zz_4181[35 : 0];
  assign _zz_4181 = _zz_4182;
  assign _zz_4182 = ($signed(_zz_4183) >>> _zz_254);
  assign _zz_4183 = _zz_4184;
  assign _zz_4184 = ($signed(_zz_4186) - $signed(_zz_252));
  assign _zz_4185 = ({9'd0,data_mid_1_36_imag} <<< 9);
  assign _zz_4186 = {{9{_zz_4185[26]}}, _zz_4185};
  assign _zz_4187 = fixTo_303_dout;
  assign _zz_4188 = _zz_4189[35 : 0];
  assign _zz_4189 = _zz_4190;
  assign _zz_4190 = ($signed(_zz_4191) >>> _zz_255);
  assign _zz_4191 = _zz_4192;
  assign _zz_4192 = ($signed(_zz_4194) + $signed(_zz_251));
  assign _zz_4193 = ({9'd0,data_mid_1_36_real} <<< 9);
  assign _zz_4194 = {{9{_zz_4193[26]}}, _zz_4193};
  assign _zz_4195 = fixTo_304_dout;
  assign _zz_4196 = _zz_4197[35 : 0];
  assign _zz_4197 = _zz_4198;
  assign _zz_4198 = ($signed(_zz_4199) >>> _zz_255);
  assign _zz_4199 = _zz_4200;
  assign _zz_4200 = ($signed(_zz_4202) + $signed(_zz_252));
  assign _zz_4201 = ({9'd0,data_mid_1_36_imag} <<< 9);
  assign _zz_4202 = {{9{_zz_4201[26]}}, _zz_4201};
  assign _zz_4203 = fixTo_305_dout;
  assign _zz_4204 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_4205 = ($signed(_zz_258) - $signed(_zz_4206));
  assign _zz_4206 = ($signed(_zz_4207) * $signed(twiddle_factor_table_2_imag));
  assign _zz_4207 = ($signed(data_mid_1_39_real) + $signed(data_mid_1_39_imag));
  assign _zz_4208 = fixTo_306_dout;
  assign _zz_4209 = ($signed(_zz_258) + $signed(_zz_4210));
  assign _zz_4210 = ($signed(_zz_4211) * $signed(twiddle_factor_table_2_real));
  assign _zz_4211 = ($signed(data_mid_1_39_imag) - $signed(data_mid_1_39_real));
  assign _zz_4212 = fixTo_307_dout;
  assign _zz_4213 = _zz_4214[35 : 0];
  assign _zz_4214 = _zz_4215;
  assign _zz_4215 = ($signed(_zz_4216) >>> _zz_259);
  assign _zz_4216 = _zz_4217;
  assign _zz_4217 = ($signed(_zz_4219) - $signed(_zz_256));
  assign _zz_4218 = ({9'd0,data_mid_1_37_real} <<< 9);
  assign _zz_4219 = {{9{_zz_4218[26]}}, _zz_4218};
  assign _zz_4220 = fixTo_308_dout;
  assign _zz_4221 = _zz_4222[35 : 0];
  assign _zz_4222 = _zz_4223;
  assign _zz_4223 = ($signed(_zz_4224) >>> _zz_259);
  assign _zz_4224 = _zz_4225;
  assign _zz_4225 = ($signed(_zz_4227) - $signed(_zz_257));
  assign _zz_4226 = ({9'd0,data_mid_1_37_imag} <<< 9);
  assign _zz_4227 = {{9{_zz_4226[26]}}, _zz_4226};
  assign _zz_4228 = fixTo_309_dout;
  assign _zz_4229 = _zz_4230[35 : 0];
  assign _zz_4230 = _zz_4231;
  assign _zz_4231 = ($signed(_zz_4232) >>> _zz_260);
  assign _zz_4232 = _zz_4233;
  assign _zz_4233 = ($signed(_zz_4235) + $signed(_zz_256));
  assign _zz_4234 = ({9'd0,data_mid_1_37_real} <<< 9);
  assign _zz_4235 = {{9{_zz_4234[26]}}, _zz_4234};
  assign _zz_4236 = fixTo_310_dout;
  assign _zz_4237 = _zz_4238[35 : 0];
  assign _zz_4238 = _zz_4239;
  assign _zz_4239 = ($signed(_zz_4240) >>> _zz_260);
  assign _zz_4240 = _zz_4241;
  assign _zz_4241 = ($signed(_zz_4243) + $signed(_zz_257));
  assign _zz_4242 = ({9'd0,data_mid_1_37_imag} <<< 9);
  assign _zz_4243 = {{9{_zz_4242[26]}}, _zz_4242};
  assign _zz_4244 = fixTo_311_dout;
  assign _zz_4245 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_4246 = ($signed(_zz_263) - $signed(_zz_4247));
  assign _zz_4247 = ($signed(_zz_4248) * $signed(twiddle_factor_table_1_imag));
  assign _zz_4248 = ($signed(data_mid_1_42_real) + $signed(data_mid_1_42_imag));
  assign _zz_4249 = fixTo_312_dout;
  assign _zz_4250 = ($signed(_zz_263) + $signed(_zz_4251));
  assign _zz_4251 = ($signed(_zz_4252) * $signed(twiddle_factor_table_1_real));
  assign _zz_4252 = ($signed(data_mid_1_42_imag) - $signed(data_mid_1_42_real));
  assign _zz_4253 = fixTo_313_dout;
  assign _zz_4254 = _zz_4255[35 : 0];
  assign _zz_4255 = _zz_4256;
  assign _zz_4256 = ($signed(_zz_4257) >>> _zz_264);
  assign _zz_4257 = _zz_4258;
  assign _zz_4258 = ($signed(_zz_4260) - $signed(_zz_261));
  assign _zz_4259 = ({9'd0,data_mid_1_40_real} <<< 9);
  assign _zz_4260 = {{9{_zz_4259[26]}}, _zz_4259};
  assign _zz_4261 = fixTo_314_dout;
  assign _zz_4262 = _zz_4263[35 : 0];
  assign _zz_4263 = _zz_4264;
  assign _zz_4264 = ($signed(_zz_4265) >>> _zz_264);
  assign _zz_4265 = _zz_4266;
  assign _zz_4266 = ($signed(_zz_4268) - $signed(_zz_262));
  assign _zz_4267 = ({9'd0,data_mid_1_40_imag} <<< 9);
  assign _zz_4268 = {{9{_zz_4267[26]}}, _zz_4267};
  assign _zz_4269 = fixTo_315_dout;
  assign _zz_4270 = _zz_4271[35 : 0];
  assign _zz_4271 = _zz_4272;
  assign _zz_4272 = ($signed(_zz_4273) >>> _zz_265);
  assign _zz_4273 = _zz_4274;
  assign _zz_4274 = ($signed(_zz_4276) + $signed(_zz_261));
  assign _zz_4275 = ({9'd0,data_mid_1_40_real} <<< 9);
  assign _zz_4276 = {{9{_zz_4275[26]}}, _zz_4275};
  assign _zz_4277 = fixTo_316_dout;
  assign _zz_4278 = _zz_4279[35 : 0];
  assign _zz_4279 = _zz_4280;
  assign _zz_4280 = ($signed(_zz_4281) >>> _zz_265);
  assign _zz_4281 = _zz_4282;
  assign _zz_4282 = ($signed(_zz_4284) + $signed(_zz_262));
  assign _zz_4283 = ({9'd0,data_mid_1_40_imag} <<< 9);
  assign _zz_4284 = {{9{_zz_4283[26]}}, _zz_4283};
  assign _zz_4285 = fixTo_317_dout;
  assign _zz_4286 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_4287 = ($signed(_zz_268) - $signed(_zz_4288));
  assign _zz_4288 = ($signed(_zz_4289) * $signed(twiddle_factor_table_2_imag));
  assign _zz_4289 = ($signed(data_mid_1_43_real) + $signed(data_mid_1_43_imag));
  assign _zz_4290 = fixTo_318_dout;
  assign _zz_4291 = ($signed(_zz_268) + $signed(_zz_4292));
  assign _zz_4292 = ($signed(_zz_4293) * $signed(twiddle_factor_table_2_real));
  assign _zz_4293 = ($signed(data_mid_1_43_imag) - $signed(data_mid_1_43_real));
  assign _zz_4294 = fixTo_319_dout;
  assign _zz_4295 = _zz_4296[35 : 0];
  assign _zz_4296 = _zz_4297;
  assign _zz_4297 = ($signed(_zz_4298) >>> _zz_269);
  assign _zz_4298 = _zz_4299;
  assign _zz_4299 = ($signed(_zz_4301) - $signed(_zz_266));
  assign _zz_4300 = ({9'd0,data_mid_1_41_real} <<< 9);
  assign _zz_4301 = {{9{_zz_4300[26]}}, _zz_4300};
  assign _zz_4302 = fixTo_320_dout;
  assign _zz_4303 = _zz_4304[35 : 0];
  assign _zz_4304 = _zz_4305;
  assign _zz_4305 = ($signed(_zz_4306) >>> _zz_269);
  assign _zz_4306 = _zz_4307;
  assign _zz_4307 = ($signed(_zz_4309) - $signed(_zz_267));
  assign _zz_4308 = ({9'd0,data_mid_1_41_imag} <<< 9);
  assign _zz_4309 = {{9{_zz_4308[26]}}, _zz_4308};
  assign _zz_4310 = fixTo_321_dout;
  assign _zz_4311 = _zz_4312[35 : 0];
  assign _zz_4312 = _zz_4313;
  assign _zz_4313 = ($signed(_zz_4314) >>> _zz_270);
  assign _zz_4314 = _zz_4315;
  assign _zz_4315 = ($signed(_zz_4317) + $signed(_zz_266));
  assign _zz_4316 = ({9'd0,data_mid_1_41_real} <<< 9);
  assign _zz_4317 = {{9{_zz_4316[26]}}, _zz_4316};
  assign _zz_4318 = fixTo_322_dout;
  assign _zz_4319 = _zz_4320[35 : 0];
  assign _zz_4320 = _zz_4321;
  assign _zz_4321 = ($signed(_zz_4322) >>> _zz_270);
  assign _zz_4322 = _zz_4323;
  assign _zz_4323 = ($signed(_zz_4325) + $signed(_zz_267));
  assign _zz_4324 = ({9'd0,data_mid_1_41_imag} <<< 9);
  assign _zz_4325 = {{9{_zz_4324[26]}}, _zz_4324};
  assign _zz_4326 = fixTo_323_dout;
  assign _zz_4327 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_4328 = ($signed(_zz_273) - $signed(_zz_4329));
  assign _zz_4329 = ($signed(_zz_4330) * $signed(twiddle_factor_table_1_imag));
  assign _zz_4330 = ($signed(data_mid_1_46_real) + $signed(data_mid_1_46_imag));
  assign _zz_4331 = fixTo_324_dout;
  assign _zz_4332 = ($signed(_zz_273) + $signed(_zz_4333));
  assign _zz_4333 = ($signed(_zz_4334) * $signed(twiddle_factor_table_1_real));
  assign _zz_4334 = ($signed(data_mid_1_46_imag) - $signed(data_mid_1_46_real));
  assign _zz_4335 = fixTo_325_dout;
  assign _zz_4336 = _zz_4337[35 : 0];
  assign _zz_4337 = _zz_4338;
  assign _zz_4338 = ($signed(_zz_4339) >>> _zz_274);
  assign _zz_4339 = _zz_4340;
  assign _zz_4340 = ($signed(_zz_4342) - $signed(_zz_271));
  assign _zz_4341 = ({9'd0,data_mid_1_44_real} <<< 9);
  assign _zz_4342 = {{9{_zz_4341[26]}}, _zz_4341};
  assign _zz_4343 = fixTo_326_dout;
  assign _zz_4344 = _zz_4345[35 : 0];
  assign _zz_4345 = _zz_4346;
  assign _zz_4346 = ($signed(_zz_4347) >>> _zz_274);
  assign _zz_4347 = _zz_4348;
  assign _zz_4348 = ($signed(_zz_4350) - $signed(_zz_272));
  assign _zz_4349 = ({9'd0,data_mid_1_44_imag} <<< 9);
  assign _zz_4350 = {{9{_zz_4349[26]}}, _zz_4349};
  assign _zz_4351 = fixTo_327_dout;
  assign _zz_4352 = _zz_4353[35 : 0];
  assign _zz_4353 = _zz_4354;
  assign _zz_4354 = ($signed(_zz_4355) >>> _zz_275);
  assign _zz_4355 = _zz_4356;
  assign _zz_4356 = ($signed(_zz_4358) + $signed(_zz_271));
  assign _zz_4357 = ({9'd0,data_mid_1_44_real} <<< 9);
  assign _zz_4358 = {{9{_zz_4357[26]}}, _zz_4357};
  assign _zz_4359 = fixTo_328_dout;
  assign _zz_4360 = _zz_4361[35 : 0];
  assign _zz_4361 = _zz_4362;
  assign _zz_4362 = ($signed(_zz_4363) >>> _zz_275);
  assign _zz_4363 = _zz_4364;
  assign _zz_4364 = ($signed(_zz_4366) + $signed(_zz_272));
  assign _zz_4365 = ({9'd0,data_mid_1_44_imag} <<< 9);
  assign _zz_4366 = {{9{_zz_4365[26]}}, _zz_4365};
  assign _zz_4367 = fixTo_329_dout;
  assign _zz_4368 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_4369 = ($signed(_zz_278) - $signed(_zz_4370));
  assign _zz_4370 = ($signed(_zz_4371) * $signed(twiddle_factor_table_2_imag));
  assign _zz_4371 = ($signed(data_mid_1_47_real) + $signed(data_mid_1_47_imag));
  assign _zz_4372 = fixTo_330_dout;
  assign _zz_4373 = ($signed(_zz_278) + $signed(_zz_4374));
  assign _zz_4374 = ($signed(_zz_4375) * $signed(twiddle_factor_table_2_real));
  assign _zz_4375 = ($signed(data_mid_1_47_imag) - $signed(data_mid_1_47_real));
  assign _zz_4376 = fixTo_331_dout;
  assign _zz_4377 = _zz_4378[35 : 0];
  assign _zz_4378 = _zz_4379;
  assign _zz_4379 = ($signed(_zz_4380) >>> _zz_279);
  assign _zz_4380 = _zz_4381;
  assign _zz_4381 = ($signed(_zz_4383) - $signed(_zz_276));
  assign _zz_4382 = ({9'd0,data_mid_1_45_real} <<< 9);
  assign _zz_4383 = {{9{_zz_4382[26]}}, _zz_4382};
  assign _zz_4384 = fixTo_332_dout;
  assign _zz_4385 = _zz_4386[35 : 0];
  assign _zz_4386 = _zz_4387;
  assign _zz_4387 = ($signed(_zz_4388) >>> _zz_279);
  assign _zz_4388 = _zz_4389;
  assign _zz_4389 = ($signed(_zz_4391) - $signed(_zz_277));
  assign _zz_4390 = ({9'd0,data_mid_1_45_imag} <<< 9);
  assign _zz_4391 = {{9{_zz_4390[26]}}, _zz_4390};
  assign _zz_4392 = fixTo_333_dout;
  assign _zz_4393 = _zz_4394[35 : 0];
  assign _zz_4394 = _zz_4395;
  assign _zz_4395 = ($signed(_zz_4396) >>> _zz_280);
  assign _zz_4396 = _zz_4397;
  assign _zz_4397 = ($signed(_zz_4399) + $signed(_zz_276));
  assign _zz_4398 = ({9'd0,data_mid_1_45_real} <<< 9);
  assign _zz_4399 = {{9{_zz_4398[26]}}, _zz_4398};
  assign _zz_4400 = fixTo_334_dout;
  assign _zz_4401 = _zz_4402[35 : 0];
  assign _zz_4402 = _zz_4403;
  assign _zz_4403 = ($signed(_zz_4404) >>> _zz_280);
  assign _zz_4404 = _zz_4405;
  assign _zz_4405 = ($signed(_zz_4407) + $signed(_zz_277));
  assign _zz_4406 = ({9'd0,data_mid_1_45_imag} <<< 9);
  assign _zz_4407 = {{9{_zz_4406[26]}}, _zz_4406};
  assign _zz_4408 = fixTo_335_dout;
  assign _zz_4409 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_4410 = ($signed(_zz_283) - $signed(_zz_4411));
  assign _zz_4411 = ($signed(_zz_4412) * $signed(twiddle_factor_table_1_imag));
  assign _zz_4412 = ($signed(data_mid_1_50_real) + $signed(data_mid_1_50_imag));
  assign _zz_4413 = fixTo_336_dout;
  assign _zz_4414 = ($signed(_zz_283) + $signed(_zz_4415));
  assign _zz_4415 = ($signed(_zz_4416) * $signed(twiddle_factor_table_1_real));
  assign _zz_4416 = ($signed(data_mid_1_50_imag) - $signed(data_mid_1_50_real));
  assign _zz_4417 = fixTo_337_dout;
  assign _zz_4418 = _zz_4419[35 : 0];
  assign _zz_4419 = _zz_4420;
  assign _zz_4420 = ($signed(_zz_4421) >>> _zz_284);
  assign _zz_4421 = _zz_4422;
  assign _zz_4422 = ($signed(_zz_4424) - $signed(_zz_281));
  assign _zz_4423 = ({9'd0,data_mid_1_48_real} <<< 9);
  assign _zz_4424 = {{9{_zz_4423[26]}}, _zz_4423};
  assign _zz_4425 = fixTo_338_dout;
  assign _zz_4426 = _zz_4427[35 : 0];
  assign _zz_4427 = _zz_4428;
  assign _zz_4428 = ($signed(_zz_4429) >>> _zz_284);
  assign _zz_4429 = _zz_4430;
  assign _zz_4430 = ($signed(_zz_4432) - $signed(_zz_282));
  assign _zz_4431 = ({9'd0,data_mid_1_48_imag} <<< 9);
  assign _zz_4432 = {{9{_zz_4431[26]}}, _zz_4431};
  assign _zz_4433 = fixTo_339_dout;
  assign _zz_4434 = _zz_4435[35 : 0];
  assign _zz_4435 = _zz_4436;
  assign _zz_4436 = ($signed(_zz_4437) >>> _zz_285);
  assign _zz_4437 = _zz_4438;
  assign _zz_4438 = ($signed(_zz_4440) + $signed(_zz_281));
  assign _zz_4439 = ({9'd0,data_mid_1_48_real} <<< 9);
  assign _zz_4440 = {{9{_zz_4439[26]}}, _zz_4439};
  assign _zz_4441 = fixTo_340_dout;
  assign _zz_4442 = _zz_4443[35 : 0];
  assign _zz_4443 = _zz_4444;
  assign _zz_4444 = ($signed(_zz_4445) >>> _zz_285);
  assign _zz_4445 = _zz_4446;
  assign _zz_4446 = ($signed(_zz_4448) + $signed(_zz_282));
  assign _zz_4447 = ({9'd0,data_mid_1_48_imag} <<< 9);
  assign _zz_4448 = {{9{_zz_4447[26]}}, _zz_4447};
  assign _zz_4449 = fixTo_341_dout;
  assign _zz_4450 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_4451 = ($signed(_zz_288) - $signed(_zz_4452));
  assign _zz_4452 = ($signed(_zz_4453) * $signed(twiddle_factor_table_2_imag));
  assign _zz_4453 = ($signed(data_mid_1_51_real) + $signed(data_mid_1_51_imag));
  assign _zz_4454 = fixTo_342_dout;
  assign _zz_4455 = ($signed(_zz_288) + $signed(_zz_4456));
  assign _zz_4456 = ($signed(_zz_4457) * $signed(twiddle_factor_table_2_real));
  assign _zz_4457 = ($signed(data_mid_1_51_imag) - $signed(data_mid_1_51_real));
  assign _zz_4458 = fixTo_343_dout;
  assign _zz_4459 = _zz_4460[35 : 0];
  assign _zz_4460 = _zz_4461;
  assign _zz_4461 = ($signed(_zz_4462) >>> _zz_289);
  assign _zz_4462 = _zz_4463;
  assign _zz_4463 = ($signed(_zz_4465) - $signed(_zz_286));
  assign _zz_4464 = ({9'd0,data_mid_1_49_real} <<< 9);
  assign _zz_4465 = {{9{_zz_4464[26]}}, _zz_4464};
  assign _zz_4466 = fixTo_344_dout;
  assign _zz_4467 = _zz_4468[35 : 0];
  assign _zz_4468 = _zz_4469;
  assign _zz_4469 = ($signed(_zz_4470) >>> _zz_289);
  assign _zz_4470 = _zz_4471;
  assign _zz_4471 = ($signed(_zz_4473) - $signed(_zz_287));
  assign _zz_4472 = ({9'd0,data_mid_1_49_imag} <<< 9);
  assign _zz_4473 = {{9{_zz_4472[26]}}, _zz_4472};
  assign _zz_4474 = fixTo_345_dout;
  assign _zz_4475 = _zz_4476[35 : 0];
  assign _zz_4476 = _zz_4477;
  assign _zz_4477 = ($signed(_zz_4478) >>> _zz_290);
  assign _zz_4478 = _zz_4479;
  assign _zz_4479 = ($signed(_zz_4481) + $signed(_zz_286));
  assign _zz_4480 = ({9'd0,data_mid_1_49_real} <<< 9);
  assign _zz_4481 = {{9{_zz_4480[26]}}, _zz_4480};
  assign _zz_4482 = fixTo_346_dout;
  assign _zz_4483 = _zz_4484[35 : 0];
  assign _zz_4484 = _zz_4485;
  assign _zz_4485 = ($signed(_zz_4486) >>> _zz_290);
  assign _zz_4486 = _zz_4487;
  assign _zz_4487 = ($signed(_zz_4489) + $signed(_zz_287));
  assign _zz_4488 = ({9'd0,data_mid_1_49_imag} <<< 9);
  assign _zz_4489 = {{9{_zz_4488[26]}}, _zz_4488};
  assign _zz_4490 = fixTo_347_dout;
  assign _zz_4491 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_4492 = ($signed(_zz_293) - $signed(_zz_4493));
  assign _zz_4493 = ($signed(_zz_4494) * $signed(twiddle_factor_table_1_imag));
  assign _zz_4494 = ($signed(data_mid_1_54_real) + $signed(data_mid_1_54_imag));
  assign _zz_4495 = fixTo_348_dout;
  assign _zz_4496 = ($signed(_zz_293) + $signed(_zz_4497));
  assign _zz_4497 = ($signed(_zz_4498) * $signed(twiddle_factor_table_1_real));
  assign _zz_4498 = ($signed(data_mid_1_54_imag) - $signed(data_mid_1_54_real));
  assign _zz_4499 = fixTo_349_dout;
  assign _zz_4500 = _zz_4501[35 : 0];
  assign _zz_4501 = _zz_4502;
  assign _zz_4502 = ($signed(_zz_4503) >>> _zz_294);
  assign _zz_4503 = _zz_4504;
  assign _zz_4504 = ($signed(_zz_4506) - $signed(_zz_291));
  assign _zz_4505 = ({9'd0,data_mid_1_52_real} <<< 9);
  assign _zz_4506 = {{9{_zz_4505[26]}}, _zz_4505};
  assign _zz_4507 = fixTo_350_dout;
  assign _zz_4508 = _zz_4509[35 : 0];
  assign _zz_4509 = _zz_4510;
  assign _zz_4510 = ($signed(_zz_4511) >>> _zz_294);
  assign _zz_4511 = _zz_4512;
  assign _zz_4512 = ($signed(_zz_4514) - $signed(_zz_292));
  assign _zz_4513 = ({9'd0,data_mid_1_52_imag} <<< 9);
  assign _zz_4514 = {{9{_zz_4513[26]}}, _zz_4513};
  assign _zz_4515 = fixTo_351_dout;
  assign _zz_4516 = _zz_4517[35 : 0];
  assign _zz_4517 = _zz_4518;
  assign _zz_4518 = ($signed(_zz_4519) >>> _zz_295);
  assign _zz_4519 = _zz_4520;
  assign _zz_4520 = ($signed(_zz_4522) + $signed(_zz_291));
  assign _zz_4521 = ({9'd0,data_mid_1_52_real} <<< 9);
  assign _zz_4522 = {{9{_zz_4521[26]}}, _zz_4521};
  assign _zz_4523 = fixTo_352_dout;
  assign _zz_4524 = _zz_4525[35 : 0];
  assign _zz_4525 = _zz_4526;
  assign _zz_4526 = ($signed(_zz_4527) >>> _zz_295);
  assign _zz_4527 = _zz_4528;
  assign _zz_4528 = ($signed(_zz_4530) + $signed(_zz_292));
  assign _zz_4529 = ({9'd0,data_mid_1_52_imag} <<< 9);
  assign _zz_4530 = {{9{_zz_4529[26]}}, _zz_4529};
  assign _zz_4531 = fixTo_353_dout;
  assign _zz_4532 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_4533 = ($signed(_zz_298) - $signed(_zz_4534));
  assign _zz_4534 = ($signed(_zz_4535) * $signed(twiddle_factor_table_2_imag));
  assign _zz_4535 = ($signed(data_mid_1_55_real) + $signed(data_mid_1_55_imag));
  assign _zz_4536 = fixTo_354_dout;
  assign _zz_4537 = ($signed(_zz_298) + $signed(_zz_4538));
  assign _zz_4538 = ($signed(_zz_4539) * $signed(twiddle_factor_table_2_real));
  assign _zz_4539 = ($signed(data_mid_1_55_imag) - $signed(data_mid_1_55_real));
  assign _zz_4540 = fixTo_355_dout;
  assign _zz_4541 = _zz_4542[35 : 0];
  assign _zz_4542 = _zz_4543;
  assign _zz_4543 = ($signed(_zz_4544) >>> _zz_299);
  assign _zz_4544 = _zz_4545;
  assign _zz_4545 = ($signed(_zz_4547) - $signed(_zz_296));
  assign _zz_4546 = ({9'd0,data_mid_1_53_real} <<< 9);
  assign _zz_4547 = {{9{_zz_4546[26]}}, _zz_4546};
  assign _zz_4548 = fixTo_356_dout;
  assign _zz_4549 = _zz_4550[35 : 0];
  assign _zz_4550 = _zz_4551;
  assign _zz_4551 = ($signed(_zz_4552) >>> _zz_299);
  assign _zz_4552 = _zz_4553;
  assign _zz_4553 = ($signed(_zz_4555) - $signed(_zz_297));
  assign _zz_4554 = ({9'd0,data_mid_1_53_imag} <<< 9);
  assign _zz_4555 = {{9{_zz_4554[26]}}, _zz_4554};
  assign _zz_4556 = fixTo_357_dout;
  assign _zz_4557 = _zz_4558[35 : 0];
  assign _zz_4558 = _zz_4559;
  assign _zz_4559 = ($signed(_zz_4560) >>> _zz_300);
  assign _zz_4560 = _zz_4561;
  assign _zz_4561 = ($signed(_zz_4563) + $signed(_zz_296));
  assign _zz_4562 = ({9'd0,data_mid_1_53_real} <<< 9);
  assign _zz_4563 = {{9{_zz_4562[26]}}, _zz_4562};
  assign _zz_4564 = fixTo_358_dout;
  assign _zz_4565 = _zz_4566[35 : 0];
  assign _zz_4566 = _zz_4567;
  assign _zz_4567 = ($signed(_zz_4568) >>> _zz_300);
  assign _zz_4568 = _zz_4569;
  assign _zz_4569 = ($signed(_zz_4571) + $signed(_zz_297));
  assign _zz_4570 = ({9'd0,data_mid_1_53_imag} <<< 9);
  assign _zz_4571 = {{9{_zz_4570[26]}}, _zz_4570};
  assign _zz_4572 = fixTo_359_dout;
  assign _zz_4573 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_4574 = ($signed(_zz_303) - $signed(_zz_4575));
  assign _zz_4575 = ($signed(_zz_4576) * $signed(twiddle_factor_table_1_imag));
  assign _zz_4576 = ($signed(data_mid_1_58_real) + $signed(data_mid_1_58_imag));
  assign _zz_4577 = fixTo_360_dout;
  assign _zz_4578 = ($signed(_zz_303) + $signed(_zz_4579));
  assign _zz_4579 = ($signed(_zz_4580) * $signed(twiddle_factor_table_1_real));
  assign _zz_4580 = ($signed(data_mid_1_58_imag) - $signed(data_mid_1_58_real));
  assign _zz_4581 = fixTo_361_dout;
  assign _zz_4582 = _zz_4583[35 : 0];
  assign _zz_4583 = _zz_4584;
  assign _zz_4584 = ($signed(_zz_4585) >>> _zz_304);
  assign _zz_4585 = _zz_4586;
  assign _zz_4586 = ($signed(_zz_4588) - $signed(_zz_301));
  assign _zz_4587 = ({9'd0,data_mid_1_56_real} <<< 9);
  assign _zz_4588 = {{9{_zz_4587[26]}}, _zz_4587};
  assign _zz_4589 = fixTo_362_dout;
  assign _zz_4590 = _zz_4591[35 : 0];
  assign _zz_4591 = _zz_4592;
  assign _zz_4592 = ($signed(_zz_4593) >>> _zz_304);
  assign _zz_4593 = _zz_4594;
  assign _zz_4594 = ($signed(_zz_4596) - $signed(_zz_302));
  assign _zz_4595 = ({9'd0,data_mid_1_56_imag} <<< 9);
  assign _zz_4596 = {{9{_zz_4595[26]}}, _zz_4595};
  assign _zz_4597 = fixTo_363_dout;
  assign _zz_4598 = _zz_4599[35 : 0];
  assign _zz_4599 = _zz_4600;
  assign _zz_4600 = ($signed(_zz_4601) >>> _zz_305);
  assign _zz_4601 = _zz_4602;
  assign _zz_4602 = ($signed(_zz_4604) + $signed(_zz_301));
  assign _zz_4603 = ({9'd0,data_mid_1_56_real} <<< 9);
  assign _zz_4604 = {{9{_zz_4603[26]}}, _zz_4603};
  assign _zz_4605 = fixTo_364_dout;
  assign _zz_4606 = _zz_4607[35 : 0];
  assign _zz_4607 = _zz_4608;
  assign _zz_4608 = ($signed(_zz_4609) >>> _zz_305);
  assign _zz_4609 = _zz_4610;
  assign _zz_4610 = ($signed(_zz_4612) + $signed(_zz_302));
  assign _zz_4611 = ({9'd0,data_mid_1_56_imag} <<< 9);
  assign _zz_4612 = {{9{_zz_4611[26]}}, _zz_4611};
  assign _zz_4613 = fixTo_365_dout;
  assign _zz_4614 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_4615 = ($signed(_zz_308) - $signed(_zz_4616));
  assign _zz_4616 = ($signed(_zz_4617) * $signed(twiddle_factor_table_2_imag));
  assign _zz_4617 = ($signed(data_mid_1_59_real) + $signed(data_mid_1_59_imag));
  assign _zz_4618 = fixTo_366_dout;
  assign _zz_4619 = ($signed(_zz_308) + $signed(_zz_4620));
  assign _zz_4620 = ($signed(_zz_4621) * $signed(twiddle_factor_table_2_real));
  assign _zz_4621 = ($signed(data_mid_1_59_imag) - $signed(data_mid_1_59_real));
  assign _zz_4622 = fixTo_367_dout;
  assign _zz_4623 = _zz_4624[35 : 0];
  assign _zz_4624 = _zz_4625;
  assign _zz_4625 = ($signed(_zz_4626) >>> _zz_309);
  assign _zz_4626 = _zz_4627;
  assign _zz_4627 = ($signed(_zz_4629) - $signed(_zz_306));
  assign _zz_4628 = ({9'd0,data_mid_1_57_real} <<< 9);
  assign _zz_4629 = {{9{_zz_4628[26]}}, _zz_4628};
  assign _zz_4630 = fixTo_368_dout;
  assign _zz_4631 = _zz_4632[35 : 0];
  assign _zz_4632 = _zz_4633;
  assign _zz_4633 = ($signed(_zz_4634) >>> _zz_309);
  assign _zz_4634 = _zz_4635;
  assign _zz_4635 = ($signed(_zz_4637) - $signed(_zz_307));
  assign _zz_4636 = ({9'd0,data_mid_1_57_imag} <<< 9);
  assign _zz_4637 = {{9{_zz_4636[26]}}, _zz_4636};
  assign _zz_4638 = fixTo_369_dout;
  assign _zz_4639 = _zz_4640[35 : 0];
  assign _zz_4640 = _zz_4641;
  assign _zz_4641 = ($signed(_zz_4642) >>> _zz_310);
  assign _zz_4642 = _zz_4643;
  assign _zz_4643 = ($signed(_zz_4645) + $signed(_zz_306));
  assign _zz_4644 = ({9'd0,data_mid_1_57_real} <<< 9);
  assign _zz_4645 = {{9{_zz_4644[26]}}, _zz_4644};
  assign _zz_4646 = fixTo_370_dout;
  assign _zz_4647 = _zz_4648[35 : 0];
  assign _zz_4648 = _zz_4649;
  assign _zz_4649 = ($signed(_zz_4650) >>> _zz_310);
  assign _zz_4650 = _zz_4651;
  assign _zz_4651 = ($signed(_zz_4653) + $signed(_zz_307));
  assign _zz_4652 = ({9'd0,data_mid_1_57_imag} <<< 9);
  assign _zz_4653 = {{9{_zz_4652[26]}}, _zz_4652};
  assign _zz_4654 = fixTo_371_dout;
  assign _zz_4655 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_4656 = ($signed(_zz_313) - $signed(_zz_4657));
  assign _zz_4657 = ($signed(_zz_4658) * $signed(twiddle_factor_table_1_imag));
  assign _zz_4658 = ($signed(data_mid_1_62_real) + $signed(data_mid_1_62_imag));
  assign _zz_4659 = fixTo_372_dout;
  assign _zz_4660 = ($signed(_zz_313) + $signed(_zz_4661));
  assign _zz_4661 = ($signed(_zz_4662) * $signed(twiddle_factor_table_1_real));
  assign _zz_4662 = ($signed(data_mid_1_62_imag) - $signed(data_mid_1_62_real));
  assign _zz_4663 = fixTo_373_dout;
  assign _zz_4664 = _zz_4665[35 : 0];
  assign _zz_4665 = _zz_4666;
  assign _zz_4666 = ($signed(_zz_4667) >>> _zz_314);
  assign _zz_4667 = _zz_4668;
  assign _zz_4668 = ($signed(_zz_4670) - $signed(_zz_311));
  assign _zz_4669 = ({9'd0,data_mid_1_60_real} <<< 9);
  assign _zz_4670 = {{9{_zz_4669[26]}}, _zz_4669};
  assign _zz_4671 = fixTo_374_dout;
  assign _zz_4672 = _zz_4673[35 : 0];
  assign _zz_4673 = _zz_4674;
  assign _zz_4674 = ($signed(_zz_4675) >>> _zz_314);
  assign _zz_4675 = _zz_4676;
  assign _zz_4676 = ($signed(_zz_4678) - $signed(_zz_312));
  assign _zz_4677 = ({9'd0,data_mid_1_60_imag} <<< 9);
  assign _zz_4678 = {{9{_zz_4677[26]}}, _zz_4677};
  assign _zz_4679 = fixTo_375_dout;
  assign _zz_4680 = _zz_4681[35 : 0];
  assign _zz_4681 = _zz_4682;
  assign _zz_4682 = ($signed(_zz_4683) >>> _zz_315);
  assign _zz_4683 = _zz_4684;
  assign _zz_4684 = ($signed(_zz_4686) + $signed(_zz_311));
  assign _zz_4685 = ({9'd0,data_mid_1_60_real} <<< 9);
  assign _zz_4686 = {{9{_zz_4685[26]}}, _zz_4685};
  assign _zz_4687 = fixTo_376_dout;
  assign _zz_4688 = _zz_4689[35 : 0];
  assign _zz_4689 = _zz_4690;
  assign _zz_4690 = ($signed(_zz_4691) >>> _zz_315);
  assign _zz_4691 = _zz_4692;
  assign _zz_4692 = ($signed(_zz_4694) + $signed(_zz_312));
  assign _zz_4693 = ({9'd0,data_mid_1_60_imag} <<< 9);
  assign _zz_4694 = {{9{_zz_4693[26]}}, _zz_4693};
  assign _zz_4695 = fixTo_377_dout;
  assign _zz_4696 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_4697 = ($signed(_zz_318) - $signed(_zz_4698));
  assign _zz_4698 = ($signed(_zz_4699) * $signed(twiddle_factor_table_2_imag));
  assign _zz_4699 = ($signed(data_mid_1_63_real) + $signed(data_mid_1_63_imag));
  assign _zz_4700 = fixTo_378_dout;
  assign _zz_4701 = ($signed(_zz_318) + $signed(_zz_4702));
  assign _zz_4702 = ($signed(_zz_4703) * $signed(twiddle_factor_table_2_real));
  assign _zz_4703 = ($signed(data_mid_1_63_imag) - $signed(data_mid_1_63_real));
  assign _zz_4704 = fixTo_379_dout;
  assign _zz_4705 = _zz_4706[35 : 0];
  assign _zz_4706 = _zz_4707;
  assign _zz_4707 = ($signed(_zz_4708) >>> _zz_319);
  assign _zz_4708 = _zz_4709;
  assign _zz_4709 = ($signed(_zz_4711) - $signed(_zz_316));
  assign _zz_4710 = ({9'd0,data_mid_1_61_real} <<< 9);
  assign _zz_4711 = {{9{_zz_4710[26]}}, _zz_4710};
  assign _zz_4712 = fixTo_380_dout;
  assign _zz_4713 = _zz_4714[35 : 0];
  assign _zz_4714 = _zz_4715;
  assign _zz_4715 = ($signed(_zz_4716) >>> _zz_319);
  assign _zz_4716 = _zz_4717;
  assign _zz_4717 = ($signed(_zz_4719) - $signed(_zz_317));
  assign _zz_4718 = ({9'd0,data_mid_1_61_imag} <<< 9);
  assign _zz_4719 = {{9{_zz_4718[26]}}, _zz_4718};
  assign _zz_4720 = fixTo_381_dout;
  assign _zz_4721 = _zz_4722[35 : 0];
  assign _zz_4722 = _zz_4723;
  assign _zz_4723 = ($signed(_zz_4724) >>> _zz_320);
  assign _zz_4724 = _zz_4725;
  assign _zz_4725 = ($signed(_zz_4727) + $signed(_zz_316));
  assign _zz_4726 = ({9'd0,data_mid_1_61_real} <<< 9);
  assign _zz_4727 = {{9{_zz_4726[26]}}, _zz_4726};
  assign _zz_4728 = fixTo_382_dout;
  assign _zz_4729 = _zz_4730[35 : 0];
  assign _zz_4730 = _zz_4731;
  assign _zz_4731 = ($signed(_zz_4732) >>> _zz_320);
  assign _zz_4732 = _zz_4733;
  assign _zz_4733 = ($signed(_zz_4735) + $signed(_zz_317));
  assign _zz_4734 = ({9'd0,data_mid_1_61_imag} <<< 9);
  assign _zz_4735 = {{9{_zz_4734[26]}}, _zz_4734};
  assign _zz_4736 = fixTo_383_dout;
  assign _zz_4737 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_4738 = ($signed(_zz_323) - $signed(_zz_4739));
  assign _zz_4739 = ($signed(_zz_4740) * $signed(twiddle_factor_table_3_imag));
  assign _zz_4740 = ($signed(data_mid_2_4_real) + $signed(data_mid_2_4_imag));
  assign _zz_4741 = fixTo_384_dout;
  assign _zz_4742 = ($signed(_zz_323) + $signed(_zz_4743));
  assign _zz_4743 = ($signed(_zz_4744) * $signed(twiddle_factor_table_3_real));
  assign _zz_4744 = ($signed(data_mid_2_4_imag) - $signed(data_mid_2_4_real));
  assign _zz_4745 = fixTo_385_dout;
  assign _zz_4746 = _zz_4747[35 : 0];
  assign _zz_4747 = _zz_4748;
  assign _zz_4748 = ($signed(_zz_4749) >>> _zz_324);
  assign _zz_4749 = _zz_4750;
  assign _zz_4750 = ($signed(_zz_4752) - $signed(_zz_321));
  assign _zz_4751 = ({9'd0,data_mid_2_0_real} <<< 9);
  assign _zz_4752 = {{9{_zz_4751[26]}}, _zz_4751};
  assign _zz_4753 = fixTo_386_dout;
  assign _zz_4754 = _zz_4755[35 : 0];
  assign _zz_4755 = _zz_4756;
  assign _zz_4756 = ($signed(_zz_4757) >>> _zz_324);
  assign _zz_4757 = _zz_4758;
  assign _zz_4758 = ($signed(_zz_4760) - $signed(_zz_322));
  assign _zz_4759 = ({9'd0,data_mid_2_0_imag} <<< 9);
  assign _zz_4760 = {{9{_zz_4759[26]}}, _zz_4759};
  assign _zz_4761 = fixTo_387_dout;
  assign _zz_4762 = _zz_4763[35 : 0];
  assign _zz_4763 = _zz_4764;
  assign _zz_4764 = ($signed(_zz_4765) >>> _zz_325);
  assign _zz_4765 = _zz_4766;
  assign _zz_4766 = ($signed(_zz_4768) + $signed(_zz_321));
  assign _zz_4767 = ({9'd0,data_mid_2_0_real} <<< 9);
  assign _zz_4768 = {{9{_zz_4767[26]}}, _zz_4767};
  assign _zz_4769 = fixTo_388_dout;
  assign _zz_4770 = _zz_4771[35 : 0];
  assign _zz_4771 = _zz_4772;
  assign _zz_4772 = ($signed(_zz_4773) >>> _zz_325);
  assign _zz_4773 = _zz_4774;
  assign _zz_4774 = ($signed(_zz_4776) + $signed(_zz_322));
  assign _zz_4775 = ({9'd0,data_mid_2_0_imag} <<< 9);
  assign _zz_4776 = {{9{_zz_4775[26]}}, _zz_4775};
  assign _zz_4777 = fixTo_389_dout;
  assign _zz_4778 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_4779 = ($signed(_zz_328) - $signed(_zz_4780));
  assign _zz_4780 = ($signed(_zz_4781) * $signed(twiddle_factor_table_4_imag));
  assign _zz_4781 = ($signed(data_mid_2_5_real) + $signed(data_mid_2_5_imag));
  assign _zz_4782 = fixTo_390_dout;
  assign _zz_4783 = ($signed(_zz_328) + $signed(_zz_4784));
  assign _zz_4784 = ($signed(_zz_4785) * $signed(twiddle_factor_table_4_real));
  assign _zz_4785 = ($signed(data_mid_2_5_imag) - $signed(data_mid_2_5_real));
  assign _zz_4786 = fixTo_391_dout;
  assign _zz_4787 = _zz_4788[35 : 0];
  assign _zz_4788 = _zz_4789;
  assign _zz_4789 = ($signed(_zz_4790) >>> _zz_329);
  assign _zz_4790 = _zz_4791;
  assign _zz_4791 = ($signed(_zz_4793) - $signed(_zz_326));
  assign _zz_4792 = ({9'd0,data_mid_2_1_real} <<< 9);
  assign _zz_4793 = {{9{_zz_4792[26]}}, _zz_4792};
  assign _zz_4794 = fixTo_392_dout;
  assign _zz_4795 = _zz_4796[35 : 0];
  assign _zz_4796 = _zz_4797;
  assign _zz_4797 = ($signed(_zz_4798) >>> _zz_329);
  assign _zz_4798 = _zz_4799;
  assign _zz_4799 = ($signed(_zz_4801) - $signed(_zz_327));
  assign _zz_4800 = ({9'd0,data_mid_2_1_imag} <<< 9);
  assign _zz_4801 = {{9{_zz_4800[26]}}, _zz_4800};
  assign _zz_4802 = fixTo_393_dout;
  assign _zz_4803 = _zz_4804[35 : 0];
  assign _zz_4804 = _zz_4805;
  assign _zz_4805 = ($signed(_zz_4806) >>> _zz_330);
  assign _zz_4806 = _zz_4807;
  assign _zz_4807 = ($signed(_zz_4809) + $signed(_zz_326));
  assign _zz_4808 = ({9'd0,data_mid_2_1_real} <<< 9);
  assign _zz_4809 = {{9{_zz_4808[26]}}, _zz_4808};
  assign _zz_4810 = fixTo_394_dout;
  assign _zz_4811 = _zz_4812[35 : 0];
  assign _zz_4812 = _zz_4813;
  assign _zz_4813 = ($signed(_zz_4814) >>> _zz_330);
  assign _zz_4814 = _zz_4815;
  assign _zz_4815 = ($signed(_zz_4817) + $signed(_zz_327));
  assign _zz_4816 = ({9'd0,data_mid_2_1_imag} <<< 9);
  assign _zz_4817 = {{9{_zz_4816[26]}}, _zz_4816};
  assign _zz_4818 = fixTo_395_dout;
  assign _zz_4819 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_4820 = ($signed(_zz_333) - $signed(_zz_4821));
  assign _zz_4821 = ($signed(_zz_4822) * $signed(twiddle_factor_table_5_imag));
  assign _zz_4822 = ($signed(data_mid_2_6_real) + $signed(data_mid_2_6_imag));
  assign _zz_4823 = fixTo_396_dout;
  assign _zz_4824 = ($signed(_zz_333) + $signed(_zz_4825));
  assign _zz_4825 = ($signed(_zz_4826) * $signed(twiddle_factor_table_5_real));
  assign _zz_4826 = ($signed(data_mid_2_6_imag) - $signed(data_mid_2_6_real));
  assign _zz_4827 = fixTo_397_dout;
  assign _zz_4828 = _zz_4829[35 : 0];
  assign _zz_4829 = _zz_4830;
  assign _zz_4830 = ($signed(_zz_4831) >>> _zz_334);
  assign _zz_4831 = _zz_4832;
  assign _zz_4832 = ($signed(_zz_4834) - $signed(_zz_331));
  assign _zz_4833 = ({9'd0,data_mid_2_2_real} <<< 9);
  assign _zz_4834 = {{9{_zz_4833[26]}}, _zz_4833};
  assign _zz_4835 = fixTo_398_dout;
  assign _zz_4836 = _zz_4837[35 : 0];
  assign _zz_4837 = _zz_4838;
  assign _zz_4838 = ($signed(_zz_4839) >>> _zz_334);
  assign _zz_4839 = _zz_4840;
  assign _zz_4840 = ($signed(_zz_4842) - $signed(_zz_332));
  assign _zz_4841 = ({9'd0,data_mid_2_2_imag} <<< 9);
  assign _zz_4842 = {{9{_zz_4841[26]}}, _zz_4841};
  assign _zz_4843 = fixTo_399_dout;
  assign _zz_4844 = _zz_4845[35 : 0];
  assign _zz_4845 = _zz_4846;
  assign _zz_4846 = ($signed(_zz_4847) >>> _zz_335);
  assign _zz_4847 = _zz_4848;
  assign _zz_4848 = ($signed(_zz_4850) + $signed(_zz_331));
  assign _zz_4849 = ({9'd0,data_mid_2_2_real} <<< 9);
  assign _zz_4850 = {{9{_zz_4849[26]}}, _zz_4849};
  assign _zz_4851 = fixTo_400_dout;
  assign _zz_4852 = _zz_4853[35 : 0];
  assign _zz_4853 = _zz_4854;
  assign _zz_4854 = ($signed(_zz_4855) >>> _zz_335);
  assign _zz_4855 = _zz_4856;
  assign _zz_4856 = ($signed(_zz_4858) + $signed(_zz_332));
  assign _zz_4857 = ({9'd0,data_mid_2_2_imag} <<< 9);
  assign _zz_4858 = {{9{_zz_4857[26]}}, _zz_4857};
  assign _zz_4859 = fixTo_401_dout;
  assign _zz_4860 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_4861 = ($signed(_zz_338) - $signed(_zz_4862));
  assign _zz_4862 = ($signed(_zz_4863) * $signed(twiddle_factor_table_6_imag));
  assign _zz_4863 = ($signed(data_mid_2_7_real) + $signed(data_mid_2_7_imag));
  assign _zz_4864 = fixTo_402_dout;
  assign _zz_4865 = ($signed(_zz_338) + $signed(_zz_4866));
  assign _zz_4866 = ($signed(_zz_4867) * $signed(twiddle_factor_table_6_real));
  assign _zz_4867 = ($signed(data_mid_2_7_imag) - $signed(data_mid_2_7_real));
  assign _zz_4868 = fixTo_403_dout;
  assign _zz_4869 = _zz_4870[35 : 0];
  assign _zz_4870 = _zz_4871;
  assign _zz_4871 = ($signed(_zz_4872) >>> _zz_339);
  assign _zz_4872 = _zz_4873;
  assign _zz_4873 = ($signed(_zz_4875) - $signed(_zz_336));
  assign _zz_4874 = ({9'd0,data_mid_2_3_real} <<< 9);
  assign _zz_4875 = {{9{_zz_4874[26]}}, _zz_4874};
  assign _zz_4876 = fixTo_404_dout;
  assign _zz_4877 = _zz_4878[35 : 0];
  assign _zz_4878 = _zz_4879;
  assign _zz_4879 = ($signed(_zz_4880) >>> _zz_339);
  assign _zz_4880 = _zz_4881;
  assign _zz_4881 = ($signed(_zz_4883) - $signed(_zz_337));
  assign _zz_4882 = ({9'd0,data_mid_2_3_imag} <<< 9);
  assign _zz_4883 = {{9{_zz_4882[26]}}, _zz_4882};
  assign _zz_4884 = fixTo_405_dout;
  assign _zz_4885 = _zz_4886[35 : 0];
  assign _zz_4886 = _zz_4887;
  assign _zz_4887 = ($signed(_zz_4888) >>> _zz_340);
  assign _zz_4888 = _zz_4889;
  assign _zz_4889 = ($signed(_zz_4891) + $signed(_zz_336));
  assign _zz_4890 = ({9'd0,data_mid_2_3_real} <<< 9);
  assign _zz_4891 = {{9{_zz_4890[26]}}, _zz_4890};
  assign _zz_4892 = fixTo_406_dout;
  assign _zz_4893 = _zz_4894[35 : 0];
  assign _zz_4894 = _zz_4895;
  assign _zz_4895 = ($signed(_zz_4896) >>> _zz_340);
  assign _zz_4896 = _zz_4897;
  assign _zz_4897 = ($signed(_zz_4899) + $signed(_zz_337));
  assign _zz_4898 = ({9'd0,data_mid_2_3_imag} <<< 9);
  assign _zz_4899 = {{9{_zz_4898[26]}}, _zz_4898};
  assign _zz_4900 = fixTo_407_dout;
  assign _zz_4901 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_4902 = ($signed(_zz_343) - $signed(_zz_4903));
  assign _zz_4903 = ($signed(_zz_4904) * $signed(twiddle_factor_table_3_imag));
  assign _zz_4904 = ($signed(data_mid_2_12_real) + $signed(data_mid_2_12_imag));
  assign _zz_4905 = fixTo_408_dout;
  assign _zz_4906 = ($signed(_zz_343) + $signed(_zz_4907));
  assign _zz_4907 = ($signed(_zz_4908) * $signed(twiddle_factor_table_3_real));
  assign _zz_4908 = ($signed(data_mid_2_12_imag) - $signed(data_mid_2_12_real));
  assign _zz_4909 = fixTo_409_dout;
  assign _zz_4910 = _zz_4911[35 : 0];
  assign _zz_4911 = _zz_4912;
  assign _zz_4912 = ($signed(_zz_4913) >>> _zz_344);
  assign _zz_4913 = _zz_4914;
  assign _zz_4914 = ($signed(_zz_4916) - $signed(_zz_341));
  assign _zz_4915 = ({9'd0,data_mid_2_8_real} <<< 9);
  assign _zz_4916 = {{9{_zz_4915[26]}}, _zz_4915};
  assign _zz_4917 = fixTo_410_dout;
  assign _zz_4918 = _zz_4919[35 : 0];
  assign _zz_4919 = _zz_4920;
  assign _zz_4920 = ($signed(_zz_4921) >>> _zz_344);
  assign _zz_4921 = _zz_4922;
  assign _zz_4922 = ($signed(_zz_4924) - $signed(_zz_342));
  assign _zz_4923 = ({9'd0,data_mid_2_8_imag} <<< 9);
  assign _zz_4924 = {{9{_zz_4923[26]}}, _zz_4923};
  assign _zz_4925 = fixTo_411_dout;
  assign _zz_4926 = _zz_4927[35 : 0];
  assign _zz_4927 = _zz_4928;
  assign _zz_4928 = ($signed(_zz_4929) >>> _zz_345);
  assign _zz_4929 = _zz_4930;
  assign _zz_4930 = ($signed(_zz_4932) + $signed(_zz_341));
  assign _zz_4931 = ({9'd0,data_mid_2_8_real} <<< 9);
  assign _zz_4932 = {{9{_zz_4931[26]}}, _zz_4931};
  assign _zz_4933 = fixTo_412_dout;
  assign _zz_4934 = _zz_4935[35 : 0];
  assign _zz_4935 = _zz_4936;
  assign _zz_4936 = ($signed(_zz_4937) >>> _zz_345);
  assign _zz_4937 = _zz_4938;
  assign _zz_4938 = ($signed(_zz_4940) + $signed(_zz_342));
  assign _zz_4939 = ({9'd0,data_mid_2_8_imag} <<< 9);
  assign _zz_4940 = {{9{_zz_4939[26]}}, _zz_4939};
  assign _zz_4941 = fixTo_413_dout;
  assign _zz_4942 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_4943 = ($signed(_zz_348) - $signed(_zz_4944));
  assign _zz_4944 = ($signed(_zz_4945) * $signed(twiddle_factor_table_4_imag));
  assign _zz_4945 = ($signed(data_mid_2_13_real) + $signed(data_mid_2_13_imag));
  assign _zz_4946 = fixTo_414_dout;
  assign _zz_4947 = ($signed(_zz_348) + $signed(_zz_4948));
  assign _zz_4948 = ($signed(_zz_4949) * $signed(twiddle_factor_table_4_real));
  assign _zz_4949 = ($signed(data_mid_2_13_imag) - $signed(data_mid_2_13_real));
  assign _zz_4950 = fixTo_415_dout;
  assign _zz_4951 = _zz_4952[35 : 0];
  assign _zz_4952 = _zz_4953;
  assign _zz_4953 = ($signed(_zz_4954) >>> _zz_349);
  assign _zz_4954 = _zz_4955;
  assign _zz_4955 = ($signed(_zz_4957) - $signed(_zz_346));
  assign _zz_4956 = ({9'd0,data_mid_2_9_real} <<< 9);
  assign _zz_4957 = {{9{_zz_4956[26]}}, _zz_4956};
  assign _zz_4958 = fixTo_416_dout;
  assign _zz_4959 = _zz_4960[35 : 0];
  assign _zz_4960 = _zz_4961;
  assign _zz_4961 = ($signed(_zz_4962) >>> _zz_349);
  assign _zz_4962 = _zz_4963;
  assign _zz_4963 = ($signed(_zz_4965) - $signed(_zz_347));
  assign _zz_4964 = ({9'd0,data_mid_2_9_imag} <<< 9);
  assign _zz_4965 = {{9{_zz_4964[26]}}, _zz_4964};
  assign _zz_4966 = fixTo_417_dout;
  assign _zz_4967 = _zz_4968[35 : 0];
  assign _zz_4968 = _zz_4969;
  assign _zz_4969 = ($signed(_zz_4970) >>> _zz_350);
  assign _zz_4970 = _zz_4971;
  assign _zz_4971 = ($signed(_zz_4973) + $signed(_zz_346));
  assign _zz_4972 = ({9'd0,data_mid_2_9_real} <<< 9);
  assign _zz_4973 = {{9{_zz_4972[26]}}, _zz_4972};
  assign _zz_4974 = fixTo_418_dout;
  assign _zz_4975 = _zz_4976[35 : 0];
  assign _zz_4976 = _zz_4977;
  assign _zz_4977 = ($signed(_zz_4978) >>> _zz_350);
  assign _zz_4978 = _zz_4979;
  assign _zz_4979 = ($signed(_zz_4981) + $signed(_zz_347));
  assign _zz_4980 = ({9'd0,data_mid_2_9_imag} <<< 9);
  assign _zz_4981 = {{9{_zz_4980[26]}}, _zz_4980};
  assign _zz_4982 = fixTo_419_dout;
  assign _zz_4983 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_4984 = ($signed(_zz_353) - $signed(_zz_4985));
  assign _zz_4985 = ($signed(_zz_4986) * $signed(twiddle_factor_table_5_imag));
  assign _zz_4986 = ($signed(data_mid_2_14_real) + $signed(data_mid_2_14_imag));
  assign _zz_4987 = fixTo_420_dout;
  assign _zz_4988 = ($signed(_zz_353) + $signed(_zz_4989));
  assign _zz_4989 = ($signed(_zz_4990) * $signed(twiddle_factor_table_5_real));
  assign _zz_4990 = ($signed(data_mid_2_14_imag) - $signed(data_mid_2_14_real));
  assign _zz_4991 = fixTo_421_dout;
  assign _zz_4992 = _zz_4993[35 : 0];
  assign _zz_4993 = _zz_4994;
  assign _zz_4994 = ($signed(_zz_4995) >>> _zz_354);
  assign _zz_4995 = _zz_4996;
  assign _zz_4996 = ($signed(_zz_4998) - $signed(_zz_351));
  assign _zz_4997 = ({9'd0,data_mid_2_10_real} <<< 9);
  assign _zz_4998 = {{9{_zz_4997[26]}}, _zz_4997};
  assign _zz_4999 = fixTo_422_dout;
  assign _zz_5000 = _zz_5001[35 : 0];
  assign _zz_5001 = _zz_5002;
  assign _zz_5002 = ($signed(_zz_5003) >>> _zz_354);
  assign _zz_5003 = _zz_5004;
  assign _zz_5004 = ($signed(_zz_5006) - $signed(_zz_352));
  assign _zz_5005 = ({9'd0,data_mid_2_10_imag} <<< 9);
  assign _zz_5006 = {{9{_zz_5005[26]}}, _zz_5005};
  assign _zz_5007 = fixTo_423_dout;
  assign _zz_5008 = _zz_5009[35 : 0];
  assign _zz_5009 = _zz_5010;
  assign _zz_5010 = ($signed(_zz_5011) >>> _zz_355);
  assign _zz_5011 = _zz_5012;
  assign _zz_5012 = ($signed(_zz_5014) + $signed(_zz_351));
  assign _zz_5013 = ({9'd0,data_mid_2_10_real} <<< 9);
  assign _zz_5014 = {{9{_zz_5013[26]}}, _zz_5013};
  assign _zz_5015 = fixTo_424_dout;
  assign _zz_5016 = _zz_5017[35 : 0];
  assign _zz_5017 = _zz_5018;
  assign _zz_5018 = ($signed(_zz_5019) >>> _zz_355);
  assign _zz_5019 = _zz_5020;
  assign _zz_5020 = ($signed(_zz_5022) + $signed(_zz_352));
  assign _zz_5021 = ({9'd0,data_mid_2_10_imag} <<< 9);
  assign _zz_5022 = {{9{_zz_5021[26]}}, _zz_5021};
  assign _zz_5023 = fixTo_425_dout;
  assign _zz_5024 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_5025 = ($signed(_zz_358) - $signed(_zz_5026));
  assign _zz_5026 = ($signed(_zz_5027) * $signed(twiddle_factor_table_6_imag));
  assign _zz_5027 = ($signed(data_mid_2_15_real) + $signed(data_mid_2_15_imag));
  assign _zz_5028 = fixTo_426_dout;
  assign _zz_5029 = ($signed(_zz_358) + $signed(_zz_5030));
  assign _zz_5030 = ($signed(_zz_5031) * $signed(twiddle_factor_table_6_real));
  assign _zz_5031 = ($signed(data_mid_2_15_imag) - $signed(data_mid_2_15_real));
  assign _zz_5032 = fixTo_427_dout;
  assign _zz_5033 = _zz_5034[35 : 0];
  assign _zz_5034 = _zz_5035;
  assign _zz_5035 = ($signed(_zz_5036) >>> _zz_359);
  assign _zz_5036 = _zz_5037;
  assign _zz_5037 = ($signed(_zz_5039) - $signed(_zz_356));
  assign _zz_5038 = ({9'd0,data_mid_2_11_real} <<< 9);
  assign _zz_5039 = {{9{_zz_5038[26]}}, _zz_5038};
  assign _zz_5040 = fixTo_428_dout;
  assign _zz_5041 = _zz_5042[35 : 0];
  assign _zz_5042 = _zz_5043;
  assign _zz_5043 = ($signed(_zz_5044) >>> _zz_359);
  assign _zz_5044 = _zz_5045;
  assign _zz_5045 = ($signed(_zz_5047) - $signed(_zz_357));
  assign _zz_5046 = ({9'd0,data_mid_2_11_imag} <<< 9);
  assign _zz_5047 = {{9{_zz_5046[26]}}, _zz_5046};
  assign _zz_5048 = fixTo_429_dout;
  assign _zz_5049 = _zz_5050[35 : 0];
  assign _zz_5050 = _zz_5051;
  assign _zz_5051 = ($signed(_zz_5052) >>> _zz_360);
  assign _zz_5052 = _zz_5053;
  assign _zz_5053 = ($signed(_zz_5055) + $signed(_zz_356));
  assign _zz_5054 = ({9'd0,data_mid_2_11_real} <<< 9);
  assign _zz_5055 = {{9{_zz_5054[26]}}, _zz_5054};
  assign _zz_5056 = fixTo_430_dout;
  assign _zz_5057 = _zz_5058[35 : 0];
  assign _zz_5058 = _zz_5059;
  assign _zz_5059 = ($signed(_zz_5060) >>> _zz_360);
  assign _zz_5060 = _zz_5061;
  assign _zz_5061 = ($signed(_zz_5063) + $signed(_zz_357));
  assign _zz_5062 = ({9'd0,data_mid_2_11_imag} <<< 9);
  assign _zz_5063 = {{9{_zz_5062[26]}}, _zz_5062};
  assign _zz_5064 = fixTo_431_dout;
  assign _zz_5065 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_5066 = ($signed(_zz_363) - $signed(_zz_5067));
  assign _zz_5067 = ($signed(_zz_5068) * $signed(twiddle_factor_table_3_imag));
  assign _zz_5068 = ($signed(data_mid_2_20_real) + $signed(data_mid_2_20_imag));
  assign _zz_5069 = fixTo_432_dout;
  assign _zz_5070 = ($signed(_zz_363) + $signed(_zz_5071));
  assign _zz_5071 = ($signed(_zz_5072) * $signed(twiddle_factor_table_3_real));
  assign _zz_5072 = ($signed(data_mid_2_20_imag) - $signed(data_mid_2_20_real));
  assign _zz_5073 = fixTo_433_dout;
  assign _zz_5074 = _zz_5075[35 : 0];
  assign _zz_5075 = _zz_5076;
  assign _zz_5076 = ($signed(_zz_5077) >>> _zz_364);
  assign _zz_5077 = _zz_5078;
  assign _zz_5078 = ($signed(_zz_5080) - $signed(_zz_361));
  assign _zz_5079 = ({9'd0,data_mid_2_16_real} <<< 9);
  assign _zz_5080 = {{9{_zz_5079[26]}}, _zz_5079};
  assign _zz_5081 = fixTo_434_dout;
  assign _zz_5082 = _zz_5083[35 : 0];
  assign _zz_5083 = _zz_5084;
  assign _zz_5084 = ($signed(_zz_5085) >>> _zz_364);
  assign _zz_5085 = _zz_5086;
  assign _zz_5086 = ($signed(_zz_5088) - $signed(_zz_362));
  assign _zz_5087 = ({9'd0,data_mid_2_16_imag} <<< 9);
  assign _zz_5088 = {{9{_zz_5087[26]}}, _zz_5087};
  assign _zz_5089 = fixTo_435_dout;
  assign _zz_5090 = _zz_5091[35 : 0];
  assign _zz_5091 = _zz_5092;
  assign _zz_5092 = ($signed(_zz_5093) >>> _zz_365);
  assign _zz_5093 = _zz_5094;
  assign _zz_5094 = ($signed(_zz_5096) + $signed(_zz_361));
  assign _zz_5095 = ({9'd0,data_mid_2_16_real} <<< 9);
  assign _zz_5096 = {{9{_zz_5095[26]}}, _zz_5095};
  assign _zz_5097 = fixTo_436_dout;
  assign _zz_5098 = _zz_5099[35 : 0];
  assign _zz_5099 = _zz_5100;
  assign _zz_5100 = ($signed(_zz_5101) >>> _zz_365);
  assign _zz_5101 = _zz_5102;
  assign _zz_5102 = ($signed(_zz_5104) + $signed(_zz_362));
  assign _zz_5103 = ({9'd0,data_mid_2_16_imag} <<< 9);
  assign _zz_5104 = {{9{_zz_5103[26]}}, _zz_5103};
  assign _zz_5105 = fixTo_437_dout;
  assign _zz_5106 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_5107 = ($signed(_zz_368) - $signed(_zz_5108));
  assign _zz_5108 = ($signed(_zz_5109) * $signed(twiddle_factor_table_4_imag));
  assign _zz_5109 = ($signed(data_mid_2_21_real) + $signed(data_mid_2_21_imag));
  assign _zz_5110 = fixTo_438_dout;
  assign _zz_5111 = ($signed(_zz_368) + $signed(_zz_5112));
  assign _zz_5112 = ($signed(_zz_5113) * $signed(twiddle_factor_table_4_real));
  assign _zz_5113 = ($signed(data_mid_2_21_imag) - $signed(data_mid_2_21_real));
  assign _zz_5114 = fixTo_439_dout;
  assign _zz_5115 = _zz_5116[35 : 0];
  assign _zz_5116 = _zz_5117;
  assign _zz_5117 = ($signed(_zz_5118) >>> _zz_369);
  assign _zz_5118 = _zz_5119;
  assign _zz_5119 = ($signed(_zz_5121) - $signed(_zz_366));
  assign _zz_5120 = ({9'd0,data_mid_2_17_real} <<< 9);
  assign _zz_5121 = {{9{_zz_5120[26]}}, _zz_5120};
  assign _zz_5122 = fixTo_440_dout;
  assign _zz_5123 = _zz_5124[35 : 0];
  assign _zz_5124 = _zz_5125;
  assign _zz_5125 = ($signed(_zz_5126) >>> _zz_369);
  assign _zz_5126 = _zz_5127;
  assign _zz_5127 = ($signed(_zz_5129) - $signed(_zz_367));
  assign _zz_5128 = ({9'd0,data_mid_2_17_imag} <<< 9);
  assign _zz_5129 = {{9{_zz_5128[26]}}, _zz_5128};
  assign _zz_5130 = fixTo_441_dout;
  assign _zz_5131 = _zz_5132[35 : 0];
  assign _zz_5132 = _zz_5133;
  assign _zz_5133 = ($signed(_zz_5134) >>> _zz_370);
  assign _zz_5134 = _zz_5135;
  assign _zz_5135 = ($signed(_zz_5137) + $signed(_zz_366));
  assign _zz_5136 = ({9'd0,data_mid_2_17_real} <<< 9);
  assign _zz_5137 = {{9{_zz_5136[26]}}, _zz_5136};
  assign _zz_5138 = fixTo_442_dout;
  assign _zz_5139 = _zz_5140[35 : 0];
  assign _zz_5140 = _zz_5141;
  assign _zz_5141 = ($signed(_zz_5142) >>> _zz_370);
  assign _zz_5142 = _zz_5143;
  assign _zz_5143 = ($signed(_zz_5145) + $signed(_zz_367));
  assign _zz_5144 = ({9'd0,data_mid_2_17_imag} <<< 9);
  assign _zz_5145 = {{9{_zz_5144[26]}}, _zz_5144};
  assign _zz_5146 = fixTo_443_dout;
  assign _zz_5147 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_5148 = ($signed(_zz_373) - $signed(_zz_5149));
  assign _zz_5149 = ($signed(_zz_5150) * $signed(twiddle_factor_table_5_imag));
  assign _zz_5150 = ($signed(data_mid_2_22_real) + $signed(data_mid_2_22_imag));
  assign _zz_5151 = fixTo_444_dout;
  assign _zz_5152 = ($signed(_zz_373) + $signed(_zz_5153));
  assign _zz_5153 = ($signed(_zz_5154) * $signed(twiddle_factor_table_5_real));
  assign _zz_5154 = ($signed(data_mid_2_22_imag) - $signed(data_mid_2_22_real));
  assign _zz_5155 = fixTo_445_dout;
  assign _zz_5156 = _zz_5157[35 : 0];
  assign _zz_5157 = _zz_5158;
  assign _zz_5158 = ($signed(_zz_5159) >>> _zz_374);
  assign _zz_5159 = _zz_5160;
  assign _zz_5160 = ($signed(_zz_5162) - $signed(_zz_371));
  assign _zz_5161 = ({9'd0,data_mid_2_18_real} <<< 9);
  assign _zz_5162 = {{9{_zz_5161[26]}}, _zz_5161};
  assign _zz_5163 = fixTo_446_dout;
  assign _zz_5164 = _zz_5165[35 : 0];
  assign _zz_5165 = _zz_5166;
  assign _zz_5166 = ($signed(_zz_5167) >>> _zz_374);
  assign _zz_5167 = _zz_5168;
  assign _zz_5168 = ($signed(_zz_5170) - $signed(_zz_372));
  assign _zz_5169 = ({9'd0,data_mid_2_18_imag} <<< 9);
  assign _zz_5170 = {{9{_zz_5169[26]}}, _zz_5169};
  assign _zz_5171 = fixTo_447_dout;
  assign _zz_5172 = _zz_5173[35 : 0];
  assign _zz_5173 = _zz_5174;
  assign _zz_5174 = ($signed(_zz_5175) >>> _zz_375);
  assign _zz_5175 = _zz_5176;
  assign _zz_5176 = ($signed(_zz_5178) + $signed(_zz_371));
  assign _zz_5177 = ({9'd0,data_mid_2_18_real} <<< 9);
  assign _zz_5178 = {{9{_zz_5177[26]}}, _zz_5177};
  assign _zz_5179 = fixTo_448_dout;
  assign _zz_5180 = _zz_5181[35 : 0];
  assign _zz_5181 = _zz_5182;
  assign _zz_5182 = ($signed(_zz_5183) >>> _zz_375);
  assign _zz_5183 = _zz_5184;
  assign _zz_5184 = ($signed(_zz_5186) + $signed(_zz_372));
  assign _zz_5185 = ({9'd0,data_mid_2_18_imag} <<< 9);
  assign _zz_5186 = {{9{_zz_5185[26]}}, _zz_5185};
  assign _zz_5187 = fixTo_449_dout;
  assign _zz_5188 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_5189 = ($signed(_zz_378) - $signed(_zz_5190));
  assign _zz_5190 = ($signed(_zz_5191) * $signed(twiddle_factor_table_6_imag));
  assign _zz_5191 = ($signed(data_mid_2_23_real) + $signed(data_mid_2_23_imag));
  assign _zz_5192 = fixTo_450_dout;
  assign _zz_5193 = ($signed(_zz_378) + $signed(_zz_5194));
  assign _zz_5194 = ($signed(_zz_5195) * $signed(twiddle_factor_table_6_real));
  assign _zz_5195 = ($signed(data_mid_2_23_imag) - $signed(data_mid_2_23_real));
  assign _zz_5196 = fixTo_451_dout;
  assign _zz_5197 = _zz_5198[35 : 0];
  assign _zz_5198 = _zz_5199;
  assign _zz_5199 = ($signed(_zz_5200) >>> _zz_379);
  assign _zz_5200 = _zz_5201;
  assign _zz_5201 = ($signed(_zz_5203) - $signed(_zz_376));
  assign _zz_5202 = ({9'd0,data_mid_2_19_real} <<< 9);
  assign _zz_5203 = {{9{_zz_5202[26]}}, _zz_5202};
  assign _zz_5204 = fixTo_452_dout;
  assign _zz_5205 = _zz_5206[35 : 0];
  assign _zz_5206 = _zz_5207;
  assign _zz_5207 = ($signed(_zz_5208) >>> _zz_379);
  assign _zz_5208 = _zz_5209;
  assign _zz_5209 = ($signed(_zz_5211) - $signed(_zz_377));
  assign _zz_5210 = ({9'd0,data_mid_2_19_imag} <<< 9);
  assign _zz_5211 = {{9{_zz_5210[26]}}, _zz_5210};
  assign _zz_5212 = fixTo_453_dout;
  assign _zz_5213 = _zz_5214[35 : 0];
  assign _zz_5214 = _zz_5215;
  assign _zz_5215 = ($signed(_zz_5216) >>> _zz_380);
  assign _zz_5216 = _zz_5217;
  assign _zz_5217 = ($signed(_zz_5219) + $signed(_zz_376));
  assign _zz_5218 = ({9'd0,data_mid_2_19_real} <<< 9);
  assign _zz_5219 = {{9{_zz_5218[26]}}, _zz_5218};
  assign _zz_5220 = fixTo_454_dout;
  assign _zz_5221 = _zz_5222[35 : 0];
  assign _zz_5222 = _zz_5223;
  assign _zz_5223 = ($signed(_zz_5224) >>> _zz_380);
  assign _zz_5224 = _zz_5225;
  assign _zz_5225 = ($signed(_zz_5227) + $signed(_zz_377));
  assign _zz_5226 = ({9'd0,data_mid_2_19_imag} <<< 9);
  assign _zz_5227 = {{9{_zz_5226[26]}}, _zz_5226};
  assign _zz_5228 = fixTo_455_dout;
  assign _zz_5229 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_5230 = ($signed(_zz_383) - $signed(_zz_5231));
  assign _zz_5231 = ($signed(_zz_5232) * $signed(twiddle_factor_table_3_imag));
  assign _zz_5232 = ($signed(data_mid_2_28_real) + $signed(data_mid_2_28_imag));
  assign _zz_5233 = fixTo_456_dout;
  assign _zz_5234 = ($signed(_zz_383) + $signed(_zz_5235));
  assign _zz_5235 = ($signed(_zz_5236) * $signed(twiddle_factor_table_3_real));
  assign _zz_5236 = ($signed(data_mid_2_28_imag) - $signed(data_mid_2_28_real));
  assign _zz_5237 = fixTo_457_dout;
  assign _zz_5238 = _zz_5239[35 : 0];
  assign _zz_5239 = _zz_5240;
  assign _zz_5240 = ($signed(_zz_5241) >>> _zz_384);
  assign _zz_5241 = _zz_5242;
  assign _zz_5242 = ($signed(_zz_5244) - $signed(_zz_381));
  assign _zz_5243 = ({9'd0,data_mid_2_24_real} <<< 9);
  assign _zz_5244 = {{9{_zz_5243[26]}}, _zz_5243};
  assign _zz_5245 = fixTo_458_dout;
  assign _zz_5246 = _zz_5247[35 : 0];
  assign _zz_5247 = _zz_5248;
  assign _zz_5248 = ($signed(_zz_5249) >>> _zz_384);
  assign _zz_5249 = _zz_5250;
  assign _zz_5250 = ($signed(_zz_5252) - $signed(_zz_382));
  assign _zz_5251 = ({9'd0,data_mid_2_24_imag} <<< 9);
  assign _zz_5252 = {{9{_zz_5251[26]}}, _zz_5251};
  assign _zz_5253 = fixTo_459_dout;
  assign _zz_5254 = _zz_5255[35 : 0];
  assign _zz_5255 = _zz_5256;
  assign _zz_5256 = ($signed(_zz_5257) >>> _zz_385);
  assign _zz_5257 = _zz_5258;
  assign _zz_5258 = ($signed(_zz_5260) + $signed(_zz_381));
  assign _zz_5259 = ({9'd0,data_mid_2_24_real} <<< 9);
  assign _zz_5260 = {{9{_zz_5259[26]}}, _zz_5259};
  assign _zz_5261 = fixTo_460_dout;
  assign _zz_5262 = _zz_5263[35 : 0];
  assign _zz_5263 = _zz_5264;
  assign _zz_5264 = ($signed(_zz_5265) >>> _zz_385);
  assign _zz_5265 = _zz_5266;
  assign _zz_5266 = ($signed(_zz_5268) + $signed(_zz_382));
  assign _zz_5267 = ({9'd0,data_mid_2_24_imag} <<< 9);
  assign _zz_5268 = {{9{_zz_5267[26]}}, _zz_5267};
  assign _zz_5269 = fixTo_461_dout;
  assign _zz_5270 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_5271 = ($signed(_zz_388) - $signed(_zz_5272));
  assign _zz_5272 = ($signed(_zz_5273) * $signed(twiddle_factor_table_4_imag));
  assign _zz_5273 = ($signed(data_mid_2_29_real) + $signed(data_mid_2_29_imag));
  assign _zz_5274 = fixTo_462_dout;
  assign _zz_5275 = ($signed(_zz_388) + $signed(_zz_5276));
  assign _zz_5276 = ($signed(_zz_5277) * $signed(twiddle_factor_table_4_real));
  assign _zz_5277 = ($signed(data_mid_2_29_imag) - $signed(data_mid_2_29_real));
  assign _zz_5278 = fixTo_463_dout;
  assign _zz_5279 = _zz_5280[35 : 0];
  assign _zz_5280 = _zz_5281;
  assign _zz_5281 = ($signed(_zz_5282) >>> _zz_389);
  assign _zz_5282 = _zz_5283;
  assign _zz_5283 = ($signed(_zz_5285) - $signed(_zz_386));
  assign _zz_5284 = ({9'd0,data_mid_2_25_real} <<< 9);
  assign _zz_5285 = {{9{_zz_5284[26]}}, _zz_5284};
  assign _zz_5286 = fixTo_464_dout;
  assign _zz_5287 = _zz_5288[35 : 0];
  assign _zz_5288 = _zz_5289;
  assign _zz_5289 = ($signed(_zz_5290) >>> _zz_389);
  assign _zz_5290 = _zz_5291;
  assign _zz_5291 = ($signed(_zz_5293) - $signed(_zz_387));
  assign _zz_5292 = ({9'd0,data_mid_2_25_imag} <<< 9);
  assign _zz_5293 = {{9{_zz_5292[26]}}, _zz_5292};
  assign _zz_5294 = fixTo_465_dout;
  assign _zz_5295 = _zz_5296[35 : 0];
  assign _zz_5296 = _zz_5297;
  assign _zz_5297 = ($signed(_zz_5298) >>> _zz_390);
  assign _zz_5298 = _zz_5299;
  assign _zz_5299 = ($signed(_zz_5301) + $signed(_zz_386));
  assign _zz_5300 = ({9'd0,data_mid_2_25_real} <<< 9);
  assign _zz_5301 = {{9{_zz_5300[26]}}, _zz_5300};
  assign _zz_5302 = fixTo_466_dout;
  assign _zz_5303 = _zz_5304[35 : 0];
  assign _zz_5304 = _zz_5305;
  assign _zz_5305 = ($signed(_zz_5306) >>> _zz_390);
  assign _zz_5306 = _zz_5307;
  assign _zz_5307 = ($signed(_zz_5309) + $signed(_zz_387));
  assign _zz_5308 = ({9'd0,data_mid_2_25_imag} <<< 9);
  assign _zz_5309 = {{9{_zz_5308[26]}}, _zz_5308};
  assign _zz_5310 = fixTo_467_dout;
  assign _zz_5311 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_5312 = ($signed(_zz_393) - $signed(_zz_5313));
  assign _zz_5313 = ($signed(_zz_5314) * $signed(twiddle_factor_table_5_imag));
  assign _zz_5314 = ($signed(data_mid_2_30_real) + $signed(data_mid_2_30_imag));
  assign _zz_5315 = fixTo_468_dout;
  assign _zz_5316 = ($signed(_zz_393) + $signed(_zz_5317));
  assign _zz_5317 = ($signed(_zz_5318) * $signed(twiddle_factor_table_5_real));
  assign _zz_5318 = ($signed(data_mid_2_30_imag) - $signed(data_mid_2_30_real));
  assign _zz_5319 = fixTo_469_dout;
  assign _zz_5320 = _zz_5321[35 : 0];
  assign _zz_5321 = _zz_5322;
  assign _zz_5322 = ($signed(_zz_5323) >>> _zz_394);
  assign _zz_5323 = _zz_5324;
  assign _zz_5324 = ($signed(_zz_5326) - $signed(_zz_391));
  assign _zz_5325 = ({9'd0,data_mid_2_26_real} <<< 9);
  assign _zz_5326 = {{9{_zz_5325[26]}}, _zz_5325};
  assign _zz_5327 = fixTo_470_dout;
  assign _zz_5328 = _zz_5329[35 : 0];
  assign _zz_5329 = _zz_5330;
  assign _zz_5330 = ($signed(_zz_5331) >>> _zz_394);
  assign _zz_5331 = _zz_5332;
  assign _zz_5332 = ($signed(_zz_5334) - $signed(_zz_392));
  assign _zz_5333 = ({9'd0,data_mid_2_26_imag} <<< 9);
  assign _zz_5334 = {{9{_zz_5333[26]}}, _zz_5333};
  assign _zz_5335 = fixTo_471_dout;
  assign _zz_5336 = _zz_5337[35 : 0];
  assign _zz_5337 = _zz_5338;
  assign _zz_5338 = ($signed(_zz_5339) >>> _zz_395);
  assign _zz_5339 = _zz_5340;
  assign _zz_5340 = ($signed(_zz_5342) + $signed(_zz_391));
  assign _zz_5341 = ({9'd0,data_mid_2_26_real} <<< 9);
  assign _zz_5342 = {{9{_zz_5341[26]}}, _zz_5341};
  assign _zz_5343 = fixTo_472_dout;
  assign _zz_5344 = _zz_5345[35 : 0];
  assign _zz_5345 = _zz_5346;
  assign _zz_5346 = ($signed(_zz_5347) >>> _zz_395);
  assign _zz_5347 = _zz_5348;
  assign _zz_5348 = ($signed(_zz_5350) + $signed(_zz_392));
  assign _zz_5349 = ({9'd0,data_mid_2_26_imag} <<< 9);
  assign _zz_5350 = {{9{_zz_5349[26]}}, _zz_5349};
  assign _zz_5351 = fixTo_473_dout;
  assign _zz_5352 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_5353 = ($signed(_zz_398) - $signed(_zz_5354));
  assign _zz_5354 = ($signed(_zz_5355) * $signed(twiddle_factor_table_6_imag));
  assign _zz_5355 = ($signed(data_mid_2_31_real) + $signed(data_mid_2_31_imag));
  assign _zz_5356 = fixTo_474_dout;
  assign _zz_5357 = ($signed(_zz_398) + $signed(_zz_5358));
  assign _zz_5358 = ($signed(_zz_5359) * $signed(twiddle_factor_table_6_real));
  assign _zz_5359 = ($signed(data_mid_2_31_imag) - $signed(data_mid_2_31_real));
  assign _zz_5360 = fixTo_475_dout;
  assign _zz_5361 = _zz_5362[35 : 0];
  assign _zz_5362 = _zz_5363;
  assign _zz_5363 = ($signed(_zz_5364) >>> _zz_399);
  assign _zz_5364 = _zz_5365;
  assign _zz_5365 = ($signed(_zz_5367) - $signed(_zz_396));
  assign _zz_5366 = ({9'd0,data_mid_2_27_real} <<< 9);
  assign _zz_5367 = {{9{_zz_5366[26]}}, _zz_5366};
  assign _zz_5368 = fixTo_476_dout;
  assign _zz_5369 = _zz_5370[35 : 0];
  assign _zz_5370 = _zz_5371;
  assign _zz_5371 = ($signed(_zz_5372) >>> _zz_399);
  assign _zz_5372 = _zz_5373;
  assign _zz_5373 = ($signed(_zz_5375) - $signed(_zz_397));
  assign _zz_5374 = ({9'd0,data_mid_2_27_imag} <<< 9);
  assign _zz_5375 = {{9{_zz_5374[26]}}, _zz_5374};
  assign _zz_5376 = fixTo_477_dout;
  assign _zz_5377 = _zz_5378[35 : 0];
  assign _zz_5378 = _zz_5379;
  assign _zz_5379 = ($signed(_zz_5380) >>> _zz_400);
  assign _zz_5380 = _zz_5381;
  assign _zz_5381 = ($signed(_zz_5383) + $signed(_zz_396));
  assign _zz_5382 = ({9'd0,data_mid_2_27_real} <<< 9);
  assign _zz_5383 = {{9{_zz_5382[26]}}, _zz_5382};
  assign _zz_5384 = fixTo_478_dout;
  assign _zz_5385 = _zz_5386[35 : 0];
  assign _zz_5386 = _zz_5387;
  assign _zz_5387 = ($signed(_zz_5388) >>> _zz_400);
  assign _zz_5388 = _zz_5389;
  assign _zz_5389 = ($signed(_zz_5391) + $signed(_zz_397));
  assign _zz_5390 = ({9'd0,data_mid_2_27_imag} <<< 9);
  assign _zz_5391 = {{9{_zz_5390[26]}}, _zz_5390};
  assign _zz_5392 = fixTo_479_dout;
  assign _zz_5393 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_5394 = ($signed(_zz_403) - $signed(_zz_5395));
  assign _zz_5395 = ($signed(_zz_5396) * $signed(twiddle_factor_table_3_imag));
  assign _zz_5396 = ($signed(data_mid_2_36_real) + $signed(data_mid_2_36_imag));
  assign _zz_5397 = fixTo_480_dout;
  assign _zz_5398 = ($signed(_zz_403) + $signed(_zz_5399));
  assign _zz_5399 = ($signed(_zz_5400) * $signed(twiddle_factor_table_3_real));
  assign _zz_5400 = ($signed(data_mid_2_36_imag) - $signed(data_mid_2_36_real));
  assign _zz_5401 = fixTo_481_dout;
  assign _zz_5402 = _zz_5403[35 : 0];
  assign _zz_5403 = _zz_5404;
  assign _zz_5404 = ($signed(_zz_5405) >>> _zz_404);
  assign _zz_5405 = _zz_5406;
  assign _zz_5406 = ($signed(_zz_5408) - $signed(_zz_401));
  assign _zz_5407 = ({9'd0,data_mid_2_32_real} <<< 9);
  assign _zz_5408 = {{9{_zz_5407[26]}}, _zz_5407};
  assign _zz_5409 = fixTo_482_dout;
  assign _zz_5410 = _zz_5411[35 : 0];
  assign _zz_5411 = _zz_5412;
  assign _zz_5412 = ($signed(_zz_5413) >>> _zz_404);
  assign _zz_5413 = _zz_5414;
  assign _zz_5414 = ($signed(_zz_5416) - $signed(_zz_402));
  assign _zz_5415 = ({9'd0,data_mid_2_32_imag} <<< 9);
  assign _zz_5416 = {{9{_zz_5415[26]}}, _zz_5415};
  assign _zz_5417 = fixTo_483_dout;
  assign _zz_5418 = _zz_5419[35 : 0];
  assign _zz_5419 = _zz_5420;
  assign _zz_5420 = ($signed(_zz_5421) >>> _zz_405);
  assign _zz_5421 = _zz_5422;
  assign _zz_5422 = ($signed(_zz_5424) + $signed(_zz_401));
  assign _zz_5423 = ({9'd0,data_mid_2_32_real} <<< 9);
  assign _zz_5424 = {{9{_zz_5423[26]}}, _zz_5423};
  assign _zz_5425 = fixTo_484_dout;
  assign _zz_5426 = _zz_5427[35 : 0];
  assign _zz_5427 = _zz_5428;
  assign _zz_5428 = ($signed(_zz_5429) >>> _zz_405);
  assign _zz_5429 = _zz_5430;
  assign _zz_5430 = ($signed(_zz_5432) + $signed(_zz_402));
  assign _zz_5431 = ({9'd0,data_mid_2_32_imag} <<< 9);
  assign _zz_5432 = {{9{_zz_5431[26]}}, _zz_5431};
  assign _zz_5433 = fixTo_485_dout;
  assign _zz_5434 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_5435 = ($signed(_zz_408) - $signed(_zz_5436));
  assign _zz_5436 = ($signed(_zz_5437) * $signed(twiddle_factor_table_4_imag));
  assign _zz_5437 = ($signed(data_mid_2_37_real) + $signed(data_mid_2_37_imag));
  assign _zz_5438 = fixTo_486_dout;
  assign _zz_5439 = ($signed(_zz_408) + $signed(_zz_5440));
  assign _zz_5440 = ($signed(_zz_5441) * $signed(twiddle_factor_table_4_real));
  assign _zz_5441 = ($signed(data_mid_2_37_imag) - $signed(data_mid_2_37_real));
  assign _zz_5442 = fixTo_487_dout;
  assign _zz_5443 = _zz_5444[35 : 0];
  assign _zz_5444 = _zz_5445;
  assign _zz_5445 = ($signed(_zz_5446) >>> _zz_409);
  assign _zz_5446 = _zz_5447;
  assign _zz_5447 = ($signed(_zz_5449) - $signed(_zz_406));
  assign _zz_5448 = ({9'd0,data_mid_2_33_real} <<< 9);
  assign _zz_5449 = {{9{_zz_5448[26]}}, _zz_5448};
  assign _zz_5450 = fixTo_488_dout;
  assign _zz_5451 = _zz_5452[35 : 0];
  assign _zz_5452 = _zz_5453;
  assign _zz_5453 = ($signed(_zz_5454) >>> _zz_409);
  assign _zz_5454 = _zz_5455;
  assign _zz_5455 = ($signed(_zz_5457) - $signed(_zz_407));
  assign _zz_5456 = ({9'd0,data_mid_2_33_imag} <<< 9);
  assign _zz_5457 = {{9{_zz_5456[26]}}, _zz_5456};
  assign _zz_5458 = fixTo_489_dout;
  assign _zz_5459 = _zz_5460[35 : 0];
  assign _zz_5460 = _zz_5461;
  assign _zz_5461 = ($signed(_zz_5462) >>> _zz_410);
  assign _zz_5462 = _zz_5463;
  assign _zz_5463 = ($signed(_zz_5465) + $signed(_zz_406));
  assign _zz_5464 = ({9'd0,data_mid_2_33_real} <<< 9);
  assign _zz_5465 = {{9{_zz_5464[26]}}, _zz_5464};
  assign _zz_5466 = fixTo_490_dout;
  assign _zz_5467 = _zz_5468[35 : 0];
  assign _zz_5468 = _zz_5469;
  assign _zz_5469 = ($signed(_zz_5470) >>> _zz_410);
  assign _zz_5470 = _zz_5471;
  assign _zz_5471 = ($signed(_zz_5473) + $signed(_zz_407));
  assign _zz_5472 = ({9'd0,data_mid_2_33_imag} <<< 9);
  assign _zz_5473 = {{9{_zz_5472[26]}}, _zz_5472};
  assign _zz_5474 = fixTo_491_dout;
  assign _zz_5475 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_5476 = ($signed(_zz_413) - $signed(_zz_5477));
  assign _zz_5477 = ($signed(_zz_5478) * $signed(twiddle_factor_table_5_imag));
  assign _zz_5478 = ($signed(data_mid_2_38_real) + $signed(data_mid_2_38_imag));
  assign _zz_5479 = fixTo_492_dout;
  assign _zz_5480 = ($signed(_zz_413) + $signed(_zz_5481));
  assign _zz_5481 = ($signed(_zz_5482) * $signed(twiddle_factor_table_5_real));
  assign _zz_5482 = ($signed(data_mid_2_38_imag) - $signed(data_mid_2_38_real));
  assign _zz_5483 = fixTo_493_dout;
  assign _zz_5484 = _zz_5485[35 : 0];
  assign _zz_5485 = _zz_5486;
  assign _zz_5486 = ($signed(_zz_5487) >>> _zz_414);
  assign _zz_5487 = _zz_5488;
  assign _zz_5488 = ($signed(_zz_5490) - $signed(_zz_411));
  assign _zz_5489 = ({9'd0,data_mid_2_34_real} <<< 9);
  assign _zz_5490 = {{9{_zz_5489[26]}}, _zz_5489};
  assign _zz_5491 = fixTo_494_dout;
  assign _zz_5492 = _zz_5493[35 : 0];
  assign _zz_5493 = _zz_5494;
  assign _zz_5494 = ($signed(_zz_5495) >>> _zz_414);
  assign _zz_5495 = _zz_5496;
  assign _zz_5496 = ($signed(_zz_5498) - $signed(_zz_412));
  assign _zz_5497 = ({9'd0,data_mid_2_34_imag} <<< 9);
  assign _zz_5498 = {{9{_zz_5497[26]}}, _zz_5497};
  assign _zz_5499 = fixTo_495_dout;
  assign _zz_5500 = _zz_5501[35 : 0];
  assign _zz_5501 = _zz_5502;
  assign _zz_5502 = ($signed(_zz_5503) >>> _zz_415);
  assign _zz_5503 = _zz_5504;
  assign _zz_5504 = ($signed(_zz_5506) + $signed(_zz_411));
  assign _zz_5505 = ({9'd0,data_mid_2_34_real} <<< 9);
  assign _zz_5506 = {{9{_zz_5505[26]}}, _zz_5505};
  assign _zz_5507 = fixTo_496_dout;
  assign _zz_5508 = _zz_5509[35 : 0];
  assign _zz_5509 = _zz_5510;
  assign _zz_5510 = ($signed(_zz_5511) >>> _zz_415);
  assign _zz_5511 = _zz_5512;
  assign _zz_5512 = ($signed(_zz_5514) + $signed(_zz_412));
  assign _zz_5513 = ({9'd0,data_mid_2_34_imag} <<< 9);
  assign _zz_5514 = {{9{_zz_5513[26]}}, _zz_5513};
  assign _zz_5515 = fixTo_497_dout;
  assign _zz_5516 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_5517 = ($signed(_zz_418) - $signed(_zz_5518));
  assign _zz_5518 = ($signed(_zz_5519) * $signed(twiddle_factor_table_6_imag));
  assign _zz_5519 = ($signed(data_mid_2_39_real) + $signed(data_mid_2_39_imag));
  assign _zz_5520 = fixTo_498_dout;
  assign _zz_5521 = ($signed(_zz_418) + $signed(_zz_5522));
  assign _zz_5522 = ($signed(_zz_5523) * $signed(twiddle_factor_table_6_real));
  assign _zz_5523 = ($signed(data_mid_2_39_imag) - $signed(data_mid_2_39_real));
  assign _zz_5524 = fixTo_499_dout;
  assign _zz_5525 = _zz_5526[35 : 0];
  assign _zz_5526 = _zz_5527;
  assign _zz_5527 = ($signed(_zz_5528) >>> _zz_419);
  assign _zz_5528 = _zz_5529;
  assign _zz_5529 = ($signed(_zz_5531) - $signed(_zz_416));
  assign _zz_5530 = ({9'd0,data_mid_2_35_real} <<< 9);
  assign _zz_5531 = {{9{_zz_5530[26]}}, _zz_5530};
  assign _zz_5532 = fixTo_500_dout;
  assign _zz_5533 = _zz_5534[35 : 0];
  assign _zz_5534 = _zz_5535;
  assign _zz_5535 = ($signed(_zz_5536) >>> _zz_419);
  assign _zz_5536 = _zz_5537;
  assign _zz_5537 = ($signed(_zz_5539) - $signed(_zz_417));
  assign _zz_5538 = ({9'd0,data_mid_2_35_imag} <<< 9);
  assign _zz_5539 = {{9{_zz_5538[26]}}, _zz_5538};
  assign _zz_5540 = fixTo_501_dout;
  assign _zz_5541 = _zz_5542[35 : 0];
  assign _zz_5542 = _zz_5543;
  assign _zz_5543 = ($signed(_zz_5544) >>> _zz_420);
  assign _zz_5544 = _zz_5545;
  assign _zz_5545 = ($signed(_zz_5547) + $signed(_zz_416));
  assign _zz_5546 = ({9'd0,data_mid_2_35_real} <<< 9);
  assign _zz_5547 = {{9{_zz_5546[26]}}, _zz_5546};
  assign _zz_5548 = fixTo_502_dout;
  assign _zz_5549 = _zz_5550[35 : 0];
  assign _zz_5550 = _zz_5551;
  assign _zz_5551 = ($signed(_zz_5552) >>> _zz_420);
  assign _zz_5552 = _zz_5553;
  assign _zz_5553 = ($signed(_zz_5555) + $signed(_zz_417));
  assign _zz_5554 = ({9'd0,data_mid_2_35_imag} <<< 9);
  assign _zz_5555 = {{9{_zz_5554[26]}}, _zz_5554};
  assign _zz_5556 = fixTo_503_dout;
  assign _zz_5557 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_5558 = ($signed(_zz_423) - $signed(_zz_5559));
  assign _zz_5559 = ($signed(_zz_5560) * $signed(twiddle_factor_table_3_imag));
  assign _zz_5560 = ($signed(data_mid_2_44_real) + $signed(data_mid_2_44_imag));
  assign _zz_5561 = fixTo_504_dout;
  assign _zz_5562 = ($signed(_zz_423) + $signed(_zz_5563));
  assign _zz_5563 = ($signed(_zz_5564) * $signed(twiddle_factor_table_3_real));
  assign _zz_5564 = ($signed(data_mid_2_44_imag) - $signed(data_mid_2_44_real));
  assign _zz_5565 = fixTo_505_dout;
  assign _zz_5566 = _zz_5567[35 : 0];
  assign _zz_5567 = _zz_5568;
  assign _zz_5568 = ($signed(_zz_5569) >>> _zz_424);
  assign _zz_5569 = _zz_5570;
  assign _zz_5570 = ($signed(_zz_5572) - $signed(_zz_421));
  assign _zz_5571 = ({9'd0,data_mid_2_40_real} <<< 9);
  assign _zz_5572 = {{9{_zz_5571[26]}}, _zz_5571};
  assign _zz_5573 = fixTo_506_dout;
  assign _zz_5574 = _zz_5575[35 : 0];
  assign _zz_5575 = _zz_5576;
  assign _zz_5576 = ($signed(_zz_5577) >>> _zz_424);
  assign _zz_5577 = _zz_5578;
  assign _zz_5578 = ($signed(_zz_5580) - $signed(_zz_422));
  assign _zz_5579 = ({9'd0,data_mid_2_40_imag} <<< 9);
  assign _zz_5580 = {{9{_zz_5579[26]}}, _zz_5579};
  assign _zz_5581 = fixTo_507_dout;
  assign _zz_5582 = _zz_5583[35 : 0];
  assign _zz_5583 = _zz_5584;
  assign _zz_5584 = ($signed(_zz_5585) >>> _zz_425);
  assign _zz_5585 = _zz_5586;
  assign _zz_5586 = ($signed(_zz_5588) + $signed(_zz_421));
  assign _zz_5587 = ({9'd0,data_mid_2_40_real} <<< 9);
  assign _zz_5588 = {{9{_zz_5587[26]}}, _zz_5587};
  assign _zz_5589 = fixTo_508_dout;
  assign _zz_5590 = _zz_5591[35 : 0];
  assign _zz_5591 = _zz_5592;
  assign _zz_5592 = ($signed(_zz_5593) >>> _zz_425);
  assign _zz_5593 = _zz_5594;
  assign _zz_5594 = ($signed(_zz_5596) + $signed(_zz_422));
  assign _zz_5595 = ({9'd0,data_mid_2_40_imag} <<< 9);
  assign _zz_5596 = {{9{_zz_5595[26]}}, _zz_5595};
  assign _zz_5597 = fixTo_509_dout;
  assign _zz_5598 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_5599 = ($signed(_zz_428) - $signed(_zz_5600));
  assign _zz_5600 = ($signed(_zz_5601) * $signed(twiddle_factor_table_4_imag));
  assign _zz_5601 = ($signed(data_mid_2_45_real) + $signed(data_mid_2_45_imag));
  assign _zz_5602 = fixTo_510_dout;
  assign _zz_5603 = ($signed(_zz_428) + $signed(_zz_5604));
  assign _zz_5604 = ($signed(_zz_5605) * $signed(twiddle_factor_table_4_real));
  assign _zz_5605 = ($signed(data_mid_2_45_imag) - $signed(data_mid_2_45_real));
  assign _zz_5606 = fixTo_511_dout;
  assign _zz_5607 = _zz_5608[35 : 0];
  assign _zz_5608 = _zz_5609;
  assign _zz_5609 = ($signed(_zz_5610) >>> _zz_429);
  assign _zz_5610 = _zz_5611;
  assign _zz_5611 = ($signed(_zz_5613) - $signed(_zz_426));
  assign _zz_5612 = ({9'd0,data_mid_2_41_real} <<< 9);
  assign _zz_5613 = {{9{_zz_5612[26]}}, _zz_5612};
  assign _zz_5614 = fixTo_512_dout;
  assign _zz_5615 = _zz_5616[35 : 0];
  assign _zz_5616 = _zz_5617;
  assign _zz_5617 = ($signed(_zz_5618) >>> _zz_429);
  assign _zz_5618 = _zz_5619;
  assign _zz_5619 = ($signed(_zz_5621) - $signed(_zz_427));
  assign _zz_5620 = ({9'd0,data_mid_2_41_imag} <<< 9);
  assign _zz_5621 = {{9{_zz_5620[26]}}, _zz_5620};
  assign _zz_5622 = fixTo_513_dout;
  assign _zz_5623 = _zz_5624[35 : 0];
  assign _zz_5624 = _zz_5625;
  assign _zz_5625 = ($signed(_zz_5626) >>> _zz_430);
  assign _zz_5626 = _zz_5627;
  assign _zz_5627 = ($signed(_zz_5629) + $signed(_zz_426));
  assign _zz_5628 = ({9'd0,data_mid_2_41_real} <<< 9);
  assign _zz_5629 = {{9{_zz_5628[26]}}, _zz_5628};
  assign _zz_5630 = fixTo_514_dout;
  assign _zz_5631 = _zz_5632[35 : 0];
  assign _zz_5632 = _zz_5633;
  assign _zz_5633 = ($signed(_zz_5634) >>> _zz_430);
  assign _zz_5634 = _zz_5635;
  assign _zz_5635 = ($signed(_zz_5637) + $signed(_zz_427));
  assign _zz_5636 = ({9'd0,data_mid_2_41_imag} <<< 9);
  assign _zz_5637 = {{9{_zz_5636[26]}}, _zz_5636};
  assign _zz_5638 = fixTo_515_dout;
  assign _zz_5639 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_5640 = ($signed(_zz_433) - $signed(_zz_5641));
  assign _zz_5641 = ($signed(_zz_5642) * $signed(twiddle_factor_table_5_imag));
  assign _zz_5642 = ($signed(data_mid_2_46_real) + $signed(data_mid_2_46_imag));
  assign _zz_5643 = fixTo_516_dout;
  assign _zz_5644 = ($signed(_zz_433) + $signed(_zz_5645));
  assign _zz_5645 = ($signed(_zz_5646) * $signed(twiddle_factor_table_5_real));
  assign _zz_5646 = ($signed(data_mid_2_46_imag) - $signed(data_mid_2_46_real));
  assign _zz_5647 = fixTo_517_dout;
  assign _zz_5648 = _zz_5649[35 : 0];
  assign _zz_5649 = _zz_5650;
  assign _zz_5650 = ($signed(_zz_5651) >>> _zz_434);
  assign _zz_5651 = _zz_5652;
  assign _zz_5652 = ($signed(_zz_5654) - $signed(_zz_431));
  assign _zz_5653 = ({9'd0,data_mid_2_42_real} <<< 9);
  assign _zz_5654 = {{9{_zz_5653[26]}}, _zz_5653};
  assign _zz_5655 = fixTo_518_dout;
  assign _zz_5656 = _zz_5657[35 : 0];
  assign _zz_5657 = _zz_5658;
  assign _zz_5658 = ($signed(_zz_5659) >>> _zz_434);
  assign _zz_5659 = _zz_5660;
  assign _zz_5660 = ($signed(_zz_5662) - $signed(_zz_432));
  assign _zz_5661 = ({9'd0,data_mid_2_42_imag} <<< 9);
  assign _zz_5662 = {{9{_zz_5661[26]}}, _zz_5661};
  assign _zz_5663 = fixTo_519_dout;
  assign _zz_5664 = _zz_5665[35 : 0];
  assign _zz_5665 = _zz_5666;
  assign _zz_5666 = ($signed(_zz_5667) >>> _zz_435);
  assign _zz_5667 = _zz_5668;
  assign _zz_5668 = ($signed(_zz_5670) + $signed(_zz_431));
  assign _zz_5669 = ({9'd0,data_mid_2_42_real} <<< 9);
  assign _zz_5670 = {{9{_zz_5669[26]}}, _zz_5669};
  assign _zz_5671 = fixTo_520_dout;
  assign _zz_5672 = _zz_5673[35 : 0];
  assign _zz_5673 = _zz_5674;
  assign _zz_5674 = ($signed(_zz_5675) >>> _zz_435);
  assign _zz_5675 = _zz_5676;
  assign _zz_5676 = ($signed(_zz_5678) + $signed(_zz_432));
  assign _zz_5677 = ({9'd0,data_mid_2_42_imag} <<< 9);
  assign _zz_5678 = {{9{_zz_5677[26]}}, _zz_5677};
  assign _zz_5679 = fixTo_521_dout;
  assign _zz_5680 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_5681 = ($signed(_zz_438) - $signed(_zz_5682));
  assign _zz_5682 = ($signed(_zz_5683) * $signed(twiddle_factor_table_6_imag));
  assign _zz_5683 = ($signed(data_mid_2_47_real) + $signed(data_mid_2_47_imag));
  assign _zz_5684 = fixTo_522_dout;
  assign _zz_5685 = ($signed(_zz_438) + $signed(_zz_5686));
  assign _zz_5686 = ($signed(_zz_5687) * $signed(twiddle_factor_table_6_real));
  assign _zz_5687 = ($signed(data_mid_2_47_imag) - $signed(data_mid_2_47_real));
  assign _zz_5688 = fixTo_523_dout;
  assign _zz_5689 = _zz_5690[35 : 0];
  assign _zz_5690 = _zz_5691;
  assign _zz_5691 = ($signed(_zz_5692) >>> _zz_439);
  assign _zz_5692 = _zz_5693;
  assign _zz_5693 = ($signed(_zz_5695) - $signed(_zz_436));
  assign _zz_5694 = ({9'd0,data_mid_2_43_real} <<< 9);
  assign _zz_5695 = {{9{_zz_5694[26]}}, _zz_5694};
  assign _zz_5696 = fixTo_524_dout;
  assign _zz_5697 = _zz_5698[35 : 0];
  assign _zz_5698 = _zz_5699;
  assign _zz_5699 = ($signed(_zz_5700) >>> _zz_439);
  assign _zz_5700 = _zz_5701;
  assign _zz_5701 = ($signed(_zz_5703) - $signed(_zz_437));
  assign _zz_5702 = ({9'd0,data_mid_2_43_imag} <<< 9);
  assign _zz_5703 = {{9{_zz_5702[26]}}, _zz_5702};
  assign _zz_5704 = fixTo_525_dout;
  assign _zz_5705 = _zz_5706[35 : 0];
  assign _zz_5706 = _zz_5707;
  assign _zz_5707 = ($signed(_zz_5708) >>> _zz_440);
  assign _zz_5708 = _zz_5709;
  assign _zz_5709 = ($signed(_zz_5711) + $signed(_zz_436));
  assign _zz_5710 = ({9'd0,data_mid_2_43_real} <<< 9);
  assign _zz_5711 = {{9{_zz_5710[26]}}, _zz_5710};
  assign _zz_5712 = fixTo_526_dout;
  assign _zz_5713 = _zz_5714[35 : 0];
  assign _zz_5714 = _zz_5715;
  assign _zz_5715 = ($signed(_zz_5716) >>> _zz_440);
  assign _zz_5716 = _zz_5717;
  assign _zz_5717 = ($signed(_zz_5719) + $signed(_zz_437));
  assign _zz_5718 = ({9'd0,data_mid_2_43_imag} <<< 9);
  assign _zz_5719 = {{9{_zz_5718[26]}}, _zz_5718};
  assign _zz_5720 = fixTo_527_dout;
  assign _zz_5721 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_5722 = ($signed(_zz_443) - $signed(_zz_5723));
  assign _zz_5723 = ($signed(_zz_5724) * $signed(twiddle_factor_table_3_imag));
  assign _zz_5724 = ($signed(data_mid_2_52_real) + $signed(data_mid_2_52_imag));
  assign _zz_5725 = fixTo_528_dout;
  assign _zz_5726 = ($signed(_zz_443) + $signed(_zz_5727));
  assign _zz_5727 = ($signed(_zz_5728) * $signed(twiddle_factor_table_3_real));
  assign _zz_5728 = ($signed(data_mid_2_52_imag) - $signed(data_mid_2_52_real));
  assign _zz_5729 = fixTo_529_dout;
  assign _zz_5730 = _zz_5731[35 : 0];
  assign _zz_5731 = _zz_5732;
  assign _zz_5732 = ($signed(_zz_5733) >>> _zz_444);
  assign _zz_5733 = _zz_5734;
  assign _zz_5734 = ($signed(_zz_5736) - $signed(_zz_441));
  assign _zz_5735 = ({9'd0,data_mid_2_48_real} <<< 9);
  assign _zz_5736 = {{9{_zz_5735[26]}}, _zz_5735};
  assign _zz_5737 = fixTo_530_dout;
  assign _zz_5738 = _zz_5739[35 : 0];
  assign _zz_5739 = _zz_5740;
  assign _zz_5740 = ($signed(_zz_5741) >>> _zz_444);
  assign _zz_5741 = _zz_5742;
  assign _zz_5742 = ($signed(_zz_5744) - $signed(_zz_442));
  assign _zz_5743 = ({9'd0,data_mid_2_48_imag} <<< 9);
  assign _zz_5744 = {{9{_zz_5743[26]}}, _zz_5743};
  assign _zz_5745 = fixTo_531_dout;
  assign _zz_5746 = _zz_5747[35 : 0];
  assign _zz_5747 = _zz_5748;
  assign _zz_5748 = ($signed(_zz_5749) >>> _zz_445);
  assign _zz_5749 = _zz_5750;
  assign _zz_5750 = ($signed(_zz_5752) + $signed(_zz_441));
  assign _zz_5751 = ({9'd0,data_mid_2_48_real} <<< 9);
  assign _zz_5752 = {{9{_zz_5751[26]}}, _zz_5751};
  assign _zz_5753 = fixTo_532_dout;
  assign _zz_5754 = _zz_5755[35 : 0];
  assign _zz_5755 = _zz_5756;
  assign _zz_5756 = ($signed(_zz_5757) >>> _zz_445);
  assign _zz_5757 = _zz_5758;
  assign _zz_5758 = ($signed(_zz_5760) + $signed(_zz_442));
  assign _zz_5759 = ({9'd0,data_mid_2_48_imag} <<< 9);
  assign _zz_5760 = {{9{_zz_5759[26]}}, _zz_5759};
  assign _zz_5761 = fixTo_533_dout;
  assign _zz_5762 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_5763 = ($signed(_zz_448) - $signed(_zz_5764));
  assign _zz_5764 = ($signed(_zz_5765) * $signed(twiddle_factor_table_4_imag));
  assign _zz_5765 = ($signed(data_mid_2_53_real) + $signed(data_mid_2_53_imag));
  assign _zz_5766 = fixTo_534_dout;
  assign _zz_5767 = ($signed(_zz_448) + $signed(_zz_5768));
  assign _zz_5768 = ($signed(_zz_5769) * $signed(twiddle_factor_table_4_real));
  assign _zz_5769 = ($signed(data_mid_2_53_imag) - $signed(data_mid_2_53_real));
  assign _zz_5770 = fixTo_535_dout;
  assign _zz_5771 = _zz_5772[35 : 0];
  assign _zz_5772 = _zz_5773;
  assign _zz_5773 = ($signed(_zz_5774) >>> _zz_449);
  assign _zz_5774 = _zz_5775;
  assign _zz_5775 = ($signed(_zz_5777) - $signed(_zz_446));
  assign _zz_5776 = ({9'd0,data_mid_2_49_real} <<< 9);
  assign _zz_5777 = {{9{_zz_5776[26]}}, _zz_5776};
  assign _zz_5778 = fixTo_536_dout;
  assign _zz_5779 = _zz_5780[35 : 0];
  assign _zz_5780 = _zz_5781;
  assign _zz_5781 = ($signed(_zz_5782) >>> _zz_449);
  assign _zz_5782 = _zz_5783;
  assign _zz_5783 = ($signed(_zz_5785) - $signed(_zz_447));
  assign _zz_5784 = ({9'd0,data_mid_2_49_imag} <<< 9);
  assign _zz_5785 = {{9{_zz_5784[26]}}, _zz_5784};
  assign _zz_5786 = fixTo_537_dout;
  assign _zz_5787 = _zz_5788[35 : 0];
  assign _zz_5788 = _zz_5789;
  assign _zz_5789 = ($signed(_zz_5790) >>> _zz_450);
  assign _zz_5790 = _zz_5791;
  assign _zz_5791 = ($signed(_zz_5793) + $signed(_zz_446));
  assign _zz_5792 = ({9'd0,data_mid_2_49_real} <<< 9);
  assign _zz_5793 = {{9{_zz_5792[26]}}, _zz_5792};
  assign _zz_5794 = fixTo_538_dout;
  assign _zz_5795 = _zz_5796[35 : 0];
  assign _zz_5796 = _zz_5797;
  assign _zz_5797 = ($signed(_zz_5798) >>> _zz_450);
  assign _zz_5798 = _zz_5799;
  assign _zz_5799 = ($signed(_zz_5801) + $signed(_zz_447));
  assign _zz_5800 = ({9'd0,data_mid_2_49_imag} <<< 9);
  assign _zz_5801 = {{9{_zz_5800[26]}}, _zz_5800};
  assign _zz_5802 = fixTo_539_dout;
  assign _zz_5803 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_5804 = ($signed(_zz_453) - $signed(_zz_5805));
  assign _zz_5805 = ($signed(_zz_5806) * $signed(twiddle_factor_table_5_imag));
  assign _zz_5806 = ($signed(data_mid_2_54_real) + $signed(data_mid_2_54_imag));
  assign _zz_5807 = fixTo_540_dout;
  assign _zz_5808 = ($signed(_zz_453) + $signed(_zz_5809));
  assign _zz_5809 = ($signed(_zz_5810) * $signed(twiddle_factor_table_5_real));
  assign _zz_5810 = ($signed(data_mid_2_54_imag) - $signed(data_mid_2_54_real));
  assign _zz_5811 = fixTo_541_dout;
  assign _zz_5812 = _zz_5813[35 : 0];
  assign _zz_5813 = _zz_5814;
  assign _zz_5814 = ($signed(_zz_5815) >>> _zz_454);
  assign _zz_5815 = _zz_5816;
  assign _zz_5816 = ($signed(_zz_5818) - $signed(_zz_451));
  assign _zz_5817 = ({9'd0,data_mid_2_50_real} <<< 9);
  assign _zz_5818 = {{9{_zz_5817[26]}}, _zz_5817};
  assign _zz_5819 = fixTo_542_dout;
  assign _zz_5820 = _zz_5821[35 : 0];
  assign _zz_5821 = _zz_5822;
  assign _zz_5822 = ($signed(_zz_5823) >>> _zz_454);
  assign _zz_5823 = _zz_5824;
  assign _zz_5824 = ($signed(_zz_5826) - $signed(_zz_452));
  assign _zz_5825 = ({9'd0,data_mid_2_50_imag} <<< 9);
  assign _zz_5826 = {{9{_zz_5825[26]}}, _zz_5825};
  assign _zz_5827 = fixTo_543_dout;
  assign _zz_5828 = _zz_5829[35 : 0];
  assign _zz_5829 = _zz_5830;
  assign _zz_5830 = ($signed(_zz_5831) >>> _zz_455);
  assign _zz_5831 = _zz_5832;
  assign _zz_5832 = ($signed(_zz_5834) + $signed(_zz_451));
  assign _zz_5833 = ({9'd0,data_mid_2_50_real} <<< 9);
  assign _zz_5834 = {{9{_zz_5833[26]}}, _zz_5833};
  assign _zz_5835 = fixTo_544_dout;
  assign _zz_5836 = _zz_5837[35 : 0];
  assign _zz_5837 = _zz_5838;
  assign _zz_5838 = ($signed(_zz_5839) >>> _zz_455);
  assign _zz_5839 = _zz_5840;
  assign _zz_5840 = ($signed(_zz_5842) + $signed(_zz_452));
  assign _zz_5841 = ({9'd0,data_mid_2_50_imag} <<< 9);
  assign _zz_5842 = {{9{_zz_5841[26]}}, _zz_5841};
  assign _zz_5843 = fixTo_545_dout;
  assign _zz_5844 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_5845 = ($signed(_zz_458) - $signed(_zz_5846));
  assign _zz_5846 = ($signed(_zz_5847) * $signed(twiddle_factor_table_6_imag));
  assign _zz_5847 = ($signed(data_mid_2_55_real) + $signed(data_mid_2_55_imag));
  assign _zz_5848 = fixTo_546_dout;
  assign _zz_5849 = ($signed(_zz_458) + $signed(_zz_5850));
  assign _zz_5850 = ($signed(_zz_5851) * $signed(twiddle_factor_table_6_real));
  assign _zz_5851 = ($signed(data_mid_2_55_imag) - $signed(data_mid_2_55_real));
  assign _zz_5852 = fixTo_547_dout;
  assign _zz_5853 = _zz_5854[35 : 0];
  assign _zz_5854 = _zz_5855;
  assign _zz_5855 = ($signed(_zz_5856) >>> _zz_459);
  assign _zz_5856 = _zz_5857;
  assign _zz_5857 = ($signed(_zz_5859) - $signed(_zz_456));
  assign _zz_5858 = ({9'd0,data_mid_2_51_real} <<< 9);
  assign _zz_5859 = {{9{_zz_5858[26]}}, _zz_5858};
  assign _zz_5860 = fixTo_548_dout;
  assign _zz_5861 = _zz_5862[35 : 0];
  assign _zz_5862 = _zz_5863;
  assign _zz_5863 = ($signed(_zz_5864) >>> _zz_459);
  assign _zz_5864 = _zz_5865;
  assign _zz_5865 = ($signed(_zz_5867) - $signed(_zz_457));
  assign _zz_5866 = ({9'd0,data_mid_2_51_imag} <<< 9);
  assign _zz_5867 = {{9{_zz_5866[26]}}, _zz_5866};
  assign _zz_5868 = fixTo_549_dout;
  assign _zz_5869 = _zz_5870[35 : 0];
  assign _zz_5870 = _zz_5871;
  assign _zz_5871 = ($signed(_zz_5872) >>> _zz_460);
  assign _zz_5872 = _zz_5873;
  assign _zz_5873 = ($signed(_zz_5875) + $signed(_zz_456));
  assign _zz_5874 = ({9'd0,data_mid_2_51_real} <<< 9);
  assign _zz_5875 = {{9{_zz_5874[26]}}, _zz_5874};
  assign _zz_5876 = fixTo_550_dout;
  assign _zz_5877 = _zz_5878[35 : 0];
  assign _zz_5878 = _zz_5879;
  assign _zz_5879 = ($signed(_zz_5880) >>> _zz_460);
  assign _zz_5880 = _zz_5881;
  assign _zz_5881 = ($signed(_zz_5883) + $signed(_zz_457));
  assign _zz_5882 = ({9'd0,data_mid_2_51_imag} <<< 9);
  assign _zz_5883 = {{9{_zz_5882[26]}}, _zz_5882};
  assign _zz_5884 = fixTo_551_dout;
  assign _zz_5885 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_5886 = ($signed(_zz_463) - $signed(_zz_5887));
  assign _zz_5887 = ($signed(_zz_5888) * $signed(twiddle_factor_table_3_imag));
  assign _zz_5888 = ($signed(data_mid_2_60_real) + $signed(data_mid_2_60_imag));
  assign _zz_5889 = fixTo_552_dout;
  assign _zz_5890 = ($signed(_zz_463) + $signed(_zz_5891));
  assign _zz_5891 = ($signed(_zz_5892) * $signed(twiddle_factor_table_3_real));
  assign _zz_5892 = ($signed(data_mid_2_60_imag) - $signed(data_mid_2_60_real));
  assign _zz_5893 = fixTo_553_dout;
  assign _zz_5894 = _zz_5895[35 : 0];
  assign _zz_5895 = _zz_5896;
  assign _zz_5896 = ($signed(_zz_5897) >>> _zz_464);
  assign _zz_5897 = _zz_5898;
  assign _zz_5898 = ($signed(_zz_5900) - $signed(_zz_461));
  assign _zz_5899 = ({9'd0,data_mid_2_56_real} <<< 9);
  assign _zz_5900 = {{9{_zz_5899[26]}}, _zz_5899};
  assign _zz_5901 = fixTo_554_dout;
  assign _zz_5902 = _zz_5903[35 : 0];
  assign _zz_5903 = _zz_5904;
  assign _zz_5904 = ($signed(_zz_5905) >>> _zz_464);
  assign _zz_5905 = _zz_5906;
  assign _zz_5906 = ($signed(_zz_5908) - $signed(_zz_462));
  assign _zz_5907 = ({9'd0,data_mid_2_56_imag} <<< 9);
  assign _zz_5908 = {{9{_zz_5907[26]}}, _zz_5907};
  assign _zz_5909 = fixTo_555_dout;
  assign _zz_5910 = _zz_5911[35 : 0];
  assign _zz_5911 = _zz_5912;
  assign _zz_5912 = ($signed(_zz_5913) >>> _zz_465);
  assign _zz_5913 = _zz_5914;
  assign _zz_5914 = ($signed(_zz_5916) + $signed(_zz_461));
  assign _zz_5915 = ({9'd0,data_mid_2_56_real} <<< 9);
  assign _zz_5916 = {{9{_zz_5915[26]}}, _zz_5915};
  assign _zz_5917 = fixTo_556_dout;
  assign _zz_5918 = _zz_5919[35 : 0];
  assign _zz_5919 = _zz_5920;
  assign _zz_5920 = ($signed(_zz_5921) >>> _zz_465);
  assign _zz_5921 = _zz_5922;
  assign _zz_5922 = ($signed(_zz_5924) + $signed(_zz_462));
  assign _zz_5923 = ({9'd0,data_mid_2_56_imag} <<< 9);
  assign _zz_5924 = {{9{_zz_5923[26]}}, _zz_5923};
  assign _zz_5925 = fixTo_557_dout;
  assign _zz_5926 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_5927 = ($signed(_zz_468) - $signed(_zz_5928));
  assign _zz_5928 = ($signed(_zz_5929) * $signed(twiddle_factor_table_4_imag));
  assign _zz_5929 = ($signed(data_mid_2_61_real) + $signed(data_mid_2_61_imag));
  assign _zz_5930 = fixTo_558_dout;
  assign _zz_5931 = ($signed(_zz_468) + $signed(_zz_5932));
  assign _zz_5932 = ($signed(_zz_5933) * $signed(twiddle_factor_table_4_real));
  assign _zz_5933 = ($signed(data_mid_2_61_imag) - $signed(data_mid_2_61_real));
  assign _zz_5934 = fixTo_559_dout;
  assign _zz_5935 = _zz_5936[35 : 0];
  assign _zz_5936 = _zz_5937;
  assign _zz_5937 = ($signed(_zz_5938) >>> _zz_469);
  assign _zz_5938 = _zz_5939;
  assign _zz_5939 = ($signed(_zz_5941) - $signed(_zz_466));
  assign _zz_5940 = ({9'd0,data_mid_2_57_real} <<< 9);
  assign _zz_5941 = {{9{_zz_5940[26]}}, _zz_5940};
  assign _zz_5942 = fixTo_560_dout;
  assign _zz_5943 = _zz_5944[35 : 0];
  assign _zz_5944 = _zz_5945;
  assign _zz_5945 = ($signed(_zz_5946) >>> _zz_469);
  assign _zz_5946 = _zz_5947;
  assign _zz_5947 = ($signed(_zz_5949) - $signed(_zz_467));
  assign _zz_5948 = ({9'd0,data_mid_2_57_imag} <<< 9);
  assign _zz_5949 = {{9{_zz_5948[26]}}, _zz_5948};
  assign _zz_5950 = fixTo_561_dout;
  assign _zz_5951 = _zz_5952[35 : 0];
  assign _zz_5952 = _zz_5953;
  assign _zz_5953 = ($signed(_zz_5954) >>> _zz_470);
  assign _zz_5954 = _zz_5955;
  assign _zz_5955 = ($signed(_zz_5957) + $signed(_zz_466));
  assign _zz_5956 = ({9'd0,data_mid_2_57_real} <<< 9);
  assign _zz_5957 = {{9{_zz_5956[26]}}, _zz_5956};
  assign _zz_5958 = fixTo_562_dout;
  assign _zz_5959 = _zz_5960[35 : 0];
  assign _zz_5960 = _zz_5961;
  assign _zz_5961 = ($signed(_zz_5962) >>> _zz_470);
  assign _zz_5962 = _zz_5963;
  assign _zz_5963 = ($signed(_zz_5965) + $signed(_zz_467));
  assign _zz_5964 = ({9'd0,data_mid_2_57_imag} <<< 9);
  assign _zz_5965 = {{9{_zz_5964[26]}}, _zz_5964};
  assign _zz_5966 = fixTo_563_dout;
  assign _zz_5967 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_5968 = ($signed(_zz_473) - $signed(_zz_5969));
  assign _zz_5969 = ($signed(_zz_5970) * $signed(twiddle_factor_table_5_imag));
  assign _zz_5970 = ($signed(data_mid_2_62_real) + $signed(data_mid_2_62_imag));
  assign _zz_5971 = fixTo_564_dout;
  assign _zz_5972 = ($signed(_zz_473) + $signed(_zz_5973));
  assign _zz_5973 = ($signed(_zz_5974) * $signed(twiddle_factor_table_5_real));
  assign _zz_5974 = ($signed(data_mid_2_62_imag) - $signed(data_mid_2_62_real));
  assign _zz_5975 = fixTo_565_dout;
  assign _zz_5976 = _zz_5977[35 : 0];
  assign _zz_5977 = _zz_5978;
  assign _zz_5978 = ($signed(_zz_5979) >>> _zz_474);
  assign _zz_5979 = _zz_5980;
  assign _zz_5980 = ($signed(_zz_5982) - $signed(_zz_471));
  assign _zz_5981 = ({9'd0,data_mid_2_58_real} <<< 9);
  assign _zz_5982 = {{9{_zz_5981[26]}}, _zz_5981};
  assign _zz_5983 = fixTo_566_dout;
  assign _zz_5984 = _zz_5985[35 : 0];
  assign _zz_5985 = _zz_5986;
  assign _zz_5986 = ($signed(_zz_5987) >>> _zz_474);
  assign _zz_5987 = _zz_5988;
  assign _zz_5988 = ($signed(_zz_5990) - $signed(_zz_472));
  assign _zz_5989 = ({9'd0,data_mid_2_58_imag} <<< 9);
  assign _zz_5990 = {{9{_zz_5989[26]}}, _zz_5989};
  assign _zz_5991 = fixTo_567_dout;
  assign _zz_5992 = _zz_5993[35 : 0];
  assign _zz_5993 = _zz_5994;
  assign _zz_5994 = ($signed(_zz_5995) >>> _zz_475);
  assign _zz_5995 = _zz_5996;
  assign _zz_5996 = ($signed(_zz_5998) + $signed(_zz_471));
  assign _zz_5997 = ({9'd0,data_mid_2_58_real} <<< 9);
  assign _zz_5998 = {{9{_zz_5997[26]}}, _zz_5997};
  assign _zz_5999 = fixTo_568_dout;
  assign _zz_6000 = _zz_6001[35 : 0];
  assign _zz_6001 = _zz_6002;
  assign _zz_6002 = ($signed(_zz_6003) >>> _zz_475);
  assign _zz_6003 = _zz_6004;
  assign _zz_6004 = ($signed(_zz_6006) + $signed(_zz_472));
  assign _zz_6005 = ({9'd0,data_mid_2_58_imag} <<< 9);
  assign _zz_6006 = {{9{_zz_6005[26]}}, _zz_6005};
  assign _zz_6007 = fixTo_569_dout;
  assign _zz_6008 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_6009 = ($signed(_zz_478) - $signed(_zz_6010));
  assign _zz_6010 = ($signed(_zz_6011) * $signed(twiddle_factor_table_6_imag));
  assign _zz_6011 = ($signed(data_mid_2_63_real) + $signed(data_mid_2_63_imag));
  assign _zz_6012 = fixTo_570_dout;
  assign _zz_6013 = ($signed(_zz_478) + $signed(_zz_6014));
  assign _zz_6014 = ($signed(_zz_6015) * $signed(twiddle_factor_table_6_real));
  assign _zz_6015 = ($signed(data_mid_2_63_imag) - $signed(data_mid_2_63_real));
  assign _zz_6016 = fixTo_571_dout;
  assign _zz_6017 = _zz_6018[35 : 0];
  assign _zz_6018 = _zz_6019;
  assign _zz_6019 = ($signed(_zz_6020) >>> _zz_479);
  assign _zz_6020 = _zz_6021;
  assign _zz_6021 = ($signed(_zz_6023) - $signed(_zz_476));
  assign _zz_6022 = ({9'd0,data_mid_2_59_real} <<< 9);
  assign _zz_6023 = {{9{_zz_6022[26]}}, _zz_6022};
  assign _zz_6024 = fixTo_572_dout;
  assign _zz_6025 = _zz_6026[35 : 0];
  assign _zz_6026 = _zz_6027;
  assign _zz_6027 = ($signed(_zz_6028) >>> _zz_479);
  assign _zz_6028 = _zz_6029;
  assign _zz_6029 = ($signed(_zz_6031) - $signed(_zz_477));
  assign _zz_6030 = ({9'd0,data_mid_2_59_imag} <<< 9);
  assign _zz_6031 = {{9{_zz_6030[26]}}, _zz_6030};
  assign _zz_6032 = fixTo_573_dout;
  assign _zz_6033 = _zz_6034[35 : 0];
  assign _zz_6034 = _zz_6035;
  assign _zz_6035 = ($signed(_zz_6036) >>> _zz_480);
  assign _zz_6036 = _zz_6037;
  assign _zz_6037 = ($signed(_zz_6039) + $signed(_zz_476));
  assign _zz_6038 = ({9'd0,data_mid_2_59_real} <<< 9);
  assign _zz_6039 = {{9{_zz_6038[26]}}, _zz_6038};
  assign _zz_6040 = fixTo_574_dout;
  assign _zz_6041 = _zz_6042[35 : 0];
  assign _zz_6042 = _zz_6043;
  assign _zz_6043 = ($signed(_zz_6044) >>> _zz_480);
  assign _zz_6044 = _zz_6045;
  assign _zz_6045 = ($signed(_zz_6047) + $signed(_zz_477));
  assign _zz_6046 = ({9'd0,data_mid_2_59_imag} <<< 9);
  assign _zz_6047 = {{9{_zz_6046[26]}}, _zz_6046};
  assign _zz_6048 = fixTo_575_dout;
  assign _zz_6049 = ($signed(twiddle_factor_table_7_real) + $signed(twiddle_factor_table_7_imag));
  assign _zz_6050 = ($signed(_zz_483) - $signed(_zz_6051));
  assign _zz_6051 = ($signed(_zz_6052) * $signed(twiddle_factor_table_7_imag));
  assign _zz_6052 = ($signed(data_mid_3_8_real) + $signed(data_mid_3_8_imag));
  assign _zz_6053 = fixTo_576_dout;
  assign _zz_6054 = ($signed(_zz_483) + $signed(_zz_6055));
  assign _zz_6055 = ($signed(_zz_6056) * $signed(twiddle_factor_table_7_real));
  assign _zz_6056 = ($signed(data_mid_3_8_imag) - $signed(data_mid_3_8_real));
  assign _zz_6057 = fixTo_577_dout;
  assign _zz_6058 = _zz_6059[35 : 0];
  assign _zz_6059 = _zz_6060;
  assign _zz_6060 = ($signed(_zz_6061) >>> _zz_484);
  assign _zz_6061 = _zz_6062;
  assign _zz_6062 = ($signed(_zz_6064) - $signed(_zz_481));
  assign _zz_6063 = ({9'd0,data_mid_3_0_real} <<< 9);
  assign _zz_6064 = {{9{_zz_6063[26]}}, _zz_6063};
  assign _zz_6065 = fixTo_578_dout;
  assign _zz_6066 = _zz_6067[35 : 0];
  assign _zz_6067 = _zz_6068;
  assign _zz_6068 = ($signed(_zz_6069) >>> _zz_484);
  assign _zz_6069 = _zz_6070;
  assign _zz_6070 = ($signed(_zz_6072) - $signed(_zz_482));
  assign _zz_6071 = ({9'd0,data_mid_3_0_imag} <<< 9);
  assign _zz_6072 = {{9{_zz_6071[26]}}, _zz_6071};
  assign _zz_6073 = fixTo_579_dout;
  assign _zz_6074 = _zz_6075[35 : 0];
  assign _zz_6075 = _zz_6076;
  assign _zz_6076 = ($signed(_zz_6077) >>> _zz_485);
  assign _zz_6077 = _zz_6078;
  assign _zz_6078 = ($signed(_zz_6080) + $signed(_zz_481));
  assign _zz_6079 = ({9'd0,data_mid_3_0_real} <<< 9);
  assign _zz_6080 = {{9{_zz_6079[26]}}, _zz_6079};
  assign _zz_6081 = fixTo_580_dout;
  assign _zz_6082 = _zz_6083[35 : 0];
  assign _zz_6083 = _zz_6084;
  assign _zz_6084 = ($signed(_zz_6085) >>> _zz_485);
  assign _zz_6085 = _zz_6086;
  assign _zz_6086 = ($signed(_zz_6088) + $signed(_zz_482));
  assign _zz_6087 = ({9'd0,data_mid_3_0_imag} <<< 9);
  assign _zz_6088 = {{9{_zz_6087[26]}}, _zz_6087};
  assign _zz_6089 = fixTo_581_dout;
  assign _zz_6090 = ($signed(twiddle_factor_table_8_real) + $signed(twiddle_factor_table_8_imag));
  assign _zz_6091 = ($signed(_zz_488) - $signed(_zz_6092));
  assign _zz_6092 = ($signed(_zz_6093) * $signed(twiddle_factor_table_8_imag));
  assign _zz_6093 = ($signed(data_mid_3_9_real) + $signed(data_mid_3_9_imag));
  assign _zz_6094 = fixTo_582_dout;
  assign _zz_6095 = ($signed(_zz_488) + $signed(_zz_6096));
  assign _zz_6096 = ($signed(_zz_6097) * $signed(twiddle_factor_table_8_real));
  assign _zz_6097 = ($signed(data_mid_3_9_imag) - $signed(data_mid_3_9_real));
  assign _zz_6098 = fixTo_583_dout;
  assign _zz_6099 = _zz_6100[35 : 0];
  assign _zz_6100 = _zz_6101;
  assign _zz_6101 = ($signed(_zz_6102) >>> _zz_489);
  assign _zz_6102 = _zz_6103;
  assign _zz_6103 = ($signed(_zz_6105) - $signed(_zz_486));
  assign _zz_6104 = ({9'd0,data_mid_3_1_real} <<< 9);
  assign _zz_6105 = {{9{_zz_6104[26]}}, _zz_6104};
  assign _zz_6106 = fixTo_584_dout;
  assign _zz_6107 = _zz_6108[35 : 0];
  assign _zz_6108 = _zz_6109;
  assign _zz_6109 = ($signed(_zz_6110) >>> _zz_489);
  assign _zz_6110 = _zz_6111;
  assign _zz_6111 = ($signed(_zz_6113) - $signed(_zz_487));
  assign _zz_6112 = ({9'd0,data_mid_3_1_imag} <<< 9);
  assign _zz_6113 = {{9{_zz_6112[26]}}, _zz_6112};
  assign _zz_6114 = fixTo_585_dout;
  assign _zz_6115 = _zz_6116[35 : 0];
  assign _zz_6116 = _zz_6117;
  assign _zz_6117 = ($signed(_zz_6118) >>> _zz_490);
  assign _zz_6118 = _zz_6119;
  assign _zz_6119 = ($signed(_zz_6121) + $signed(_zz_486));
  assign _zz_6120 = ({9'd0,data_mid_3_1_real} <<< 9);
  assign _zz_6121 = {{9{_zz_6120[26]}}, _zz_6120};
  assign _zz_6122 = fixTo_586_dout;
  assign _zz_6123 = _zz_6124[35 : 0];
  assign _zz_6124 = _zz_6125;
  assign _zz_6125 = ($signed(_zz_6126) >>> _zz_490);
  assign _zz_6126 = _zz_6127;
  assign _zz_6127 = ($signed(_zz_6129) + $signed(_zz_487));
  assign _zz_6128 = ({9'd0,data_mid_3_1_imag} <<< 9);
  assign _zz_6129 = {{9{_zz_6128[26]}}, _zz_6128};
  assign _zz_6130 = fixTo_587_dout;
  assign _zz_6131 = ($signed(twiddle_factor_table_9_real) + $signed(twiddle_factor_table_9_imag));
  assign _zz_6132 = ($signed(_zz_493) - $signed(_zz_6133));
  assign _zz_6133 = ($signed(_zz_6134) * $signed(twiddle_factor_table_9_imag));
  assign _zz_6134 = ($signed(data_mid_3_10_real) + $signed(data_mid_3_10_imag));
  assign _zz_6135 = fixTo_588_dout;
  assign _zz_6136 = ($signed(_zz_493) + $signed(_zz_6137));
  assign _zz_6137 = ($signed(_zz_6138) * $signed(twiddle_factor_table_9_real));
  assign _zz_6138 = ($signed(data_mid_3_10_imag) - $signed(data_mid_3_10_real));
  assign _zz_6139 = fixTo_589_dout;
  assign _zz_6140 = _zz_6141[35 : 0];
  assign _zz_6141 = _zz_6142;
  assign _zz_6142 = ($signed(_zz_6143) >>> _zz_494);
  assign _zz_6143 = _zz_6144;
  assign _zz_6144 = ($signed(_zz_6146) - $signed(_zz_491));
  assign _zz_6145 = ({9'd0,data_mid_3_2_real} <<< 9);
  assign _zz_6146 = {{9{_zz_6145[26]}}, _zz_6145};
  assign _zz_6147 = fixTo_590_dout;
  assign _zz_6148 = _zz_6149[35 : 0];
  assign _zz_6149 = _zz_6150;
  assign _zz_6150 = ($signed(_zz_6151) >>> _zz_494);
  assign _zz_6151 = _zz_6152;
  assign _zz_6152 = ($signed(_zz_6154) - $signed(_zz_492));
  assign _zz_6153 = ({9'd0,data_mid_3_2_imag} <<< 9);
  assign _zz_6154 = {{9{_zz_6153[26]}}, _zz_6153};
  assign _zz_6155 = fixTo_591_dout;
  assign _zz_6156 = _zz_6157[35 : 0];
  assign _zz_6157 = _zz_6158;
  assign _zz_6158 = ($signed(_zz_6159) >>> _zz_495);
  assign _zz_6159 = _zz_6160;
  assign _zz_6160 = ($signed(_zz_6162) + $signed(_zz_491));
  assign _zz_6161 = ({9'd0,data_mid_3_2_real} <<< 9);
  assign _zz_6162 = {{9{_zz_6161[26]}}, _zz_6161};
  assign _zz_6163 = fixTo_592_dout;
  assign _zz_6164 = _zz_6165[35 : 0];
  assign _zz_6165 = _zz_6166;
  assign _zz_6166 = ($signed(_zz_6167) >>> _zz_495);
  assign _zz_6167 = _zz_6168;
  assign _zz_6168 = ($signed(_zz_6170) + $signed(_zz_492));
  assign _zz_6169 = ({9'd0,data_mid_3_2_imag} <<< 9);
  assign _zz_6170 = {{9{_zz_6169[26]}}, _zz_6169};
  assign _zz_6171 = fixTo_593_dout;
  assign _zz_6172 = ($signed(twiddle_factor_table_10_real) + $signed(twiddle_factor_table_10_imag));
  assign _zz_6173 = ($signed(_zz_498) - $signed(_zz_6174));
  assign _zz_6174 = ($signed(_zz_6175) * $signed(twiddle_factor_table_10_imag));
  assign _zz_6175 = ($signed(data_mid_3_11_real) + $signed(data_mid_3_11_imag));
  assign _zz_6176 = fixTo_594_dout;
  assign _zz_6177 = ($signed(_zz_498) + $signed(_zz_6178));
  assign _zz_6178 = ($signed(_zz_6179) * $signed(twiddle_factor_table_10_real));
  assign _zz_6179 = ($signed(data_mid_3_11_imag) - $signed(data_mid_3_11_real));
  assign _zz_6180 = fixTo_595_dout;
  assign _zz_6181 = _zz_6182[35 : 0];
  assign _zz_6182 = _zz_6183;
  assign _zz_6183 = ($signed(_zz_6184) >>> _zz_499);
  assign _zz_6184 = _zz_6185;
  assign _zz_6185 = ($signed(_zz_6187) - $signed(_zz_496));
  assign _zz_6186 = ({9'd0,data_mid_3_3_real} <<< 9);
  assign _zz_6187 = {{9{_zz_6186[26]}}, _zz_6186};
  assign _zz_6188 = fixTo_596_dout;
  assign _zz_6189 = _zz_6190[35 : 0];
  assign _zz_6190 = _zz_6191;
  assign _zz_6191 = ($signed(_zz_6192) >>> _zz_499);
  assign _zz_6192 = _zz_6193;
  assign _zz_6193 = ($signed(_zz_6195) - $signed(_zz_497));
  assign _zz_6194 = ({9'd0,data_mid_3_3_imag} <<< 9);
  assign _zz_6195 = {{9{_zz_6194[26]}}, _zz_6194};
  assign _zz_6196 = fixTo_597_dout;
  assign _zz_6197 = _zz_6198[35 : 0];
  assign _zz_6198 = _zz_6199;
  assign _zz_6199 = ($signed(_zz_6200) >>> _zz_500);
  assign _zz_6200 = _zz_6201;
  assign _zz_6201 = ($signed(_zz_6203) + $signed(_zz_496));
  assign _zz_6202 = ({9'd0,data_mid_3_3_real} <<< 9);
  assign _zz_6203 = {{9{_zz_6202[26]}}, _zz_6202};
  assign _zz_6204 = fixTo_598_dout;
  assign _zz_6205 = _zz_6206[35 : 0];
  assign _zz_6206 = _zz_6207;
  assign _zz_6207 = ($signed(_zz_6208) >>> _zz_500);
  assign _zz_6208 = _zz_6209;
  assign _zz_6209 = ($signed(_zz_6211) + $signed(_zz_497));
  assign _zz_6210 = ({9'd0,data_mid_3_3_imag} <<< 9);
  assign _zz_6211 = {{9{_zz_6210[26]}}, _zz_6210};
  assign _zz_6212 = fixTo_599_dout;
  assign _zz_6213 = ($signed(twiddle_factor_table_11_real) + $signed(twiddle_factor_table_11_imag));
  assign _zz_6214 = ($signed(_zz_503) - $signed(_zz_6215));
  assign _zz_6215 = ($signed(_zz_6216) * $signed(twiddle_factor_table_11_imag));
  assign _zz_6216 = ($signed(data_mid_3_12_real) + $signed(data_mid_3_12_imag));
  assign _zz_6217 = fixTo_600_dout;
  assign _zz_6218 = ($signed(_zz_503) + $signed(_zz_6219));
  assign _zz_6219 = ($signed(_zz_6220) * $signed(twiddle_factor_table_11_real));
  assign _zz_6220 = ($signed(data_mid_3_12_imag) - $signed(data_mid_3_12_real));
  assign _zz_6221 = fixTo_601_dout;
  assign _zz_6222 = _zz_6223[35 : 0];
  assign _zz_6223 = _zz_6224;
  assign _zz_6224 = ($signed(_zz_6225) >>> _zz_504);
  assign _zz_6225 = _zz_6226;
  assign _zz_6226 = ($signed(_zz_6228) - $signed(_zz_501));
  assign _zz_6227 = ({9'd0,data_mid_3_4_real} <<< 9);
  assign _zz_6228 = {{9{_zz_6227[26]}}, _zz_6227};
  assign _zz_6229 = fixTo_602_dout;
  assign _zz_6230 = _zz_6231[35 : 0];
  assign _zz_6231 = _zz_6232;
  assign _zz_6232 = ($signed(_zz_6233) >>> _zz_504);
  assign _zz_6233 = _zz_6234;
  assign _zz_6234 = ($signed(_zz_6236) - $signed(_zz_502));
  assign _zz_6235 = ({9'd0,data_mid_3_4_imag} <<< 9);
  assign _zz_6236 = {{9{_zz_6235[26]}}, _zz_6235};
  assign _zz_6237 = fixTo_603_dout;
  assign _zz_6238 = _zz_6239[35 : 0];
  assign _zz_6239 = _zz_6240;
  assign _zz_6240 = ($signed(_zz_6241) >>> _zz_505);
  assign _zz_6241 = _zz_6242;
  assign _zz_6242 = ($signed(_zz_6244) + $signed(_zz_501));
  assign _zz_6243 = ({9'd0,data_mid_3_4_real} <<< 9);
  assign _zz_6244 = {{9{_zz_6243[26]}}, _zz_6243};
  assign _zz_6245 = fixTo_604_dout;
  assign _zz_6246 = _zz_6247[35 : 0];
  assign _zz_6247 = _zz_6248;
  assign _zz_6248 = ($signed(_zz_6249) >>> _zz_505);
  assign _zz_6249 = _zz_6250;
  assign _zz_6250 = ($signed(_zz_6252) + $signed(_zz_502));
  assign _zz_6251 = ({9'd0,data_mid_3_4_imag} <<< 9);
  assign _zz_6252 = {{9{_zz_6251[26]}}, _zz_6251};
  assign _zz_6253 = fixTo_605_dout;
  assign _zz_6254 = ($signed(twiddle_factor_table_12_real) + $signed(twiddle_factor_table_12_imag));
  assign _zz_6255 = ($signed(_zz_508) - $signed(_zz_6256));
  assign _zz_6256 = ($signed(_zz_6257) * $signed(twiddle_factor_table_12_imag));
  assign _zz_6257 = ($signed(data_mid_3_13_real) + $signed(data_mid_3_13_imag));
  assign _zz_6258 = fixTo_606_dout;
  assign _zz_6259 = ($signed(_zz_508) + $signed(_zz_6260));
  assign _zz_6260 = ($signed(_zz_6261) * $signed(twiddle_factor_table_12_real));
  assign _zz_6261 = ($signed(data_mid_3_13_imag) - $signed(data_mid_3_13_real));
  assign _zz_6262 = fixTo_607_dout;
  assign _zz_6263 = _zz_6264[35 : 0];
  assign _zz_6264 = _zz_6265;
  assign _zz_6265 = ($signed(_zz_6266) >>> _zz_509);
  assign _zz_6266 = _zz_6267;
  assign _zz_6267 = ($signed(_zz_6269) - $signed(_zz_506));
  assign _zz_6268 = ({9'd0,data_mid_3_5_real} <<< 9);
  assign _zz_6269 = {{9{_zz_6268[26]}}, _zz_6268};
  assign _zz_6270 = fixTo_608_dout;
  assign _zz_6271 = _zz_6272[35 : 0];
  assign _zz_6272 = _zz_6273;
  assign _zz_6273 = ($signed(_zz_6274) >>> _zz_509);
  assign _zz_6274 = _zz_6275;
  assign _zz_6275 = ($signed(_zz_6277) - $signed(_zz_507));
  assign _zz_6276 = ({9'd0,data_mid_3_5_imag} <<< 9);
  assign _zz_6277 = {{9{_zz_6276[26]}}, _zz_6276};
  assign _zz_6278 = fixTo_609_dout;
  assign _zz_6279 = _zz_6280[35 : 0];
  assign _zz_6280 = _zz_6281;
  assign _zz_6281 = ($signed(_zz_6282) >>> _zz_510);
  assign _zz_6282 = _zz_6283;
  assign _zz_6283 = ($signed(_zz_6285) + $signed(_zz_506));
  assign _zz_6284 = ({9'd0,data_mid_3_5_real} <<< 9);
  assign _zz_6285 = {{9{_zz_6284[26]}}, _zz_6284};
  assign _zz_6286 = fixTo_610_dout;
  assign _zz_6287 = _zz_6288[35 : 0];
  assign _zz_6288 = _zz_6289;
  assign _zz_6289 = ($signed(_zz_6290) >>> _zz_510);
  assign _zz_6290 = _zz_6291;
  assign _zz_6291 = ($signed(_zz_6293) + $signed(_zz_507));
  assign _zz_6292 = ({9'd0,data_mid_3_5_imag} <<< 9);
  assign _zz_6293 = {{9{_zz_6292[26]}}, _zz_6292};
  assign _zz_6294 = fixTo_611_dout;
  assign _zz_6295 = ($signed(twiddle_factor_table_13_real) + $signed(twiddle_factor_table_13_imag));
  assign _zz_6296 = ($signed(_zz_513) - $signed(_zz_6297));
  assign _zz_6297 = ($signed(_zz_6298) * $signed(twiddle_factor_table_13_imag));
  assign _zz_6298 = ($signed(data_mid_3_14_real) + $signed(data_mid_3_14_imag));
  assign _zz_6299 = fixTo_612_dout;
  assign _zz_6300 = ($signed(_zz_513) + $signed(_zz_6301));
  assign _zz_6301 = ($signed(_zz_6302) * $signed(twiddle_factor_table_13_real));
  assign _zz_6302 = ($signed(data_mid_3_14_imag) - $signed(data_mid_3_14_real));
  assign _zz_6303 = fixTo_613_dout;
  assign _zz_6304 = _zz_6305[35 : 0];
  assign _zz_6305 = _zz_6306;
  assign _zz_6306 = ($signed(_zz_6307) >>> _zz_514);
  assign _zz_6307 = _zz_6308;
  assign _zz_6308 = ($signed(_zz_6310) - $signed(_zz_511));
  assign _zz_6309 = ({9'd0,data_mid_3_6_real} <<< 9);
  assign _zz_6310 = {{9{_zz_6309[26]}}, _zz_6309};
  assign _zz_6311 = fixTo_614_dout;
  assign _zz_6312 = _zz_6313[35 : 0];
  assign _zz_6313 = _zz_6314;
  assign _zz_6314 = ($signed(_zz_6315) >>> _zz_514);
  assign _zz_6315 = _zz_6316;
  assign _zz_6316 = ($signed(_zz_6318) - $signed(_zz_512));
  assign _zz_6317 = ({9'd0,data_mid_3_6_imag} <<< 9);
  assign _zz_6318 = {{9{_zz_6317[26]}}, _zz_6317};
  assign _zz_6319 = fixTo_615_dout;
  assign _zz_6320 = _zz_6321[35 : 0];
  assign _zz_6321 = _zz_6322;
  assign _zz_6322 = ($signed(_zz_6323) >>> _zz_515);
  assign _zz_6323 = _zz_6324;
  assign _zz_6324 = ($signed(_zz_6326) + $signed(_zz_511));
  assign _zz_6325 = ({9'd0,data_mid_3_6_real} <<< 9);
  assign _zz_6326 = {{9{_zz_6325[26]}}, _zz_6325};
  assign _zz_6327 = fixTo_616_dout;
  assign _zz_6328 = _zz_6329[35 : 0];
  assign _zz_6329 = _zz_6330;
  assign _zz_6330 = ($signed(_zz_6331) >>> _zz_515);
  assign _zz_6331 = _zz_6332;
  assign _zz_6332 = ($signed(_zz_6334) + $signed(_zz_512));
  assign _zz_6333 = ({9'd0,data_mid_3_6_imag} <<< 9);
  assign _zz_6334 = {{9{_zz_6333[26]}}, _zz_6333};
  assign _zz_6335 = fixTo_617_dout;
  assign _zz_6336 = ($signed(twiddle_factor_table_14_real) + $signed(twiddle_factor_table_14_imag));
  assign _zz_6337 = ($signed(_zz_518) - $signed(_zz_6338));
  assign _zz_6338 = ($signed(_zz_6339) * $signed(twiddle_factor_table_14_imag));
  assign _zz_6339 = ($signed(data_mid_3_15_real) + $signed(data_mid_3_15_imag));
  assign _zz_6340 = fixTo_618_dout;
  assign _zz_6341 = ($signed(_zz_518) + $signed(_zz_6342));
  assign _zz_6342 = ($signed(_zz_6343) * $signed(twiddle_factor_table_14_real));
  assign _zz_6343 = ($signed(data_mid_3_15_imag) - $signed(data_mid_3_15_real));
  assign _zz_6344 = fixTo_619_dout;
  assign _zz_6345 = _zz_6346[35 : 0];
  assign _zz_6346 = _zz_6347;
  assign _zz_6347 = ($signed(_zz_6348) >>> _zz_519);
  assign _zz_6348 = _zz_6349;
  assign _zz_6349 = ($signed(_zz_6351) - $signed(_zz_516));
  assign _zz_6350 = ({9'd0,data_mid_3_7_real} <<< 9);
  assign _zz_6351 = {{9{_zz_6350[26]}}, _zz_6350};
  assign _zz_6352 = fixTo_620_dout;
  assign _zz_6353 = _zz_6354[35 : 0];
  assign _zz_6354 = _zz_6355;
  assign _zz_6355 = ($signed(_zz_6356) >>> _zz_519);
  assign _zz_6356 = _zz_6357;
  assign _zz_6357 = ($signed(_zz_6359) - $signed(_zz_517));
  assign _zz_6358 = ({9'd0,data_mid_3_7_imag} <<< 9);
  assign _zz_6359 = {{9{_zz_6358[26]}}, _zz_6358};
  assign _zz_6360 = fixTo_621_dout;
  assign _zz_6361 = _zz_6362[35 : 0];
  assign _zz_6362 = _zz_6363;
  assign _zz_6363 = ($signed(_zz_6364) >>> _zz_520);
  assign _zz_6364 = _zz_6365;
  assign _zz_6365 = ($signed(_zz_6367) + $signed(_zz_516));
  assign _zz_6366 = ({9'd0,data_mid_3_7_real} <<< 9);
  assign _zz_6367 = {{9{_zz_6366[26]}}, _zz_6366};
  assign _zz_6368 = fixTo_622_dout;
  assign _zz_6369 = _zz_6370[35 : 0];
  assign _zz_6370 = _zz_6371;
  assign _zz_6371 = ($signed(_zz_6372) >>> _zz_520);
  assign _zz_6372 = _zz_6373;
  assign _zz_6373 = ($signed(_zz_6375) + $signed(_zz_517));
  assign _zz_6374 = ({9'd0,data_mid_3_7_imag} <<< 9);
  assign _zz_6375 = {{9{_zz_6374[26]}}, _zz_6374};
  assign _zz_6376 = fixTo_623_dout;
  assign _zz_6377 = ($signed(twiddle_factor_table_7_real) + $signed(twiddle_factor_table_7_imag));
  assign _zz_6378 = ($signed(_zz_523) - $signed(_zz_6379));
  assign _zz_6379 = ($signed(_zz_6380) * $signed(twiddle_factor_table_7_imag));
  assign _zz_6380 = ($signed(data_mid_3_24_real) + $signed(data_mid_3_24_imag));
  assign _zz_6381 = fixTo_624_dout;
  assign _zz_6382 = ($signed(_zz_523) + $signed(_zz_6383));
  assign _zz_6383 = ($signed(_zz_6384) * $signed(twiddle_factor_table_7_real));
  assign _zz_6384 = ($signed(data_mid_3_24_imag) - $signed(data_mid_3_24_real));
  assign _zz_6385 = fixTo_625_dout;
  assign _zz_6386 = _zz_6387[35 : 0];
  assign _zz_6387 = _zz_6388;
  assign _zz_6388 = ($signed(_zz_6389) >>> _zz_524);
  assign _zz_6389 = _zz_6390;
  assign _zz_6390 = ($signed(_zz_6392) - $signed(_zz_521));
  assign _zz_6391 = ({9'd0,data_mid_3_16_real} <<< 9);
  assign _zz_6392 = {{9{_zz_6391[26]}}, _zz_6391};
  assign _zz_6393 = fixTo_626_dout;
  assign _zz_6394 = _zz_6395[35 : 0];
  assign _zz_6395 = _zz_6396;
  assign _zz_6396 = ($signed(_zz_6397) >>> _zz_524);
  assign _zz_6397 = _zz_6398;
  assign _zz_6398 = ($signed(_zz_6400) - $signed(_zz_522));
  assign _zz_6399 = ({9'd0,data_mid_3_16_imag} <<< 9);
  assign _zz_6400 = {{9{_zz_6399[26]}}, _zz_6399};
  assign _zz_6401 = fixTo_627_dout;
  assign _zz_6402 = _zz_6403[35 : 0];
  assign _zz_6403 = _zz_6404;
  assign _zz_6404 = ($signed(_zz_6405) >>> _zz_525);
  assign _zz_6405 = _zz_6406;
  assign _zz_6406 = ($signed(_zz_6408) + $signed(_zz_521));
  assign _zz_6407 = ({9'd0,data_mid_3_16_real} <<< 9);
  assign _zz_6408 = {{9{_zz_6407[26]}}, _zz_6407};
  assign _zz_6409 = fixTo_628_dout;
  assign _zz_6410 = _zz_6411[35 : 0];
  assign _zz_6411 = _zz_6412;
  assign _zz_6412 = ($signed(_zz_6413) >>> _zz_525);
  assign _zz_6413 = _zz_6414;
  assign _zz_6414 = ($signed(_zz_6416) + $signed(_zz_522));
  assign _zz_6415 = ({9'd0,data_mid_3_16_imag} <<< 9);
  assign _zz_6416 = {{9{_zz_6415[26]}}, _zz_6415};
  assign _zz_6417 = fixTo_629_dout;
  assign _zz_6418 = ($signed(twiddle_factor_table_8_real) + $signed(twiddle_factor_table_8_imag));
  assign _zz_6419 = ($signed(_zz_528) - $signed(_zz_6420));
  assign _zz_6420 = ($signed(_zz_6421) * $signed(twiddle_factor_table_8_imag));
  assign _zz_6421 = ($signed(data_mid_3_25_real) + $signed(data_mid_3_25_imag));
  assign _zz_6422 = fixTo_630_dout;
  assign _zz_6423 = ($signed(_zz_528) + $signed(_zz_6424));
  assign _zz_6424 = ($signed(_zz_6425) * $signed(twiddle_factor_table_8_real));
  assign _zz_6425 = ($signed(data_mid_3_25_imag) - $signed(data_mid_3_25_real));
  assign _zz_6426 = fixTo_631_dout;
  assign _zz_6427 = _zz_6428[35 : 0];
  assign _zz_6428 = _zz_6429;
  assign _zz_6429 = ($signed(_zz_6430) >>> _zz_529);
  assign _zz_6430 = _zz_6431;
  assign _zz_6431 = ($signed(_zz_6433) - $signed(_zz_526));
  assign _zz_6432 = ({9'd0,data_mid_3_17_real} <<< 9);
  assign _zz_6433 = {{9{_zz_6432[26]}}, _zz_6432};
  assign _zz_6434 = fixTo_632_dout;
  assign _zz_6435 = _zz_6436[35 : 0];
  assign _zz_6436 = _zz_6437;
  assign _zz_6437 = ($signed(_zz_6438) >>> _zz_529);
  assign _zz_6438 = _zz_6439;
  assign _zz_6439 = ($signed(_zz_6441) - $signed(_zz_527));
  assign _zz_6440 = ({9'd0,data_mid_3_17_imag} <<< 9);
  assign _zz_6441 = {{9{_zz_6440[26]}}, _zz_6440};
  assign _zz_6442 = fixTo_633_dout;
  assign _zz_6443 = _zz_6444[35 : 0];
  assign _zz_6444 = _zz_6445;
  assign _zz_6445 = ($signed(_zz_6446) >>> _zz_530);
  assign _zz_6446 = _zz_6447;
  assign _zz_6447 = ($signed(_zz_6449) + $signed(_zz_526));
  assign _zz_6448 = ({9'd0,data_mid_3_17_real} <<< 9);
  assign _zz_6449 = {{9{_zz_6448[26]}}, _zz_6448};
  assign _zz_6450 = fixTo_634_dout;
  assign _zz_6451 = _zz_6452[35 : 0];
  assign _zz_6452 = _zz_6453;
  assign _zz_6453 = ($signed(_zz_6454) >>> _zz_530);
  assign _zz_6454 = _zz_6455;
  assign _zz_6455 = ($signed(_zz_6457) + $signed(_zz_527));
  assign _zz_6456 = ({9'd0,data_mid_3_17_imag} <<< 9);
  assign _zz_6457 = {{9{_zz_6456[26]}}, _zz_6456};
  assign _zz_6458 = fixTo_635_dout;
  assign _zz_6459 = ($signed(twiddle_factor_table_9_real) + $signed(twiddle_factor_table_9_imag));
  assign _zz_6460 = ($signed(_zz_533) - $signed(_zz_6461));
  assign _zz_6461 = ($signed(_zz_6462) * $signed(twiddle_factor_table_9_imag));
  assign _zz_6462 = ($signed(data_mid_3_26_real) + $signed(data_mid_3_26_imag));
  assign _zz_6463 = fixTo_636_dout;
  assign _zz_6464 = ($signed(_zz_533) + $signed(_zz_6465));
  assign _zz_6465 = ($signed(_zz_6466) * $signed(twiddle_factor_table_9_real));
  assign _zz_6466 = ($signed(data_mid_3_26_imag) - $signed(data_mid_3_26_real));
  assign _zz_6467 = fixTo_637_dout;
  assign _zz_6468 = _zz_6469[35 : 0];
  assign _zz_6469 = _zz_6470;
  assign _zz_6470 = ($signed(_zz_6471) >>> _zz_534);
  assign _zz_6471 = _zz_6472;
  assign _zz_6472 = ($signed(_zz_6474) - $signed(_zz_531));
  assign _zz_6473 = ({9'd0,data_mid_3_18_real} <<< 9);
  assign _zz_6474 = {{9{_zz_6473[26]}}, _zz_6473};
  assign _zz_6475 = fixTo_638_dout;
  assign _zz_6476 = _zz_6477[35 : 0];
  assign _zz_6477 = _zz_6478;
  assign _zz_6478 = ($signed(_zz_6479) >>> _zz_534);
  assign _zz_6479 = _zz_6480;
  assign _zz_6480 = ($signed(_zz_6482) - $signed(_zz_532));
  assign _zz_6481 = ({9'd0,data_mid_3_18_imag} <<< 9);
  assign _zz_6482 = {{9{_zz_6481[26]}}, _zz_6481};
  assign _zz_6483 = fixTo_639_dout;
  assign _zz_6484 = _zz_6485[35 : 0];
  assign _zz_6485 = _zz_6486;
  assign _zz_6486 = ($signed(_zz_6487) >>> _zz_535);
  assign _zz_6487 = _zz_6488;
  assign _zz_6488 = ($signed(_zz_6490) + $signed(_zz_531));
  assign _zz_6489 = ({9'd0,data_mid_3_18_real} <<< 9);
  assign _zz_6490 = {{9{_zz_6489[26]}}, _zz_6489};
  assign _zz_6491 = fixTo_640_dout;
  assign _zz_6492 = _zz_6493[35 : 0];
  assign _zz_6493 = _zz_6494;
  assign _zz_6494 = ($signed(_zz_6495) >>> _zz_535);
  assign _zz_6495 = _zz_6496;
  assign _zz_6496 = ($signed(_zz_6498) + $signed(_zz_532));
  assign _zz_6497 = ({9'd0,data_mid_3_18_imag} <<< 9);
  assign _zz_6498 = {{9{_zz_6497[26]}}, _zz_6497};
  assign _zz_6499 = fixTo_641_dout;
  assign _zz_6500 = ($signed(twiddle_factor_table_10_real) + $signed(twiddle_factor_table_10_imag));
  assign _zz_6501 = ($signed(_zz_538) - $signed(_zz_6502));
  assign _zz_6502 = ($signed(_zz_6503) * $signed(twiddle_factor_table_10_imag));
  assign _zz_6503 = ($signed(data_mid_3_27_real) + $signed(data_mid_3_27_imag));
  assign _zz_6504 = fixTo_642_dout;
  assign _zz_6505 = ($signed(_zz_538) + $signed(_zz_6506));
  assign _zz_6506 = ($signed(_zz_6507) * $signed(twiddle_factor_table_10_real));
  assign _zz_6507 = ($signed(data_mid_3_27_imag) - $signed(data_mid_3_27_real));
  assign _zz_6508 = fixTo_643_dout;
  assign _zz_6509 = _zz_6510[35 : 0];
  assign _zz_6510 = _zz_6511;
  assign _zz_6511 = ($signed(_zz_6512) >>> _zz_539);
  assign _zz_6512 = _zz_6513;
  assign _zz_6513 = ($signed(_zz_6515) - $signed(_zz_536));
  assign _zz_6514 = ({9'd0,data_mid_3_19_real} <<< 9);
  assign _zz_6515 = {{9{_zz_6514[26]}}, _zz_6514};
  assign _zz_6516 = fixTo_644_dout;
  assign _zz_6517 = _zz_6518[35 : 0];
  assign _zz_6518 = _zz_6519;
  assign _zz_6519 = ($signed(_zz_6520) >>> _zz_539);
  assign _zz_6520 = _zz_6521;
  assign _zz_6521 = ($signed(_zz_6523) - $signed(_zz_537));
  assign _zz_6522 = ({9'd0,data_mid_3_19_imag} <<< 9);
  assign _zz_6523 = {{9{_zz_6522[26]}}, _zz_6522};
  assign _zz_6524 = fixTo_645_dout;
  assign _zz_6525 = _zz_6526[35 : 0];
  assign _zz_6526 = _zz_6527;
  assign _zz_6527 = ($signed(_zz_6528) >>> _zz_540);
  assign _zz_6528 = _zz_6529;
  assign _zz_6529 = ($signed(_zz_6531) + $signed(_zz_536));
  assign _zz_6530 = ({9'd0,data_mid_3_19_real} <<< 9);
  assign _zz_6531 = {{9{_zz_6530[26]}}, _zz_6530};
  assign _zz_6532 = fixTo_646_dout;
  assign _zz_6533 = _zz_6534[35 : 0];
  assign _zz_6534 = _zz_6535;
  assign _zz_6535 = ($signed(_zz_6536) >>> _zz_540);
  assign _zz_6536 = _zz_6537;
  assign _zz_6537 = ($signed(_zz_6539) + $signed(_zz_537));
  assign _zz_6538 = ({9'd0,data_mid_3_19_imag} <<< 9);
  assign _zz_6539 = {{9{_zz_6538[26]}}, _zz_6538};
  assign _zz_6540 = fixTo_647_dout;
  assign _zz_6541 = ($signed(twiddle_factor_table_11_real) + $signed(twiddle_factor_table_11_imag));
  assign _zz_6542 = ($signed(_zz_543) - $signed(_zz_6543));
  assign _zz_6543 = ($signed(_zz_6544) * $signed(twiddle_factor_table_11_imag));
  assign _zz_6544 = ($signed(data_mid_3_28_real) + $signed(data_mid_3_28_imag));
  assign _zz_6545 = fixTo_648_dout;
  assign _zz_6546 = ($signed(_zz_543) + $signed(_zz_6547));
  assign _zz_6547 = ($signed(_zz_6548) * $signed(twiddle_factor_table_11_real));
  assign _zz_6548 = ($signed(data_mid_3_28_imag) - $signed(data_mid_3_28_real));
  assign _zz_6549 = fixTo_649_dout;
  assign _zz_6550 = _zz_6551[35 : 0];
  assign _zz_6551 = _zz_6552;
  assign _zz_6552 = ($signed(_zz_6553) >>> _zz_544);
  assign _zz_6553 = _zz_6554;
  assign _zz_6554 = ($signed(_zz_6556) - $signed(_zz_541));
  assign _zz_6555 = ({9'd0,data_mid_3_20_real} <<< 9);
  assign _zz_6556 = {{9{_zz_6555[26]}}, _zz_6555};
  assign _zz_6557 = fixTo_650_dout;
  assign _zz_6558 = _zz_6559[35 : 0];
  assign _zz_6559 = _zz_6560;
  assign _zz_6560 = ($signed(_zz_6561) >>> _zz_544);
  assign _zz_6561 = _zz_6562;
  assign _zz_6562 = ($signed(_zz_6564) - $signed(_zz_542));
  assign _zz_6563 = ({9'd0,data_mid_3_20_imag} <<< 9);
  assign _zz_6564 = {{9{_zz_6563[26]}}, _zz_6563};
  assign _zz_6565 = fixTo_651_dout;
  assign _zz_6566 = _zz_6567[35 : 0];
  assign _zz_6567 = _zz_6568;
  assign _zz_6568 = ($signed(_zz_6569) >>> _zz_545);
  assign _zz_6569 = _zz_6570;
  assign _zz_6570 = ($signed(_zz_6572) + $signed(_zz_541));
  assign _zz_6571 = ({9'd0,data_mid_3_20_real} <<< 9);
  assign _zz_6572 = {{9{_zz_6571[26]}}, _zz_6571};
  assign _zz_6573 = fixTo_652_dout;
  assign _zz_6574 = _zz_6575[35 : 0];
  assign _zz_6575 = _zz_6576;
  assign _zz_6576 = ($signed(_zz_6577) >>> _zz_545);
  assign _zz_6577 = _zz_6578;
  assign _zz_6578 = ($signed(_zz_6580) + $signed(_zz_542));
  assign _zz_6579 = ({9'd0,data_mid_3_20_imag} <<< 9);
  assign _zz_6580 = {{9{_zz_6579[26]}}, _zz_6579};
  assign _zz_6581 = fixTo_653_dout;
  assign _zz_6582 = ($signed(twiddle_factor_table_12_real) + $signed(twiddle_factor_table_12_imag));
  assign _zz_6583 = ($signed(_zz_548) - $signed(_zz_6584));
  assign _zz_6584 = ($signed(_zz_6585) * $signed(twiddle_factor_table_12_imag));
  assign _zz_6585 = ($signed(data_mid_3_29_real) + $signed(data_mid_3_29_imag));
  assign _zz_6586 = fixTo_654_dout;
  assign _zz_6587 = ($signed(_zz_548) + $signed(_zz_6588));
  assign _zz_6588 = ($signed(_zz_6589) * $signed(twiddle_factor_table_12_real));
  assign _zz_6589 = ($signed(data_mid_3_29_imag) - $signed(data_mid_3_29_real));
  assign _zz_6590 = fixTo_655_dout;
  assign _zz_6591 = _zz_6592[35 : 0];
  assign _zz_6592 = _zz_6593;
  assign _zz_6593 = ($signed(_zz_6594) >>> _zz_549);
  assign _zz_6594 = _zz_6595;
  assign _zz_6595 = ($signed(_zz_6597) - $signed(_zz_546));
  assign _zz_6596 = ({9'd0,data_mid_3_21_real} <<< 9);
  assign _zz_6597 = {{9{_zz_6596[26]}}, _zz_6596};
  assign _zz_6598 = fixTo_656_dout;
  assign _zz_6599 = _zz_6600[35 : 0];
  assign _zz_6600 = _zz_6601;
  assign _zz_6601 = ($signed(_zz_6602) >>> _zz_549);
  assign _zz_6602 = _zz_6603;
  assign _zz_6603 = ($signed(_zz_6605) - $signed(_zz_547));
  assign _zz_6604 = ({9'd0,data_mid_3_21_imag} <<< 9);
  assign _zz_6605 = {{9{_zz_6604[26]}}, _zz_6604};
  assign _zz_6606 = fixTo_657_dout;
  assign _zz_6607 = _zz_6608[35 : 0];
  assign _zz_6608 = _zz_6609;
  assign _zz_6609 = ($signed(_zz_6610) >>> _zz_550);
  assign _zz_6610 = _zz_6611;
  assign _zz_6611 = ($signed(_zz_6613) + $signed(_zz_546));
  assign _zz_6612 = ({9'd0,data_mid_3_21_real} <<< 9);
  assign _zz_6613 = {{9{_zz_6612[26]}}, _zz_6612};
  assign _zz_6614 = fixTo_658_dout;
  assign _zz_6615 = _zz_6616[35 : 0];
  assign _zz_6616 = _zz_6617;
  assign _zz_6617 = ($signed(_zz_6618) >>> _zz_550);
  assign _zz_6618 = _zz_6619;
  assign _zz_6619 = ($signed(_zz_6621) + $signed(_zz_547));
  assign _zz_6620 = ({9'd0,data_mid_3_21_imag} <<< 9);
  assign _zz_6621 = {{9{_zz_6620[26]}}, _zz_6620};
  assign _zz_6622 = fixTo_659_dout;
  assign _zz_6623 = ($signed(twiddle_factor_table_13_real) + $signed(twiddle_factor_table_13_imag));
  assign _zz_6624 = ($signed(_zz_553) - $signed(_zz_6625));
  assign _zz_6625 = ($signed(_zz_6626) * $signed(twiddle_factor_table_13_imag));
  assign _zz_6626 = ($signed(data_mid_3_30_real) + $signed(data_mid_3_30_imag));
  assign _zz_6627 = fixTo_660_dout;
  assign _zz_6628 = ($signed(_zz_553) + $signed(_zz_6629));
  assign _zz_6629 = ($signed(_zz_6630) * $signed(twiddle_factor_table_13_real));
  assign _zz_6630 = ($signed(data_mid_3_30_imag) - $signed(data_mid_3_30_real));
  assign _zz_6631 = fixTo_661_dout;
  assign _zz_6632 = _zz_6633[35 : 0];
  assign _zz_6633 = _zz_6634;
  assign _zz_6634 = ($signed(_zz_6635) >>> _zz_554);
  assign _zz_6635 = _zz_6636;
  assign _zz_6636 = ($signed(_zz_6638) - $signed(_zz_551));
  assign _zz_6637 = ({9'd0,data_mid_3_22_real} <<< 9);
  assign _zz_6638 = {{9{_zz_6637[26]}}, _zz_6637};
  assign _zz_6639 = fixTo_662_dout;
  assign _zz_6640 = _zz_6641[35 : 0];
  assign _zz_6641 = _zz_6642;
  assign _zz_6642 = ($signed(_zz_6643) >>> _zz_554);
  assign _zz_6643 = _zz_6644;
  assign _zz_6644 = ($signed(_zz_6646) - $signed(_zz_552));
  assign _zz_6645 = ({9'd0,data_mid_3_22_imag} <<< 9);
  assign _zz_6646 = {{9{_zz_6645[26]}}, _zz_6645};
  assign _zz_6647 = fixTo_663_dout;
  assign _zz_6648 = _zz_6649[35 : 0];
  assign _zz_6649 = _zz_6650;
  assign _zz_6650 = ($signed(_zz_6651) >>> _zz_555);
  assign _zz_6651 = _zz_6652;
  assign _zz_6652 = ($signed(_zz_6654) + $signed(_zz_551));
  assign _zz_6653 = ({9'd0,data_mid_3_22_real} <<< 9);
  assign _zz_6654 = {{9{_zz_6653[26]}}, _zz_6653};
  assign _zz_6655 = fixTo_664_dout;
  assign _zz_6656 = _zz_6657[35 : 0];
  assign _zz_6657 = _zz_6658;
  assign _zz_6658 = ($signed(_zz_6659) >>> _zz_555);
  assign _zz_6659 = _zz_6660;
  assign _zz_6660 = ($signed(_zz_6662) + $signed(_zz_552));
  assign _zz_6661 = ({9'd0,data_mid_3_22_imag} <<< 9);
  assign _zz_6662 = {{9{_zz_6661[26]}}, _zz_6661};
  assign _zz_6663 = fixTo_665_dout;
  assign _zz_6664 = ($signed(twiddle_factor_table_14_real) + $signed(twiddle_factor_table_14_imag));
  assign _zz_6665 = ($signed(_zz_558) - $signed(_zz_6666));
  assign _zz_6666 = ($signed(_zz_6667) * $signed(twiddle_factor_table_14_imag));
  assign _zz_6667 = ($signed(data_mid_3_31_real) + $signed(data_mid_3_31_imag));
  assign _zz_6668 = fixTo_666_dout;
  assign _zz_6669 = ($signed(_zz_558) + $signed(_zz_6670));
  assign _zz_6670 = ($signed(_zz_6671) * $signed(twiddle_factor_table_14_real));
  assign _zz_6671 = ($signed(data_mid_3_31_imag) - $signed(data_mid_3_31_real));
  assign _zz_6672 = fixTo_667_dout;
  assign _zz_6673 = _zz_6674[35 : 0];
  assign _zz_6674 = _zz_6675;
  assign _zz_6675 = ($signed(_zz_6676) >>> _zz_559);
  assign _zz_6676 = _zz_6677;
  assign _zz_6677 = ($signed(_zz_6679) - $signed(_zz_556));
  assign _zz_6678 = ({9'd0,data_mid_3_23_real} <<< 9);
  assign _zz_6679 = {{9{_zz_6678[26]}}, _zz_6678};
  assign _zz_6680 = fixTo_668_dout;
  assign _zz_6681 = _zz_6682[35 : 0];
  assign _zz_6682 = _zz_6683;
  assign _zz_6683 = ($signed(_zz_6684) >>> _zz_559);
  assign _zz_6684 = _zz_6685;
  assign _zz_6685 = ($signed(_zz_6687) - $signed(_zz_557));
  assign _zz_6686 = ({9'd0,data_mid_3_23_imag} <<< 9);
  assign _zz_6687 = {{9{_zz_6686[26]}}, _zz_6686};
  assign _zz_6688 = fixTo_669_dout;
  assign _zz_6689 = _zz_6690[35 : 0];
  assign _zz_6690 = _zz_6691;
  assign _zz_6691 = ($signed(_zz_6692) >>> _zz_560);
  assign _zz_6692 = _zz_6693;
  assign _zz_6693 = ($signed(_zz_6695) + $signed(_zz_556));
  assign _zz_6694 = ({9'd0,data_mid_3_23_real} <<< 9);
  assign _zz_6695 = {{9{_zz_6694[26]}}, _zz_6694};
  assign _zz_6696 = fixTo_670_dout;
  assign _zz_6697 = _zz_6698[35 : 0];
  assign _zz_6698 = _zz_6699;
  assign _zz_6699 = ($signed(_zz_6700) >>> _zz_560);
  assign _zz_6700 = _zz_6701;
  assign _zz_6701 = ($signed(_zz_6703) + $signed(_zz_557));
  assign _zz_6702 = ({9'd0,data_mid_3_23_imag} <<< 9);
  assign _zz_6703 = {{9{_zz_6702[26]}}, _zz_6702};
  assign _zz_6704 = fixTo_671_dout;
  assign _zz_6705 = ($signed(twiddle_factor_table_7_real) + $signed(twiddle_factor_table_7_imag));
  assign _zz_6706 = ($signed(_zz_563) - $signed(_zz_6707));
  assign _zz_6707 = ($signed(_zz_6708) * $signed(twiddle_factor_table_7_imag));
  assign _zz_6708 = ($signed(data_mid_3_40_real) + $signed(data_mid_3_40_imag));
  assign _zz_6709 = fixTo_672_dout;
  assign _zz_6710 = ($signed(_zz_563) + $signed(_zz_6711));
  assign _zz_6711 = ($signed(_zz_6712) * $signed(twiddle_factor_table_7_real));
  assign _zz_6712 = ($signed(data_mid_3_40_imag) - $signed(data_mid_3_40_real));
  assign _zz_6713 = fixTo_673_dout;
  assign _zz_6714 = _zz_6715[35 : 0];
  assign _zz_6715 = _zz_6716;
  assign _zz_6716 = ($signed(_zz_6717) >>> _zz_564);
  assign _zz_6717 = _zz_6718;
  assign _zz_6718 = ($signed(_zz_6720) - $signed(_zz_561));
  assign _zz_6719 = ({9'd0,data_mid_3_32_real} <<< 9);
  assign _zz_6720 = {{9{_zz_6719[26]}}, _zz_6719};
  assign _zz_6721 = fixTo_674_dout;
  assign _zz_6722 = _zz_6723[35 : 0];
  assign _zz_6723 = _zz_6724;
  assign _zz_6724 = ($signed(_zz_6725) >>> _zz_564);
  assign _zz_6725 = _zz_6726;
  assign _zz_6726 = ($signed(_zz_6728) - $signed(_zz_562));
  assign _zz_6727 = ({9'd0,data_mid_3_32_imag} <<< 9);
  assign _zz_6728 = {{9{_zz_6727[26]}}, _zz_6727};
  assign _zz_6729 = fixTo_675_dout;
  assign _zz_6730 = _zz_6731[35 : 0];
  assign _zz_6731 = _zz_6732;
  assign _zz_6732 = ($signed(_zz_6733) >>> _zz_565);
  assign _zz_6733 = _zz_6734;
  assign _zz_6734 = ($signed(_zz_6736) + $signed(_zz_561));
  assign _zz_6735 = ({9'd0,data_mid_3_32_real} <<< 9);
  assign _zz_6736 = {{9{_zz_6735[26]}}, _zz_6735};
  assign _zz_6737 = fixTo_676_dout;
  assign _zz_6738 = _zz_6739[35 : 0];
  assign _zz_6739 = _zz_6740;
  assign _zz_6740 = ($signed(_zz_6741) >>> _zz_565);
  assign _zz_6741 = _zz_6742;
  assign _zz_6742 = ($signed(_zz_6744) + $signed(_zz_562));
  assign _zz_6743 = ({9'd0,data_mid_3_32_imag} <<< 9);
  assign _zz_6744 = {{9{_zz_6743[26]}}, _zz_6743};
  assign _zz_6745 = fixTo_677_dout;
  assign _zz_6746 = ($signed(twiddle_factor_table_8_real) + $signed(twiddle_factor_table_8_imag));
  assign _zz_6747 = ($signed(_zz_568) - $signed(_zz_6748));
  assign _zz_6748 = ($signed(_zz_6749) * $signed(twiddle_factor_table_8_imag));
  assign _zz_6749 = ($signed(data_mid_3_41_real) + $signed(data_mid_3_41_imag));
  assign _zz_6750 = fixTo_678_dout;
  assign _zz_6751 = ($signed(_zz_568) + $signed(_zz_6752));
  assign _zz_6752 = ($signed(_zz_6753) * $signed(twiddle_factor_table_8_real));
  assign _zz_6753 = ($signed(data_mid_3_41_imag) - $signed(data_mid_3_41_real));
  assign _zz_6754 = fixTo_679_dout;
  assign _zz_6755 = _zz_6756[35 : 0];
  assign _zz_6756 = _zz_6757;
  assign _zz_6757 = ($signed(_zz_6758) >>> _zz_569);
  assign _zz_6758 = _zz_6759;
  assign _zz_6759 = ($signed(_zz_6761) - $signed(_zz_566));
  assign _zz_6760 = ({9'd0,data_mid_3_33_real} <<< 9);
  assign _zz_6761 = {{9{_zz_6760[26]}}, _zz_6760};
  assign _zz_6762 = fixTo_680_dout;
  assign _zz_6763 = _zz_6764[35 : 0];
  assign _zz_6764 = _zz_6765;
  assign _zz_6765 = ($signed(_zz_6766) >>> _zz_569);
  assign _zz_6766 = _zz_6767;
  assign _zz_6767 = ($signed(_zz_6769) - $signed(_zz_567));
  assign _zz_6768 = ({9'd0,data_mid_3_33_imag} <<< 9);
  assign _zz_6769 = {{9{_zz_6768[26]}}, _zz_6768};
  assign _zz_6770 = fixTo_681_dout;
  assign _zz_6771 = _zz_6772[35 : 0];
  assign _zz_6772 = _zz_6773;
  assign _zz_6773 = ($signed(_zz_6774) >>> _zz_570);
  assign _zz_6774 = _zz_6775;
  assign _zz_6775 = ($signed(_zz_6777) + $signed(_zz_566));
  assign _zz_6776 = ({9'd0,data_mid_3_33_real} <<< 9);
  assign _zz_6777 = {{9{_zz_6776[26]}}, _zz_6776};
  assign _zz_6778 = fixTo_682_dout;
  assign _zz_6779 = _zz_6780[35 : 0];
  assign _zz_6780 = _zz_6781;
  assign _zz_6781 = ($signed(_zz_6782) >>> _zz_570);
  assign _zz_6782 = _zz_6783;
  assign _zz_6783 = ($signed(_zz_6785) + $signed(_zz_567));
  assign _zz_6784 = ({9'd0,data_mid_3_33_imag} <<< 9);
  assign _zz_6785 = {{9{_zz_6784[26]}}, _zz_6784};
  assign _zz_6786 = fixTo_683_dout;
  assign _zz_6787 = ($signed(twiddle_factor_table_9_real) + $signed(twiddle_factor_table_9_imag));
  assign _zz_6788 = ($signed(_zz_573) - $signed(_zz_6789));
  assign _zz_6789 = ($signed(_zz_6790) * $signed(twiddle_factor_table_9_imag));
  assign _zz_6790 = ($signed(data_mid_3_42_real) + $signed(data_mid_3_42_imag));
  assign _zz_6791 = fixTo_684_dout;
  assign _zz_6792 = ($signed(_zz_573) + $signed(_zz_6793));
  assign _zz_6793 = ($signed(_zz_6794) * $signed(twiddle_factor_table_9_real));
  assign _zz_6794 = ($signed(data_mid_3_42_imag) - $signed(data_mid_3_42_real));
  assign _zz_6795 = fixTo_685_dout;
  assign _zz_6796 = _zz_6797[35 : 0];
  assign _zz_6797 = _zz_6798;
  assign _zz_6798 = ($signed(_zz_6799) >>> _zz_574);
  assign _zz_6799 = _zz_6800;
  assign _zz_6800 = ($signed(_zz_6802) - $signed(_zz_571));
  assign _zz_6801 = ({9'd0,data_mid_3_34_real} <<< 9);
  assign _zz_6802 = {{9{_zz_6801[26]}}, _zz_6801};
  assign _zz_6803 = fixTo_686_dout;
  assign _zz_6804 = _zz_6805[35 : 0];
  assign _zz_6805 = _zz_6806;
  assign _zz_6806 = ($signed(_zz_6807) >>> _zz_574);
  assign _zz_6807 = _zz_6808;
  assign _zz_6808 = ($signed(_zz_6810) - $signed(_zz_572));
  assign _zz_6809 = ({9'd0,data_mid_3_34_imag} <<< 9);
  assign _zz_6810 = {{9{_zz_6809[26]}}, _zz_6809};
  assign _zz_6811 = fixTo_687_dout;
  assign _zz_6812 = _zz_6813[35 : 0];
  assign _zz_6813 = _zz_6814;
  assign _zz_6814 = ($signed(_zz_6815) >>> _zz_575);
  assign _zz_6815 = _zz_6816;
  assign _zz_6816 = ($signed(_zz_6818) + $signed(_zz_571));
  assign _zz_6817 = ({9'd0,data_mid_3_34_real} <<< 9);
  assign _zz_6818 = {{9{_zz_6817[26]}}, _zz_6817};
  assign _zz_6819 = fixTo_688_dout;
  assign _zz_6820 = _zz_6821[35 : 0];
  assign _zz_6821 = _zz_6822;
  assign _zz_6822 = ($signed(_zz_6823) >>> _zz_575);
  assign _zz_6823 = _zz_6824;
  assign _zz_6824 = ($signed(_zz_6826) + $signed(_zz_572));
  assign _zz_6825 = ({9'd0,data_mid_3_34_imag} <<< 9);
  assign _zz_6826 = {{9{_zz_6825[26]}}, _zz_6825};
  assign _zz_6827 = fixTo_689_dout;
  assign _zz_6828 = ($signed(twiddle_factor_table_10_real) + $signed(twiddle_factor_table_10_imag));
  assign _zz_6829 = ($signed(_zz_578) - $signed(_zz_6830));
  assign _zz_6830 = ($signed(_zz_6831) * $signed(twiddle_factor_table_10_imag));
  assign _zz_6831 = ($signed(data_mid_3_43_real) + $signed(data_mid_3_43_imag));
  assign _zz_6832 = fixTo_690_dout;
  assign _zz_6833 = ($signed(_zz_578) + $signed(_zz_6834));
  assign _zz_6834 = ($signed(_zz_6835) * $signed(twiddle_factor_table_10_real));
  assign _zz_6835 = ($signed(data_mid_3_43_imag) - $signed(data_mid_3_43_real));
  assign _zz_6836 = fixTo_691_dout;
  assign _zz_6837 = _zz_6838[35 : 0];
  assign _zz_6838 = _zz_6839;
  assign _zz_6839 = ($signed(_zz_6840) >>> _zz_579);
  assign _zz_6840 = _zz_6841;
  assign _zz_6841 = ($signed(_zz_6843) - $signed(_zz_576));
  assign _zz_6842 = ({9'd0,data_mid_3_35_real} <<< 9);
  assign _zz_6843 = {{9{_zz_6842[26]}}, _zz_6842};
  assign _zz_6844 = fixTo_692_dout;
  assign _zz_6845 = _zz_6846[35 : 0];
  assign _zz_6846 = _zz_6847;
  assign _zz_6847 = ($signed(_zz_6848) >>> _zz_579);
  assign _zz_6848 = _zz_6849;
  assign _zz_6849 = ($signed(_zz_6851) - $signed(_zz_577));
  assign _zz_6850 = ({9'd0,data_mid_3_35_imag} <<< 9);
  assign _zz_6851 = {{9{_zz_6850[26]}}, _zz_6850};
  assign _zz_6852 = fixTo_693_dout;
  assign _zz_6853 = _zz_6854[35 : 0];
  assign _zz_6854 = _zz_6855;
  assign _zz_6855 = ($signed(_zz_6856) >>> _zz_580);
  assign _zz_6856 = _zz_6857;
  assign _zz_6857 = ($signed(_zz_6859) + $signed(_zz_576));
  assign _zz_6858 = ({9'd0,data_mid_3_35_real} <<< 9);
  assign _zz_6859 = {{9{_zz_6858[26]}}, _zz_6858};
  assign _zz_6860 = fixTo_694_dout;
  assign _zz_6861 = _zz_6862[35 : 0];
  assign _zz_6862 = _zz_6863;
  assign _zz_6863 = ($signed(_zz_6864) >>> _zz_580);
  assign _zz_6864 = _zz_6865;
  assign _zz_6865 = ($signed(_zz_6867) + $signed(_zz_577));
  assign _zz_6866 = ({9'd0,data_mid_3_35_imag} <<< 9);
  assign _zz_6867 = {{9{_zz_6866[26]}}, _zz_6866};
  assign _zz_6868 = fixTo_695_dout;
  assign _zz_6869 = ($signed(twiddle_factor_table_11_real) + $signed(twiddle_factor_table_11_imag));
  assign _zz_6870 = ($signed(_zz_583) - $signed(_zz_6871));
  assign _zz_6871 = ($signed(_zz_6872) * $signed(twiddle_factor_table_11_imag));
  assign _zz_6872 = ($signed(data_mid_3_44_real) + $signed(data_mid_3_44_imag));
  assign _zz_6873 = fixTo_696_dout;
  assign _zz_6874 = ($signed(_zz_583) + $signed(_zz_6875));
  assign _zz_6875 = ($signed(_zz_6876) * $signed(twiddle_factor_table_11_real));
  assign _zz_6876 = ($signed(data_mid_3_44_imag) - $signed(data_mid_3_44_real));
  assign _zz_6877 = fixTo_697_dout;
  assign _zz_6878 = _zz_6879[35 : 0];
  assign _zz_6879 = _zz_6880;
  assign _zz_6880 = ($signed(_zz_6881) >>> _zz_584);
  assign _zz_6881 = _zz_6882;
  assign _zz_6882 = ($signed(_zz_6884) - $signed(_zz_581));
  assign _zz_6883 = ({9'd0,data_mid_3_36_real} <<< 9);
  assign _zz_6884 = {{9{_zz_6883[26]}}, _zz_6883};
  assign _zz_6885 = fixTo_698_dout;
  assign _zz_6886 = _zz_6887[35 : 0];
  assign _zz_6887 = _zz_6888;
  assign _zz_6888 = ($signed(_zz_6889) >>> _zz_584);
  assign _zz_6889 = _zz_6890;
  assign _zz_6890 = ($signed(_zz_6892) - $signed(_zz_582));
  assign _zz_6891 = ({9'd0,data_mid_3_36_imag} <<< 9);
  assign _zz_6892 = {{9{_zz_6891[26]}}, _zz_6891};
  assign _zz_6893 = fixTo_699_dout;
  assign _zz_6894 = _zz_6895[35 : 0];
  assign _zz_6895 = _zz_6896;
  assign _zz_6896 = ($signed(_zz_6897) >>> _zz_585);
  assign _zz_6897 = _zz_6898;
  assign _zz_6898 = ($signed(_zz_6900) + $signed(_zz_581));
  assign _zz_6899 = ({9'd0,data_mid_3_36_real} <<< 9);
  assign _zz_6900 = {{9{_zz_6899[26]}}, _zz_6899};
  assign _zz_6901 = fixTo_700_dout;
  assign _zz_6902 = _zz_6903[35 : 0];
  assign _zz_6903 = _zz_6904;
  assign _zz_6904 = ($signed(_zz_6905) >>> _zz_585);
  assign _zz_6905 = _zz_6906;
  assign _zz_6906 = ($signed(_zz_6908) + $signed(_zz_582));
  assign _zz_6907 = ({9'd0,data_mid_3_36_imag} <<< 9);
  assign _zz_6908 = {{9{_zz_6907[26]}}, _zz_6907};
  assign _zz_6909 = fixTo_701_dout;
  assign _zz_6910 = ($signed(twiddle_factor_table_12_real) + $signed(twiddle_factor_table_12_imag));
  assign _zz_6911 = ($signed(_zz_588) - $signed(_zz_6912));
  assign _zz_6912 = ($signed(_zz_6913) * $signed(twiddle_factor_table_12_imag));
  assign _zz_6913 = ($signed(data_mid_3_45_real) + $signed(data_mid_3_45_imag));
  assign _zz_6914 = fixTo_702_dout;
  assign _zz_6915 = ($signed(_zz_588) + $signed(_zz_6916));
  assign _zz_6916 = ($signed(_zz_6917) * $signed(twiddle_factor_table_12_real));
  assign _zz_6917 = ($signed(data_mid_3_45_imag) - $signed(data_mid_3_45_real));
  assign _zz_6918 = fixTo_703_dout;
  assign _zz_6919 = _zz_6920[35 : 0];
  assign _zz_6920 = _zz_6921;
  assign _zz_6921 = ($signed(_zz_6922) >>> _zz_589);
  assign _zz_6922 = _zz_6923;
  assign _zz_6923 = ($signed(_zz_6925) - $signed(_zz_586));
  assign _zz_6924 = ({9'd0,data_mid_3_37_real} <<< 9);
  assign _zz_6925 = {{9{_zz_6924[26]}}, _zz_6924};
  assign _zz_6926 = fixTo_704_dout;
  assign _zz_6927 = _zz_6928[35 : 0];
  assign _zz_6928 = _zz_6929;
  assign _zz_6929 = ($signed(_zz_6930) >>> _zz_589);
  assign _zz_6930 = _zz_6931;
  assign _zz_6931 = ($signed(_zz_6933) - $signed(_zz_587));
  assign _zz_6932 = ({9'd0,data_mid_3_37_imag} <<< 9);
  assign _zz_6933 = {{9{_zz_6932[26]}}, _zz_6932};
  assign _zz_6934 = fixTo_705_dout;
  assign _zz_6935 = _zz_6936[35 : 0];
  assign _zz_6936 = _zz_6937;
  assign _zz_6937 = ($signed(_zz_6938) >>> _zz_590);
  assign _zz_6938 = _zz_6939;
  assign _zz_6939 = ($signed(_zz_6941) + $signed(_zz_586));
  assign _zz_6940 = ({9'd0,data_mid_3_37_real} <<< 9);
  assign _zz_6941 = {{9{_zz_6940[26]}}, _zz_6940};
  assign _zz_6942 = fixTo_706_dout;
  assign _zz_6943 = _zz_6944[35 : 0];
  assign _zz_6944 = _zz_6945;
  assign _zz_6945 = ($signed(_zz_6946) >>> _zz_590);
  assign _zz_6946 = _zz_6947;
  assign _zz_6947 = ($signed(_zz_6949) + $signed(_zz_587));
  assign _zz_6948 = ({9'd0,data_mid_3_37_imag} <<< 9);
  assign _zz_6949 = {{9{_zz_6948[26]}}, _zz_6948};
  assign _zz_6950 = fixTo_707_dout;
  assign _zz_6951 = ($signed(twiddle_factor_table_13_real) + $signed(twiddle_factor_table_13_imag));
  assign _zz_6952 = ($signed(_zz_593) - $signed(_zz_6953));
  assign _zz_6953 = ($signed(_zz_6954) * $signed(twiddle_factor_table_13_imag));
  assign _zz_6954 = ($signed(data_mid_3_46_real) + $signed(data_mid_3_46_imag));
  assign _zz_6955 = fixTo_708_dout;
  assign _zz_6956 = ($signed(_zz_593) + $signed(_zz_6957));
  assign _zz_6957 = ($signed(_zz_6958) * $signed(twiddle_factor_table_13_real));
  assign _zz_6958 = ($signed(data_mid_3_46_imag) - $signed(data_mid_3_46_real));
  assign _zz_6959 = fixTo_709_dout;
  assign _zz_6960 = _zz_6961[35 : 0];
  assign _zz_6961 = _zz_6962;
  assign _zz_6962 = ($signed(_zz_6963) >>> _zz_594);
  assign _zz_6963 = _zz_6964;
  assign _zz_6964 = ($signed(_zz_6966) - $signed(_zz_591));
  assign _zz_6965 = ({9'd0,data_mid_3_38_real} <<< 9);
  assign _zz_6966 = {{9{_zz_6965[26]}}, _zz_6965};
  assign _zz_6967 = fixTo_710_dout;
  assign _zz_6968 = _zz_6969[35 : 0];
  assign _zz_6969 = _zz_6970;
  assign _zz_6970 = ($signed(_zz_6971) >>> _zz_594);
  assign _zz_6971 = _zz_6972;
  assign _zz_6972 = ($signed(_zz_6974) - $signed(_zz_592));
  assign _zz_6973 = ({9'd0,data_mid_3_38_imag} <<< 9);
  assign _zz_6974 = {{9{_zz_6973[26]}}, _zz_6973};
  assign _zz_6975 = fixTo_711_dout;
  assign _zz_6976 = _zz_6977[35 : 0];
  assign _zz_6977 = _zz_6978;
  assign _zz_6978 = ($signed(_zz_6979) >>> _zz_595);
  assign _zz_6979 = _zz_6980;
  assign _zz_6980 = ($signed(_zz_6982) + $signed(_zz_591));
  assign _zz_6981 = ({9'd0,data_mid_3_38_real} <<< 9);
  assign _zz_6982 = {{9{_zz_6981[26]}}, _zz_6981};
  assign _zz_6983 = fixTo_712_dout;
  assign _zz_6984 = _zz_6985[35 : 0];
  assign _zz_6985 = _zz_6986;
  assign _zz_6986 = ($signed(_zz_6987) >>> _zz_595);
  assign _zz_6987 = _zz_6988;
  assign _zz_6988 = ($signed(_zz_6990) + $signed(_zz_592));
  assign _zz_6989 = ({9'd0,data_mid_3_38_imag} <<< 9);
  assign _zz_6990 = {{9{_zz_6989[26]}}, _zz_6989};
  assign _zz_6991 = fixTo_713_dout;
  assign _zz_6992 = ($signed(twiddle_factor_table_14_real) + $signed(twiddle_factor_table_14_imag));
  assign _zz_6993 = ($signed(_zz_598) - $signed(_zz_6994));
  assign _zz_6994 = ($signed(_zz_6995) * $signed(twiddle_factor_table_14_imag));
  assign _zz_6995 = ($signed(data_mid_3_47_real) + $signed(data_mid_3_47_imag));
  assign _zz_6996 = fixTo_714_dout;
  assign _zz_6997 = ($signed(_zz_598) + $signed(_zz_6998));
  assign _zz_6998 = ($signed(_zz_6999) * $signed(twiddle_factor_table_14_real));
  assign _zz_6999 = ($signed(data_mid_3_47_imag) - $signed(data_mid_3_47_real));
  assign _zz_7000 = fixTo_715_dout;
  assign _zz_7001 = _zz_7002[35 : 0];
  assign _zz_7002 = _zz_7003;
  assign _zz_7003 = ($signed(_zz_7004) >>> _zz_599);
  assign _zz_7004 = _zz_7005;
  assign _zz_7005 = ($signed(_zz_7007) - $signed(_zz_596));
  assign _zz_7006 = ({9'd0,data_mid_3_39_real} <<< 9);
  assign _zz_7007 = {{9{_zz_7006[26]}}, _zz_7006};
  assign _zz_7008 = fixTo_716_dout;
  assign _zz_7009 = _zz_7010[35 : 0];
  assign _zz_7010 = _zz_7011;
  assign _zz_7011 = ($signed(_zz_7012) >>> _zz_599);
  assign _zz_7012 = _zz_7013;
  assign _zz_7013 = ($signed(_zz_7015) - $signed(_zz_597));
  assign _zz_7014 = ({9'd0,data_mid_3_39_imag} <<< 9);
  assign _zz_7015 = {{9{_zz_7014[26]}}, _zz_7014};
  assign _zz_7016 = fixTo_717_dout;
  assign _zz_7017 = _zz_7018[35 : 0];
  assign _zz_7018 = _zz_7019;
  assign _zz_7019 = ($signed(_zz_7020) >>> _zz_600);
  assign _zz_7020 = _zz_7021;
  assign _zz_7021 = ($signed(_zz_7023) + $signed(_zz_596));
  assign _zz_7022 = ({9'd0,data_mid_3_39_real} <<< 9);
  assign _zz_7023 = {{9{_zz_7022[26]}}, _zz_7022};
  assign _zz_7024 = fixTo_718_dout;
  assign _zz_7025 = _zz_7026[35 : 0];
  assign _zz_7026 = _zz_7027;
  assign _zz_7027 = ($signed(_zz_7028) >>> _zz_600);
  assign _zz_7028 = _zz_7029;
  assign _zz_7029 = ($signed(_zz_7031) + $signed(_zz_597));
  assign _zz_7030 = ({9'd0,data_mid_3_39_imag} <<< 9);
  assign _zz_7031 = {{9{_zz_7030[26]}}, _zz_7030};
  assign _zz_7032 = fixTo_719_dout;
  assign _zz_7033 = ($signed(twiddle_factor_table_7_real) + $signed(twiddle_factor_table_7_imag));
  assign _zz_7034 = ($signed(_zz_603) - $signed(_zz_7035));
  assign _zz_7035 = ($signed(_zz_7036) * $signed(twiddle_factor_table_7_imag));
  assign _zz_7036 = ($signed(data_mid_3_56_real) + $signed(data_mid_3_56_imag));
  assign _zz_7037 = fixTo_720_dout;
  assign _zz_7038 = ($signed(_zz_603) + $signed(_zz_7039));
  assign _zz_7039 = ($signed(_zz_7040) * $signed(twiddle_factor_table_7_real));
  assign _zz_7040 = ($signed(data_mid_3_56_imag) - $signed(data_mid_3_56_real));
  assign _zz_7041 = fixTo_721_dout;
  assign _zz_7042 = _zz_7043[35 : 0];
  assign _zz_7043 = _zz_7044;
  assign _zz_7044 = ($signed(_zz_7045) >>> _zz_604);
  assign _zz_7045 = _zz_7046;
  assign _zz_7046 = ($signed(_zz_7048) - $signed(_zz_601));
  assign _zz_7047 = ({9'd0,data_mid_3_48_real} <<< 9);
  assign _zz_7048 = {{9{_zz_7047[26]}}, _zz_7047};
  assign _zz_7049 = fixTo_722_dout;
  assign _zz_7050 = _zz_7051[35 : 0];
  assign _zz_7051 = _zz_7052;
  assign _zz_7052 = ($signed(_zz_7053) >>> _zz_604);
  assign _zz_7053 = _zz_7054;
  assign _zz_7054 = ($signed(_zz_7056) - $signed(_zz_602));
  assign _zz_7055 = ({9'd0,data_mid_3_48_imag} <<< 9);
  assign _zz_7056 = {{9{_zz_7055[26]}}, _zz_7055};
  assign _zz_7057 = fixTo_723_dout;
  assign _zz_7058 = _zz_7059[35 : 0];
  assign _zz_7059 = _zz_7060;
  assign _zz_7060 = ($signed(_zz_7061) >>> _zz_605);
  assign _zz_7061 = _zz_7062;
  assign _zz_7062 = ($signed(_zz_7064) + $signed(_zz_601));
  assign _zz_7063 = ({9'd0,data_mid_3_48_real} <<< 9);
  assign _zz_7064 = {{9{_zz_7063[26]}}, _zz_7063};
  assign _zz_7065 = fixTo_724_dout;
  assign _zz_7066 = _zz_7067[35 : 0];
  assign _zz_7067 = _zz_7068;
  assign _zz_7068 = ($signed(_zz_7069) >>> _zz_605);
  assign _zz_7069 = _zz_7070;
  assign _zz_7070 = ($signed(_zz_7072) + $signed(_zz_602));
  assign _zz_7071 = ({9'd0,data_mid_3_48_imag} <<< 9);
  assign _zz_7072 = {{9{_zz_7071[26]}}, _zz_7071};
  assign _zz_7073 = fixTo_725_dout;
  assign _zz_7074 = ($signed(twiddle_factor_table_8_real) + $signed(twiddle_factor_table_8_imag));
  assign _zz_7075 = ($signed(_zz_608) - $signed(_zz_7076));
  assign _zz_7076 = ($signed(_zz_7077) * $signed(twiddle_factor_table_8_imag));
  assign _zz_7077 = ($signed(data_mid_3_57_real) + $signed(data_mid_3_57_imag));
  assign _zz_7078 = fixTo_726_dout;
  assign _zz_7079 = ($signed(_zz_608) + $signed(_zz_7080));
  assign _zz_7080 = ($signed(_zz_7081) * $signed(twiddle_factor_table_8_real));
  assign _zz_7081 = ($signed(data_mid_3_57_imag) - $signed(data_mid_3_57_real));
  assign _zz_7082 = fixTo_727_dout;
  assign _zz_7083 = _zz_7084[35 : 0];
  assign _zz_7084 = _zz_7085;
  assign _zz_7085 = ($signed(_zz_7086) >>> _zz_609);
  assign _zz_7086 = _zz_7087;
  assign _zz_7087 = ($signed(_zz_7089) - $signed(_zz_606));
  assign _zz_7088 = ({9'd0,data_mid_3_49_real} <<< 9);
  assign _zz_7089 = {{9{_zz_7088[26]}}, _zz_7088};
  assign _zz_7090 = fixTo_728_dout;
  assign _zz_7091 = _zz_7092[35 : 0];
  assign _zz_7092 = _zz_7093;
  assign _zz_7093 = ($signed(_zz_7094) >>> _zz_609);
  assign _zz_7094 = _zz_7095;
  assign _zz_7095 = ($signed(_zz_7097) - $signed(_zz_607));
  assign _zz_7096 = ({9'd0,data_mid_3_49_imag} <<< 9);
  assign _zz_7097 = {{9{_zz_7096[26]}}, _zz_7096};
  assign _zz_7098 = fixTo_729_dout;
  assign _zz_7099 = _zz_7100[35 : 0];
  assign _zz_7100 = _zz_7101;
  assign _zz_7101 = ($signed(_zz_7102) >>> _zz_610);
  assign _zz_7102 = _zz_7103;
  assign _zz_7103 = ($signed(_zz_7105) + $signed(_zz_606));
  assign _zz_7104 = ({9'd0,data_mid_3_49_real} <<< 9);
  assign _zz_7105 = {{9{_zz_7104[26]}}, _zz_7104};
  assign _zz_7106 = fixTo_730_dout;
  assign _zz_7107 = _zz_7108[35 : 0];
  assign _zz_7108 = _zz_7109;
  assign _zz_7109 = ($signed(_zz_7110) >>> _zz_610);
  assign _zz_7110 = _zz_7111;
  assign _zz_7111 = ($signed(_zz_7113) + $signed(_zz_607));
  assign _zz_7112 = ({9'd0,data_mid_3_49_imag} <<< 9);
  assign _zz_7113 = {{9{_zz_7112[26]}}, _zz_7112};
  assign _zz_7114 = fixTo_731_dout;
  assign _zz_7115 = ($signed(twiddle_factor_table_9_real) + $signed(twiddle_factor_table_9_imag));
  assign _zz_7116 = ($signed(_zz_613) - $signed(_zz_7117));
  assign _zz_7117 = ($signed(_zz_7118) * $signed(twiddle_factor_table_9_imag));
  assign _zz_7118 = ($signed(data_mid_3_58_real) + $signed(data_mid_3_58_imag));
  assign _zz_7119 = fixTo_732_dout;
  assign _zz_7120 = ($signed(_zz_613) + $signed(_zz_7121));
  assign _zz_7121 = ($signed(_zz_7122) * $signed(twiddle_factor_table_9_real));
  assign _zz_7122 = ($signed(data_mid_3_58_imag) - $signed(data_mid_3_58_real));
  assign _zz_7123 = fixTo_733_dout;
  assign _zz_7124 = _zz_7125[35 : 0];
  assign _zz_7125 = _zz_7126;
  assign _zz_7126 = ($signed(_zz_7127) >>> _zz_614);
  assign _zz_7127 = _zz_7128;
  assign _zz_7128 = ($signed(_zz_7130) - $signed(_zz_611));
  assign _zz_7129 = ({9'd0,data_mid_3_50_real} <<< 9);
  assign _zz_7130 = {{9{_zz_7129[26]}}, _zz_7129};
  assign _zz_7131 = fixTo_734_dout;
  assign _zz_7132 = _zz_7133[35 : 0];
  assign _zz_7133 = _zz_7134;
  assign _zz_7134 = ($signed(_zz_7135) >>> _zz_614);
  assign _zz_7135 = _zz_7136;
  assign _zz_7136 = ($signed(_zz_7138) - $signed(_zz_612));
  assign _zz_7137 = ({9'd0,data_mid_3_50_imag} <<< 9);
  assign _zz_7138 = {{9{_zz_7137[26]}}, _zz_7137};
  assign _zz_7139 = fixTo_735_dout;
  assign _zz_7140 = _zz_7141[35 : 0];
  assign _zz_7141 = _zz_7142;
  assign _zz_7142 = ($signed(_zz_7143) >>> _zz_615);
  assign _zz_7143 = _zz_7144;
  assign _zz_7144 = ($signed(_zz_7146) + $signed(_zz_611));
  assign _zz_7145 = ({9'd0,data_mid_3_50_real} <<< 9);
  assign _zz_7146 = {{9{_zz_7145[26]}}, _zz_7145};
  assign _zz_7147 = fixTo_736_dout;
  assign _zz_7148 = _zz_7149[35 : 0];
  assign _zz_7149 = _zz_7150;
  assign _zz_7150 = ($signed(_zz_7151) >>> _zz_615);
  assign _zz_7151 = _zz_7152;
  assign _zz_7152 = ($signed(_zz_7154) + $signed(_zz_612));
  assign _zz_7153 = ({9'd0,data_mid_3_50_imag} <<< 9);
  assign _zz_7154 = {{9{_zz_7153[26]}}, _zz_7153};
  assign _zz_7155 = fixTo_737_dout;
  assign _zz_7156 = ($signed(twiddle_factor_table_10_real) + $signed(twiddle_factor_table_10_imag));
  assign _zz_7157 = ($signed(_zz_618) - $signed(_zz_7158));
  assign _zz_7158 = ($signed(_zz_7159) * $signed(twiddle_factor_table_10_imag));
  assign _zz_7159 = ($signed(data_mid_3_59_real) + $signed(data_mid_3_59_imag));
  assign _zz_7160 = fixTo_738_dout;
  assign _zz_7161 = ($signed(_zz_618) + $signed(_zz_7162));
  assign _zz_7162 = ($signed(_zz_7163) * $signed(twiddle_factor_table_10_real));
  assign _zz_7163 = ($signed(data_mid_3_59_imag) - $signed(data_mid_3_59_real));
  assign _zz_7164 = fixTo_739_dout;
  assign _zz_7165 = _zz_7166[35 : 0];
  assign _zz_7166 = _zz_7167;
  assign _zz_7167 = ($signed(_zz_7168) >>> _zz_619);
  assign _zz_7168 = _zz_7169;
  assign _zz_7169 = ($signed(_zz_7171) - $signed(_zz_616));
  assign _zz_7170 = ({9'd0,data_mid_3_51_real} <<< 9);
  assign _zz_7171 = {{9{_zz_7170[26]}}, _zz_7170};
  assign _zz_7172 = fixTo_740_dout;
  assign _zz_7173 = _zz_7174[35 : 0];
  assign _zz_7174 = _zz_7175;
  assign _zz_7175 = ($signed(_zz_7176) >>> _zz_619);
  assign _zz_7176 = _zz_7177;
  assign _zz_7177 = ($signed(_zz_7179) - $signed(_zz_617));
  assign _zz_7178 = ({9'd0,data_mid_3_51_imag} <<< 9);
  assign _zz_7179 = {{9{_zz_7178[26]}}, _zz_7178};
  assign _zz_7180 = fixTo_741_dout;
  assign _zz_7181 = _zz_7182[35 : 0];
  assign _zz_7182 = _zz_7183;
  assign _zz_7183 = ($signed(_zz_7184) >>> _zz_620);
  assign _zz_7184 = _zz_7185;
  assign _zz_7185 = ($signed(_zz_7187) + $signed(_zz_616));
  assign _zz_7186 = ({9'd0,data_mid_3_51_real} <<< 9);
  assign _zz_7187 = {{9{_zz_7186[26]}}, _zz_7186};
  assign _zz_7188 = fixTo_742_dout;
  assign _zz_7189 = _zz_7190[35 : 0];
  assign _zz_7190 = _zz_7191;
  assign _zz_7191 = ($signed(_zz_7192) >>> _zz_620);
  assign _zz_7192 = _zz_7193;
  assign _zz_7193 = ($signed(_zz_7195) + $signed(_zz_617));
  assign _zz_7194 = ({9'd0,data_mid_3_51_imag} <<< 9);
  assign _zz_7195 = {{9{_zz_7194[26]}}, _zz_7194};
  assign _zz_7196 = fixTo_743_dout;
  assign _zz_7197 = ($signed(twiddle_factor_table_11_real) + $signed(twiddle_factor_table_11_imag));
  assign _zz_7198 = ($signed(_zz_623) - $signed(_zz_7199));
  assign _zz_7199 = ($signed(_zz_7200) * $signed(twiddle_factor_table_11_imag));
  assign _zz_7200 = ($signed(data_mid_3_60_real) + $signed(data_mid_3_60_imag));
  assign _zz_7201 = fixTo_744_dout;
  assign _zz_7202 = ($signed(_zz_623) + $signed(_zz_7203));
  assign _zz_7203 = ($signed(_zz_7204) * $signed(twiddle_factor_table_11_real));
  assign _zz_7204 = ($signed(data_mid_3_60_imag) - $signed(data_mid_3_60_real));
  assign _zz_7205 = fixTo_745_dout;
  assign _zz_7206 = _zz_7207[35 : 0];
  assign _zz_7207 = _zz_7208;
  assign _zz_7208 = ($signed(_zz_7209) >>> _zz_624);
  assign _zz_7209 = _zz_7210;
  assign _zz_7210 = ($signed(_zz_7212) - $signed(_zz_621));
  assign _zz_7211 = ({9'd0,data_mid_3_52_real} <<< 9);
  assign _zz_7212 = {{9{_zz_7211[26]}}, _zz_7211};
  assign _zz_7213 = fixTo_746_dout;
  assign _zz_7214 = _zz_7215[35 : 0];
  assign _zz_7215 = _zz_7216;
  assign _zz_7216 = ($signed(_zz_7217) >>> _zz_624);
  assign _zz_7217 = _zz_7218;
  assign _zz_7218 = ($signed(_zz_7220) - $signed(_zz_622));
  assign _zz_7219 = ({9'd0,data_mid_3_52_imag} <<< 9);
  assign _zz_7220 = {{9{_zz_7219[26]}}, _zz_7219};
  assign _zz_7221 = fixTo_747_dout;
  assign _zz_7222 = _zz_7223[35 : 0];
  assign _zz_7223 = _zz_7224;
  assign _zz_7224 = ($signed(_zz_7225) >>> _zz_625);
  assign _zz_7225 = _zz_7226;
  assign _zz_7226 = ($signed(_zz_7228) + $signed(_zz_621));
  assign _zz_7227 = ({9'd0,data_mid_3_52_real} <<< 9);
  assign _zz_7228 = {{9{_zz_7227[26]}}, _zz_7227};
  assign _zz_7229 = fixTo_748_dout;
  assign _zz_7230 = _zz_7231[35 : 0];
  assign _zz_7231 = _zz_7232;
  assign _zz_7232 = ($signed(_zz_7233) >>> _zz_625);
  assign _zz_7233 = _zz_7234;
  assign _zz_7234 = ($signed(_zz_7236) + $signed(_zz_622));
  assign _zz_7235 = ({9'd0,data_mid_3_52_imag} <<< 9);
  assign _zz_7236 = {{9{_zz_7235[26]}}, _zz_7235};
  assign _zz_7237 = fixTo_749_dout;
  assign _zz_7238 = ($signed(twiddle_factor_table_12_real) + $signed(twiddle_factor_table_12_imag));
  assign _zz_7239 = ($signed(_zz_628) - $signed(_zz_7240));
  assign _zz_7240 = ($signed(_zz_7241) * $signed(twiddle_factor_table_12_imag));
  assign _zz_7241 = ($signed(data_mid_3_61_real) + $signed(data_mid_3_61_imag));
  assign _zz_7242 = fixTo_750_dout;
  assign _zz_7243 = ($signed(_zz_628) + $signed(_zz_7244));
  assign _zz_7244 = ($signed(_zz_7245) * $signed(twiddle_factor_table_12_real));
  assign _zz_7245 = ($signed(data_mid_3_61_imag) - $signed(data_mid_3_61_real));
  assign _zz_7246 = fixTo_751_dout;
  assign _zz_7247 = _zz_7248[35 : 0];
  assign _zz_7248 = _zz_7249;
  assign _zz_7249 = ($signed(_zz_7250) >>> _zz_629);
  assign _zz_7250 = _zz_7251;
  assign _zz_7251 = ($signed(_zz_7253) - $signed(_zz_626));
  assign _zz_7252 = ({9'd0,data_mid_3_53_real} <<< 9);
  assign _zz_7253 = {{9{_zz_7252[26]}}, _zz_7252};
  assign _zz_7254 = fixTo_752_dout;
  assign _zz_7255 = _zz_7256[35 : 0];
  assign _zz_7256 = _zz_7257;
  assign _zz_7257 = ($signed(_zz_7258) >>> _zz_629);
  assign _zz_7258 = _zz_7259;
  assign _zz_7259 = ($signed(_zz_7261) - $signed(_zz_627));
  assign _zz_7260 = ({9'd0,data_mid_3_53_imag} <<< 9);
  assign _zz_7261 = {{9{_zz_7260[26]}}, _zz_7260};
  assign _zz_7262 = fixTo_753_dout;
  assign _zz_7263 = _zz_7264[35 : 0];
  assign _zz_7264 = _zz_7265;
  assign _zz_7265 = ($signed(_zz_7266) >>> _zz_630);
  assign _zz_7266 = _zz_7267;
  assign _zz_7267 = ($signed(_zz_7269) + $signed(_zz_626));
  assign _zz_7268 = ({9'd0,data_mid_3_53_real} <<< 9);
  assign _zz_7269 = {{9{_zz_7268[26]}}, _zz_7268};
  assign _zz_7270 = fixTo_754_dout;
  assign _zz_7271 = _zz_7272[35 : 0];
  assign _zz_7272 = _zz_7273;
  assign _zz_7273 = ($signed(_zz_7274) >>> _zz_630);
  assign _zz_7274 = _zz_7275;
  assign _zz_7275 = ($signed(_zz_7277) + $signed(_zz_627));
  assign _zz_7276 = ({9'd0,data_mid_3_53_imag} <<< 9);
  assign _zz_7277 = {{9{_zz_7276[26]}}, _zz_7276};
  assign _zz_7278 = fixTo_755_dout;
  assign _zz_7279 = ($signed(twiddle_factor_table_13_real) + $signed(twiddle_factor_table_13_imag));
  assign _zz_7280 = ($signed(_zz_633) - $signed(_zz_7281));
  assign _zz_7281 = ($signed(_zz_7282) * $signed(twiddle_factor_table_13_imag));
  assign _zz_7282 = ($signed(data_mid_3_62_real) + $signed(data_mid_3_62_imag));
  assign _zz_7283 = fixTo_756_dout;
  assign _zz_7284 = ($signed(_zz_633) + $signed(_zz_7285));
  assign _zz_7285 = ($signed(_zz_7286) * $signed(twiddle_factor_table_13_real));
  assign _zz_7286 = ($signed(data_mid_3_62_imag) - $signed(data_mid_3_62_real));
  assign _zz_7287 = fixTo_757_dout;
  assign _zz_7288 = _zz_7289[35 : 0];
  assign _zz_7289 = _zz_7290;
  assign _zz_7290 = ($signed(_zz_7291) >>> _zz_634);
  assign _zz_7291 = _zz_7292;
  assign _zz_7292 = ($signed(_zz_7294) - $signed(_zz_631));
  assign _zz_7293 = ({9'd0,data_mid_3_54_real} <<< 9);
  assign _zz_7294 = {{9{_zz_7293[26]}}, _zz_7293};
  assign _zz_7295 = fixTo_758_dout;
  assign _zz_7296 = _zz_7297[35 : 0];
  assign _zz_7297 = _zz_7298;
  assign _zz_7298 = ($signed(_zz_7299) >>> _zz_634);
  assign _zz_7299 = _zz_7300;
  assign _zz_7300 = ($signed(_zz_7302) - $signed(_zz_632));
  assign _zz_7301 = ({9'd0,data_mid_3_54_imag} <<< 9);
  assign _zz_7302 = {{9{_zz_7301[26]}}, _zz_7301};
  assign _zz_7303 = fixTo_759_dout;
  assign _zz_7304 = _zz_7305[35 : 0];
  assign _zz_7305 = _zz_7306;
  assign _zz_7306 = ($signed(_zz_7307) >>> _zz_635);
  assign _zz_7307 = _zz_7308;
  assign _zz_7308 = ($signed(_zz_7310) + $signed(_zz_631));
  assign _zz_7309 = ({9'd0,data_mid_3_54_real} <<< 9);
  assign _zz_7310 = {{9{_zz_7309[26]}}, _zz_7309};
  assign _zz_7311 = fixTo_760_dout;
  assign _zz_7312 = _zz_7313[35 : 0];
  assign _zz_7313 = _zz_7314;
  assign _zz_7314 = ($signed(_zz_7315) >>> _zz_635);
  assign _zz_7315 = _zz_7316;
  assign _zz_7316 = ($signed(_zz_7318) + $signed(_zz_632));
  assign _zz_7317 = ({9'd0,data_mid_3_54_imag} <<< 9);
  assign _zz_7318 = {{9{_zz_7317[26]}}, _zz_7317};
  assign _zz_7319 = fixTo_761_dout;
  assign _zz_7320 = ($signed(twiddle_factor_table_14_real) + $signed(twiddle_factor_table_14_imag));
  assign _zz_7321 = ($signed(_zz_638) - $signed(_zz_7322));
  assign _zz_7322 = ($signed(_zz_7323) * $signed(twiddle_factor_table_14_imag));
  assign _zz_7323 = ($signed(data_mid_3_63_real) + $signed(data_mid_3_63_imag));
  assign _zz_7324 = fixTo_762_dout;
  assign _zz_7325 = ($signed(_zz_638) + $signed(_zz_7326));
  assign _zz_7326 = ($signed(_zz_7327) * $signed(twiddle_factor_table_14_real));
  assign _zz_7327 = ($signed(data_mid_3_63_imag) - $signed(data_mid_3_63_real));
  assign _zz_7328 = fixTo_763_dout;
  assign _zz_7329 = _zz_7330[35 : 0];
  assign _zz_7330 = _zz_7331;
  assign _zz_7331 = ($signed(_zz_7332) >>> _zz_639);
  assign _zz_7332 = _zz_7333;
  assign _zz_7333 = ($signed(_zz_7335) - $signed(_zz_636));
  assign _zz_7334 = ({9'd0,data_mid_3_55_real} <<< 9);
  assign _zz_7335 = {{9{_zz_7334[26]}}, _zz_7334};
  assign _zz_7336 = fixTo_764_dout;
  assign _zz_7337 = _zz_7338[35 : 0];
  assign _zz_7338 = _zz_7339;
  assign _zz_7339 = ($signed(_zz_7340) >>> _zz_639);
  assign _zz_7340 = _zz_7341;
  assign _zz_7341 = ($signed(_zz_7343) - $signed(_zz_637));
  assign _zz_7342 = ({9'd0,data_mid_3_55_imag} <<< 9);
  assign _zz_7343 = {{9{_zz_7342[26]}}, _zz_7342};
  assign _zz_7344 = fixTo_765_dout;
  assign _zz_7345 = _zz_7346[35 : 0];
  assign _zz_7346 = _zz_7347;
  assign _zz_7347 = ($signed(_zz_7348) >>> _zz_640);
  assign _zz_7348 = _zz_7349;
  assign _zz_7349 = ($signed(_zz_7351) + $signed(_zz_636));
  assign _zz_7350 = ({9'd0,data_mid_3_55_real} <<< 9);
  assign _zz_7351 = {{9{_zz_7350[26]}}, _zz_7350};
  assign _zz_7352 = fixTo_766_dout;
  assign _zz_7353 = _zz_7354[35 : 0];
  assign _zz_7354 = _zz_7355;
  assign _zz_7355 = ($signed(_zz_7356) >>> _zz_640);
  assign _zz_7356 = _zz_7357;
  assign _zz_7357 = ($signed(_zz_7359) + $signed(_zz_637));
  assign _zz_7358 = ({9'd0,data_mid_3_55_imag} <<< 9);
  assign _zz_7359 = {{9{_zz_7358[26]}}, _zz_7358};
  assign _zz_7360 = fixTo_767_dout;
  assign _zz_7361 = ($signed(twiddle_factor_table_15_real) + $signed(twiddle_factor_table_15_imag));
  assign _zz_7362 = ($signed(_zz_643) - $signed(_zz_7363));
  assign _zz_7363 = ($signed(_zz_7364) * $signed(twiddle_factor_table_15_imag));
  assign _zz_7364 = ($signed(data_mid_4_16_real) + $signed(data_mid_4_16_imag));
  assign _zz_7365 = fixTo_768_dout;
  assign _zz_7366 = ($signed(_zz_643) + $signed(_zz_7367));
  assign _zz_7367 = ($signed(_zz_7368) * $signed(twiddle_factor_table_15_real));
  assign _zz_7368 = ($signed(data_mid_4_16_imag) - $signed(data_mid_4_16_real));
  assign _zz_7369 = fixTo_769_dout;
  assign _zz_7370 = _zz_7371[35 : 0];
  assign _zz_7371 = _zz_7372;
  assign _zz_7372 = ($signed(_zz_7373) >>> _zz_644);
  assign _zz_7373 = _zz_7374;
  assign _zz_7374 = ($signed(_zz_7376) - $signed(_zz_641));
  assign _zz_7375 = ({9'd0,data_mid_4_0_real} <<< 9);
  assign _zz_7376 = {{9{_zz_7375[26]}}, _zz_7375};
  assign _zz_7377 = fixTo_770_dout;
  assign _zz_7378 = _zz_7379[35 : 0];
  assign _zz_7379 = _zz_7380;
  assign _zz_7380 = ($signed(_zz_7381) >>> _zz_644);
  assign _zz_7381 = _zz_7382;
  assign _zz_7382 = ($signed(_zz_7384) - $signed(_zz_642));
  assign _zz_7383 = ({9'd0,data_mid_4_0_imag} <<< 9);
  assign _zz_7384 = {{9{_zz_7383[26]}}, _zz_7383};
  assign _zz_7385 = fixTo_771_dout;
  assign _zz_7386 = _zz_7387[35 : 0];
  assign _zz_7387 = _zz_7388;
  assign _zz_7388 = ($signed(_zz_7389) >>> _zz_645);
  assign _zz_7389 = _zz_7390;
  assign _zz_7390 = ($signed(_zz_7392) + $signed(_zz_641));
  assign _zz_7391 = ({9'd0,data_mid_4_0_real} <<< 9);
  assign _zz_7392 = {{9{_zz_7391[26]}}, _zz_7391};
  assign _zz_7393 = fixTo_772_dout;
  assign _zz_7394 = _zz_7395[35 : 0];
  assign _zz_7395 = _zz_7396;
  assign _zz_7396 = ($signed(_zz_7397) >>> _zz_645);
  assign _zz_7397 = _zz_7398;
  assign _zz_7398 = ($signed(_zz_7400) + $signed(_zz_642));
  assign _zz_7399 = ({9'd0,data_mid_4_0_imag} <<< 9);
  assign _zz_7400 = {{9{_zz_7399[26]}}, _zz_7399};
  assign _zz_7401 = fixTo_773_dout;
  assign _zz_7402 = ($signed(twiddle_factor_table_16_real) + $signed(twiddle_factor_table_16_imag));
  assign _zz_7403 = ($signed(_zz_648) - $signed(_zz_7404));
  assign _zz_7404 = ($signed(_zz_7405) * $signed(twiddle_factor_table_16_imag));
  assign _zz_7405 = ($signed(data_mid_4_17_real) + $signed(data_mid_4_17_imag));
  assign _zz_7406 = fixTo_774_dout;
  assign _zz_7407 = ($signed(_zz_648) + $signed(_zz_7408));
  assign _zz_7408 = ($signed(_zz_7409) * $signed(twiddle_factor_table_16_real));
  assign _zz_7409 = ($signed(data_mid_4_17_imag) - $signed(data_mid_4_17_real));
  assign _zz_7410 = fixTo_775_dout;
  assign _zz_7411 = _zz_7412[35 : 0];
  assign _zz_7412 = _zz_7413;
  assign _zz_7413 = ($signed(_zz_7414) >>> _zz_649);
  assign _zz_7414 = _zz_7415;
  assign _zz_7415 = ($signed(_zz_7417) - $signed(_zz_646));
  assign _zz_7416 = ({9'd0,data_mid_4_1_real} <<< 9);
  assign _zz_7417 = {{9{_zz_7416[26]}}, _zz_7416};
  assign _zz_7418 = fixTo_776_dout;
  assign _zz_7419 = _zz_7420[35 : 0];
  assign _zz_7420 = _zz_7421;
  assign _zz_7421 = ($signed(_zz_7422) >>> _zz_649);
  assign _zz_7422 = _zz_7423;
  assign _zz_7423 = ($signed(_zz_7425) - $signed(_zz_647));
  assign _zz_7424 = ({9'd0,data_mid_4_1_imag} <<< 9);
  assign _zz_7425 = {{9{_zz_7424[26]}}, _zz_7424};
  assign _zz_7426 = fixTo_777_dout;
  assign _zz_7427 = _zz_7428[35 : 0];
  assign _zz_7428 = _zz_7429;
  assign _zz_7429 = ($signed(_zz_7430) >>> _zz_650);
  assign _zz_7430 = _zz_7431;
  assign _zz_7431 = ($signed(_zz_7433) + $signed(_zz_646));
  assign _zz_7432 = ({9'd0,data_mid_4_1_real} <<< 9);
  assign _zz_7433 = {{9{_zz_7432[26]}}, _zz_7432};
  assign _zz_7434 = fixTo_778_dout;
  assign _zz_7435 = _zz_7436[35 : 0];
  assign _zz_7436 = _zz_7437;
  assign _zz_7437 = ($signed(_zz_7438) >>> _zz_650);
  assign _zz_7438 = _zz_7439;
  assign _zz_7439 = ($signed(_zz_7441) + $signed(_zz_647));
  assign _zz_7440 = ({9'd0,data_mid_4_1_imag} <<< 9);
  assign _zz_7441 = {{9{_zz_7440[26]}}, _zz_7440};
  assign _zz_7442 = fixTo_779_dout;
  assign _zz_7443 = ($signed(twiddle_factor_table_17_real) + $signed(twiddle_factor_table_17_imag));
  assign _zz_7444 = ($signed(_zz_653) - $signed(_zz_7445));
  assign _zz_7445 = ($signed(_zz_7446) * $signed(twiddle_factor_table_17_imag));
  assign _zz_7446 = ($signed(data_mid_4_18_real) + $signed(data_mid_4_18_imag));
  assign _zz_7447 = fixTo_780_dout;
  assign _zz_7448 = ($signed(_zz_653) + $signed(_zz_7449));
  assign _zz_7449 = ($signed(_zz_7450) * $signed(twiddle_factor_table_17_real));
  assign _zz_7450 = ($signed(data_mid_4_18_imag) - $signed(data_mid_4_18_real));
  assign _zz_7451 = fixTo_781_dout;
  assign _zz_7452 = _zz_7453[35 : 0];
  assign _zz_7453 = _zz_7454;
  assign _zz_7454 = ($signed(_zz_7455) >>> _zz_654);
  assign _zz_7455 = _zz_7456;
  assign _zz_7456 = ($signed(_zz_7458) - $signed(_zz_651));
  assign _zz_7457 = ({9'd0,data_mid_4_2_real} <<< 9);
  assign _zz_7458 = {{9{_zz_7457[26]}}, _zz_7457};
  assign _zz_7459 = fixTo_782_dout;
  assign _zz_7460 = _zz_7461[35 : 0];
  assign _zz_7461 = _zz_7462;
  assign _zz_7462 = ($signed(_zz_7463) >>> _zz_654);
  assign _zz_7463 = _zz_7464;
  assign _zz_7464 = ($signed(_zz_7466) - $signed(_zz_652));
  assign _zz_7465 = ({9'd0,data_mid_4_2_imag} <<< 9);
  assign _zz_7466 = {{9{_zz_7465[26]}}, _zz_7465};
  assign _zz_7467 = fixTo_783_dout;
  assign _zz_7468 = _zz_7469[35 : 0];
  assign _zz_7469 = _zz_7470;
  assign _zz_7470 = ($signed(_zz_7471) >>> _zz_655);
  assign _zz_7471 = _zz_7472;
  assign _zz_7472 = ($signed(_zz_7474) + $signed(_zz_651));
  assign _zz_7473 = ({9'd0,data_mid_4_2_real} <<< 9);
  assign _zz_7474 = {{9{_zz_7473[26]}}, _zz_7473};
  assign _zz_7475 = fixTo_784_dout;
  assign _zz_7476 = _zz_7477[35 : 0];
  assign _zz_7477 = _zz_7478;
  assign _zz_7478 = ($signed(_zz_7479) >>> _zz_655);
  assign _zz_7479 = _zz_7480;
  assign _zz_7480 = ($signed(_zz_7482) + $signed(_zz_652));
  assign _zz_7481 = ({9'd0,data_mid_4_2_imag} <<< 9);
  assign _zz_7482 = {{9{_zz_7481[26]}}, _zz_7481};
  assign _zz_7483 = fixTo_785_dout;
  assign _zz_7484 = ($signed(twiddle_factor_table_18_real) + $signed(twiddle_factor_table_18_imag));
  assign _zz_7485 = ($signed(_zz_658) - $signed(_zz_7486));
  assign _zz_7486 = ($signed(_zz_7487) * $signed(twiddle_factor_table_18_imag));
  assign _zz_7487 = ($signed(data_mid_4_19_real) + $signed(data_mid_4_19_imag));
  assign _zz_7488 = fixTo_786_dout;
  assign _zz_7489 = ($signed(_zz_658) + $signed(_zz_7490));
  assign _zz_7490 = ($signed(_zz_7491) * $signed(twiddle_factor_table_18_real));
  assign _zz_7491 = ($signed(data_mid_4_19_imag) - $signed(data_mid_4_19_real));
  assign _zz_7492 = fixTo_787_dout;
  assign _zz_7493 = _zz_7494[35 : 0];
  assign _zz_7494 = _zz_7495;
  assign _zz_7495 = ($signed(_zz_7496) >>> _zz_659);
  assign _zz_7496 = _zz_7497;
  assign _zz_7497 = ($signed(_zz_7499) - $signed(_zz_656));
  assign _zz_7498 = ({9'd0,data_mid_4_3_real} <<< 9);
  assign _zz_7499 = {{9{_zz_7498[26]}}, _zz_7498};
  assign _zz_7500 = fixTo_788_dout;
  assign _zz_7501 = _zz_7502[35 : 0];
  assign _zz_7502 = _zz_7503;
  assign _zz_7503 = ($signed(_zz_7504) >>> _zz_659);
  assign _zz_7504 = _zz_7505;
  assign _zz_7505 = ($signed(_zz_7507) - $signed(_zz_657));
  assign _zz_7506 = ({9'd0,data_mid_4_3_imag} <<< 9);
  assign _zz_7507 = {{9{_zz_7506[26]}}, _zz_7506};
  assign _zz_7508 = fixTo_789_dout;
  assign _zz_7509 = _zz_7510[35 : 0];
  assign _zz_7510 = _zz_7511;
  assign _zz_7511 = ($signed(_zz_7512) >>> _zz_660);
  assign _zz_7512 = _zz_7513;
  assign _zz_7513 = ($signed(_zz_7515) + $signed(_zz_656));
  assign _zz_7514 = ({9'd0,data_mid_4_3_real} <<< 9);
  assign _zz_7515 = {{9{_zz_7514[26]}}, _zz_7514};
  assign _zz_7516 = fixTo_790_dout;
  assign _zz_7517 = _zz_7518[35 : 0];
  assign _zz_7518 = _zz_7519;
  assign _zz_7519 = ($signed(_zz_7520) >>> _zz_660);
  assign _zz_7520 = _zz_7521;
  assign _zz_7521 = ($signed(_zz_7523) + $signed(_zz_657));
  assign _zz_7522 = ({9'd0,data_mid_4_3_imag} <<< 9);
  assign _zz_7523 = {{9{_zz_7522[26]}}, _zz_7522};
  assign _zz_7524 = fixTo_791_dout;
  assign _zz_7525 = ($signed(twiddle_factor_table_19_real) + $signed(twiddle_factor_table_19_imag));
  assign _zz_7526 = ($signed(_zz_663) - $signed(_zz_7527));
  assign _zz_7527 = ($signed(_zz_7528) * $signed(twiddle_factor_table_19_imag));
  assign _zz_7528 = ($signed(data_mid_4_20_real) + $signed(data_mid_4_20_imag));
  assign _zz_7529 = fixTo_792_dout;
  assign _zz_7530 = ($signed(_zz_663) + $signed(_zz_7531));
  assign _zz_7531 = ($signed(_zz_7532) * $signed(twiddle_factor_table_19_real));
  assign _zz_7532 = ($signed(data_mid_4_20_imag) - $signed(data_mid_4_20_real));
  assign _zz_7533 = fixTo_793_dout;
  assign _zz_7534 = _zz_7535[35 : 0];
  assign _zz_7535 = _zz_7536;
  assign _zz_7536 = ($signed(_zz_7537) >>> _zz_664);
  assign _zz_7537 = _zz_7538;
  assign _zz_7538 = ($signed(_zz_7540) - $signed(_zz_661));
  assign _zz_7539 = ({9'd0,data_mid_4_4_real} <<< 9);
  assign _zz_7540 = {{9{_zz_7539[26]}}, _zz_7539};
  assign _zz_7541 = fixTo_794_dout;
  assign _zz_7542 = _zz_7543[35 : 0];
  assign _zz_7543 = _zz_7544;
  assign _zz_7544 = ($signed(_zz_7545) >>> _zz_664);
  assign _zz_7545 = _zz_7546;
  assign _zz_7546 = ($signed(_zz_7548) - $signed(_zz_662));
  assign _zz_7547 = ({9'd0,data_mid_4_4_imag} <<< 9);
  assign _zz_7548 = {{9{_zz_7547[26]}}, _zz_7547};
  assign _zz_7549 = fixTo_795_dout;
  assign _zz_7550 = _zz_7551[35 : 0];
  assign _zz_7551 = _zz_7552;
  assign _zz_7552 = ($signed(_zz_7553) >>> _zz_665);
  assign _zz_7553 = _zz_7554;
  assign _zz_7554 = ($signed(_zz_7556) + $signed(_zz_661));
  assign _zz_7555 = ({9'd0,data_mid_4_4_real} <<< 9);
  assign _zz_7556 = {{9{_zz_7555[26]}}, _zz_7555};
  assign _zz_7557 = fixTo_796_dout;
  assign _zz_7558 = _zz_7559[35 : 0];
  assign _zz_7559 = _zz_7560;
  assign _zz_7560 = ($signed(_zz_7561) >>> _zz_665);
  assign _zz_7561 = _zz_7562;
  assign _zz_7562 = ($signed(_zz_7564) + $signed(_zz_662));
  assign _zz_7563 = ({9'd0,data_mid_4_4_imag} <<< 9);
  assign _zz_7564 = {{9{_zz_7563[26]}}, _zz_7563};
  assign _zz_7565 = fixTo_797_dout;
  assign _zz_7566 = ($signed(twiddle_factor_table_20_real) + $signed(twiddle_factor_table_20_imag));
  assign _zz_7567 = ($signed(_zz_668) - $signed(_zz_7568));
  assign _zz_7568 = ($signed(_zz_7569) * $signed(twiddle_factor_table_20_imag));
  assign _zz_7569 = ($signed(data_mid_4_21_real) + $signed(data_mid_4_21_imag));
  assign _zz_7570 = fixTo_798_dout;
  assign _zz_7571 = ($signed(_zz_668) + $signed(_zz_7572));
  assign _zz_7572 = ($signed(_zz_7573) * $signed(twiddle_factor_table_20_real));
  assign _zz_7573 = ($signed(data_mid_4_21_imag) - $signed(data_mid_4_21_real));
  assign _zz_7574 = fixTo_799_dout;
  assign _zz_7575 = _zz_7576[35 : 0];
  assign _zz_7576 = _zz_7577;
  assign _zz_7577 = ($signed(_zz_7578) >>> _zz_669);
  assign _zz_7578 = _zz_7579;
  assign _zz_7579 = ($signed(_zz_7581) - $signed(_zz_666));
  assign _zz_7580 = ({9'd0,data_mid_4_5_real} <<< 9);
  assign _zz_7581 = {{9{_zz_7580[26]}}, _zz_7580};
  assign _zz_7582 = fixTo_800_dout;
  assign _zz_7583 = _zz_7584[35 : 0];
  assign _zz_7584 = _zz_7585;
  assign _zz_7585 = ($signed(_zz_7586) >>> _zz_669);
  assign _zz_7586 = _zz_7587;
  assign _zz_7587 = ($signed(_zz_7589) - $signed(_zz_667));
  assign _zz_7588 = ({9'd0,data_mid_4_5_imag} <<< 9);
  assign _zz_7589 = {{9{_zz_7588[26]}}, _zz_7588};
  assign _zz_7590 = fixTo_801_dout;
  assign _zz_7591 = _zz_7592[35 : 0];
  assign _zz_7592 = _zz_7593;
  assign _zz_7593 = ($signed(_zz_7594) >>> _zz_670);
  assign _zz_7594 = _zz_7595;
  assign _zz_7595 = ($signed(_zz_7597) + $signed(_zz_666));
  assign _zz_7596 = ({9'd0,data_mid_4_5_real} <<< 9);
  assign _zz_7597 = {{9{_zz_7596[26]}}, _zz_7596};
  assign _zz_7598 = fixTo_802_dout;
  assign _zz_7599 = _zz_7600[35 : 0];
  assign _zz_7600 = _zz_7601;
  assign _zz_7601 = ($signed(_zz_7602) >>> _zz_670);
  assign _zz_7602 = _zz_7603;
  assign _zz_7603 = ($signed(_zz_7605) + $signed(_zz_667));
  assign _zz_7604 = ({9'd0,data_mid_4_5_imag} <<< 9);
  assign _zz_7605 = {{9{_zz_7604[26]}}, _zz_7604};
  assign _zz_7606 = fixTo_803_dout;
  assign _zz_7607 = ($signed(twiddle_factor_table_21_real) + $signed(twiddle_factor_table_21_imag));
  assign _zz_7608 = ($signed(_zz_673) - $signed(_zz_7609));
  assign _zz_7609 = ($signed(_zz_7610) * $signed(twiddle_factor_table_21_imag));
  assign _zz_7610 = ($signed(data_mid_4_22_real) + $signed(data_mid_4_22_imag));
  assign _zz_7611 = fixTo_804_dout;
  assign _zz_7612 = ($signed(_zz_673) + $signed(_zz_7613));
  assign _zz_7613 = ($signed(_zz_7614) * $signed(twiddle_factor_table_21_real));
  assign _zz_7614 = ($signed(data_mid_4_22_imag) - $signed(data_mid_4_22_real));
  assign _zz_7615 = fixTo_805_dout;
  assign _zz_7616 = _zz_7617[35 : 0];
  assign _zz_7617 = _zz_7618;
  assign _zz_7618 = ($signed(_zz_7619) >>> _zz_674);
  assign _zz_7619 = _zz_7620;
  assign _zz_7620 = ($signed(_zz_7622) - $signed(_zz_671));
  assign _zz_7621 = ({9'd0,data_mid_4_6_real} <<< 9);
  assign _zz_7622 = {{9{_zz_7621[26]}}, _zz_7621};
  assign _zz_7623 = fixTo_806_dout;
  assign _zz_7624 = _zz_7625[35 : 0];
  assign _zz_7625 = _zz_7626;
  assign _zz_7626 = ($signed(_zz_7627) >>> _zz_674);
  assign _zz_7627 = _zz_7628;
  assign _zz_7628 = ($signed(_zz_7630) - $signed(_zz_672));
  assign _zz_7629 = ({9'd0,data_mid_4_6_imag} <<< 9);
  assign _zz_7630 = {{9{_zz_7629[26]}}, _zz_7629};
  assign _zz_7631 = fixTo_807_dout;
  assign _zz_7632 = _zz_7633[35 : 0];
  assign _zz_7633 = _zz_7634;
  assign _zz_7634 = ($signed(_zz_7635) >>> _zz_675);
  assign _zz_7635 = _zz_7636;
  assign _zz_7636 = ($signed(_zz_7638) + $signed(_zz_671));
  assign _zz_7637 = ({9'd0,data_mid_4_6_real} <<< 9);
  assign _zz_7638 = {{9{_zz_7637[26]}}, _zz_7637};
  assign _zz_7639 = fixTo_808_dout;
  assign _zz_7640 = _zz_7641[35 : 0];
  assign _zz_7641 = _zz_7642;
  assign _zz_7642 = ($signed(_zz_7643) >>> _zz_675);
  assign _zz_7643 = _zz_7644;
  assign _zz_7644 = ($signed(_zz_7646) + $signed(_zz_672));
  assign _zz_7645 = ({9'd0,data_mid_4_6_imag} <<< 9);
  assign _zz_7646 = {{9{_zz_7645[26]}}, _zz_7645};
  assign _zz_7647 = fixTo_809_dout;
  assign _zz_7648 = ($signed(twiddle_factor_table_22_real) + $signed(twiddle_factor_table_22_imag));
  assign _zz_7649 = ($signed(_zz_678) - $signed(_zz_7650));
  assign _zz_7650 = ($signed(_zz_7651) * $signed(twiddle_factor_table_22_imag));
  assign _zz_7651 = ($signed(data_mid_4_23_real) + $signed(data_mid_4_23_imag));
  assign _zz_7652 = fixTo_810_dout;
  assign _zz_7653 = ($signed(_zz_678) + $signed(_zz_7654));
  assign _zz_7654 = ($signed(_zz_7655) * $signed(twiddle_factor_table_22_real));
  assign _zz_7655 = ($signed(data_mid_4_23_imag) - $signed(data_mid_4_23_real));
  assign _zz_7656 = fixTo_811_dout;
  assign _zz_7657 = _zz_7658[35 : 0];
  assign _zz_7658 = _zz_7659;
  assign _zz_7659 = ($signed(_zz_7660) >>> _zz_679);
  assign _zz_7660 = _zz_7661;
  assign _zz_7661 = ($signed(_zz_7663) - $signed(_zz_676));
  assign _zz_7662 = ({9'd0,data_mid_4_7_real} <<< 9);
  assign _zz_7663 = {{9{_zz_7662[26]}}, _zz_7662};
  assign _zz_7664 = fixTo_812_dout;
  assign _zz_7665 = _zz_7666[35 : 0];
  assign _zz_7666 = _zz_7667;
  assign _zz_7667 = ($signed(_zz_7668) >>> _zz_679);
  assign _zz_7668 = _zz_7669;
  assign _zz_7669 = ($signed(_zz_7671) - $signed(_zz_677));
  assign _zz_7670 = ({9'd0,data_mid_4_7_imag} <<< 9);
  assign _zz_7671 = {{9{_zz_7670[26]}}, _zz_7670};
  assign _zz_7672 = fixTo_813_dout;
  assign _zz_7673 = _zz_7674[35 : 0];
  assign _zz_7674 = _zz_7675;
  assign _zz_7675 = ($signed(_zz_7676) >>> _zz_680);
  assign _zz_7676 = _zz_7677;
  assign _zz_7677 = ($signed(_zz_7679) + $signed(_zz_676));
  assign _zz_7678 = ({9'd0,data_mid_4_7_real} <<< 9);
  assign _zz_7679 = {{9{_zz_7678[26]}}, _zz_7678};
  assign _zz_7680 = fixTo_814_dout;
  assign _zz_7681 = _zz_7682[35 : 0];
  assign _zz_7682 = _zz_7683;
  assign _zz_7683 = ($signed(_zz_7684) >>> _zz_680);
  assign _zz_7684 = _zz_7685;
  assign _zz_7685 = ($signed(_zz_7687) + $signed(_zz_677));
  assign _zz_7686 = ({9'd0,data_mid_4_7_imag} <<< 9);
  assign _zz_7687 = {{9{_zz_7686[26]}}, _zz_7686};
  assign _zz_7688 = fixTo_815_dout;
  assign _zz_7689 = ($signed(twiddle_factor_table_23_real) + $signed(twiddle_factor_table_23_imag));
  assign _zz_7690 = ($signed(_zz_683) - $signed(_zz_7691));
  assign _zz_7691 = ($signed(_zz_7692) * $signed(twiddle_factor_table_23_imag));
  assign _zz_7692 = ($signed(data_mid_4_24_real) + $signed(data_mid_4_24_imag));
  assign _zz_7693 = fixTo_816_dout;
  assign _zz_7694 = ($signed(_zz_683) + $signed(_zz_7695));
  assign _zz_7695 = ($signed(_zz_7696) * $signed(twiddle_factor_table_23_real));
  assign _zz_7696 = ($signed(data_mid_4_24_imag) - $signed(data_mid_4_24_real));
  assign _zz_7697 = fixTo_817_dout;
  assign _zz_7698 = _zz_7699[35 : 0];
  assign _zz_7699 = _zz_7700;
  assign _zz_7700 = ($signed(_zz_7701) >>> _zz_684);
  assign _zz_7701 = _zz_7702;
  assign _zz_7702 = ($signed(_zz_7704) - $signed(_zz_681));
  assign _zz_7703 = ({9'd0,data_mid_4_8_real} <<< 9);
  assign _zz_7704 = {{9{_zz_7703[26]}}, _zz_7703};
  assign _zz_7705 = fixTo_818_dout;
  assign _zz_7706 = _zz_7707[35 : 0];
  assign _zz_7707 = _zz_7708;
  assign _zz_7708 = ($signed(_zz_7709) >>> _zz_684);
  assign _zz_7709 = _zz_7710;
  assign _zz_7710 = ($signed(_zz_7712) - $signed(_zz_682));
  assign _zz_7711 = ({9'd0,data_mid_4_8_imag} <<< 9);
  assign _zz_7712 = {{9{_zz_7711[26]}}, _zz_7711};
  assign _zz_7713 = fixTo_819_dout;
  assign _zz_7714 = _zz_7715[35 : 0];
  assign _zz_7715 = _zz_7716;
  assign _zz_7716 = ($signed(_zz_7717) >>> _zz_685);
  assign _zz_7717 = _zz_7718;
  assign _zz_7718 = ($signed(_zz_7720) + $signed(_zz_681));
  assign _zz_7719 = ({9'd0,data_mid_4_8_real} <<< 9);
  assign _zz_7720 = {{9{_zz_7719[26]}}, _zz_7719};
  assign _zz_7721 = fixTo_820_dout;
  assign _zz_7722 = _zz_7723[35 : 0];
  assign _zz_7723 = _zz_7724;
  assign _zz_7724 = ($signed(_zz_7725) >>> _zz_685);
  assign _zz_7725 = _zz_7726;
  assign _zz_7726 = ($signed(_zz_7728) + $signed(_zz_682));
  assign _zz_7727 = ({9'd0,data_mid_4_8_imag} <<< 9);
  assign _zz_7728 = {{9{_zz_7727[26]}}, _zz_7727};
  assign _zz_7729 = fixTo_821_dout;
  assign _zz_7730 = ($signed(twiddle_factor_table_24_real) + $signed(twiddle_factor_table_24_imag));
  assign _zz_7731 = ($signed(_zz_688) - $signed(_zz_7732));
  assign _zz_7732 = ($signed(_zz_7733) * $signed(twiddle_factor_table_24_imag));
  assign _zz_7733 = ($signed(data_mid_4_25_real) + $signed(data_mid_4_25_imag));
  assign _zz_7734 = fixTo_822_dout;
  assign _zz_7735 = ($signed(_zz_688) + $signed(_zz_7736));
  assign _zz_7736 = ($signed(_zz_7737) * $signed(twiddle_factor_table_24_real));
  assign _zz_7737 = ($signed(data_mid_4_25_imag) - $signed(data_mid_4_25_real));
  assign _zz_7738 = fixTo_823_dout;
  assign _zz_7739 = _zz_7740[35 : 0];
  assign _zz_7740 = _zz_7741;
  assign _zz_7741 = ($signed(_zz_7742) >>> _zz_689);
  assign _zz_7742 = _zz_7743;
  assign _zz_7743 = ($signed(_zz_7745) - $signed(_zz_686));
  assign _zz_7744 = ({9'd0,data_mid_4_9_real} <<< 9);
  assign _zz_7745 = {{9{_zz_7744[26]}}, _zz_7744};
  assign _zz_7746 = fixTo_824_dout;
  assign _zz_7747 = _zz_7748[35 : 0];
  assign _zz_7748 = _zz_7749;
  assign _zz_7749 = ($signed(_zz_7750) >>> _zz_689);
  assign _zz_7750 = _zz_7751;
  assign _zz_7751 = ($signed(_zz_7753) - $signed(_zz_687));
  assign _zz_7752 = ({9'd0,data_mid_4_9_imag} <<< 9);
  assign _zz_7753 = {{9{_zz_7752[26]}}, _zz_7752};
  assign _zz_7754 = fixTo_825_dout;
  assign _zz_7755 = _zz_7756[35 : 0];
  assign _zz_7756 = _zz_7757;
  assign _zz_7757 = ($signed(_zz_7758) >>> _zz_690);
  assign _zz_7758 = _zz_7759;
  assign _zz_7759 = ($signed(_zz_7761) + $signed(_zz_686));
  assign _zz_7760 = ({9'd0,data_mid_4_9_real} <<< 9);
  assign _zz_7761 = {{9{_zz_7760[26]}}, _zz_7760};
  assign _zz_7762 = fixTo_826_dout;
  assign _zz_7763 = _zz_7764[35 : 0];
  assign _zz_7764 = _zz_7765;
  assign _zz_7765 = ($signed(_zz_7766) >>> _zz_690);
  assign _zz_7766 = _zz_7767;
  assign _zz_7767 = ($signed(_zz_7769) + $signed(_zz_687));
  assign _zz_7768 = ({9'd0,data_mid_4_9_imag} <<< 9);
  assign _zz_7769 = {{9{_zz_7768[26]}}, _zz_7768};
  assign _zz_7770 = fixTo_827_dout;
  assign _zz_7771 = ($signed(twiddle_factor_table_25_real) + $signed(twiddle_factor_table_25_imag));
  assign _zz_7772 = ($signed(_zz_693) - $signed(_zz_7773));
  assign _zz_7773 = ($signed(_zz_7774) * $signed(twiddle_factor_table_25_imag));
  assign _zz_7774 = ($signed(data_mid_4_26_real) + $signed(data_mid_4_26_imag));
  assign _zz_7775 = fixTo_828_dout;
  assign _zz_7776 = ($signed(_zz_693) + $signed(_zz_7777));
  assign _zz_7777 = ($signed(_zz_7778) * $signed(twiddle_factor_table_25_real));
  assign _zz_7778 = ($signed(data_mid_4_26_imag) - $signed(data_mid_4_26_real));
  assign _zz_7779 = fixTo_829_dout;
  assign _zz_7780 = _zz_7781[35 : 0];
  assign _zz_7781 = _zz_7782;
  assign _zz_7782 = ($signed(_zz_7783) >>> _zz_694);
  assign _zz_7783 = _zz_7784;
  assign _zz_7784 = ($signed(_zz_7786) - $signed(_zz_691));
  assign _zz_7785 = ({9'd0,data_mid_4_10_real} <<< 9);
  assign _zz_7786 = {{9{_zz_7785[26]}}, _zz_7785};
  assign _zz_7787 = fixTo_830_dout;
  assign _zz_7788 = _zz_7789[35 : 0];
  assign _zz_7789 = _zz_7790;
  assign _zz_7790 = ($signed(_zz_7791) >>> _zz_694);
  assign _zz_7791 = _zz_7792;
  assign _zz_7792 = ($signed(_zz_7794) - $signed(_zz_692));
  assign _zz_7793 = ({9'd0,data_mid_4_10_imag} <<< 9);
  assign _zz_7794 = {{9{_zz_7793[26]}}, _zz_7793};
  assign _zz_7795 = fixTo_831_dout;
  assign _zz_7796 = _zz_7797[35 : 0];
  assign _zz_7797 = _zz_7798;
  assign _zz_7798 = ($signed(_zz_7799) >>> _zz_695);
  assign _zz_7799 = _zz_7800;
  assign _zz_7800 = ($signed(_zz_7802) + $signed(_zz_691));
  assign _zz_7801 = ({9'd0,data_mid_4_10_real} <<< 9);
  assign _zz_7802 = {{9{_zz_7801[26]}}, _zz_7801};
  assign _zz_7803 = fixTo_832_dout;
  assign _zz_7804 = _zz_7805[35 : 0];
  assign _zz_7805 = _zz_7806;
  assign _zz_7806 = ($signed(_zz_7807) >>> _zz_695);
  assign _zz_7807 = _zz_7808;
  assign _zz_7808 = ($signed(_zz_7810) + $signed(_zz_692));
  assign _zz_7809 = ({9'd0,data_mid_4_10_imag} <<< 9);
  assign _zz_7810 = {{9{_zz_7809[26]}}, _zz_7809};
  assign _zz_7811 = fixTo_833_dout;
  assign _zz_7812 = ($signed(twiddle_factor_table_26_real) + $signed(twiddle_factor_table_26_imag));
  assign _zz_7813 = ($signed(_zz_698) - $signed(_zz_7814));
  assign _zz_7814 = ($signed(_zz_7815) * $signed(twiddle_factor_table_26_imag));
  assign _zz_7815 = ($signed(data_mid_4_27_real) + $signed(data_mid_4_27_imag));
  assign _zz_7816 = fixTo_834_dout;
  assign _zz_7817 = ($signed(_zz_698) + $signed(_zz_7818));
  assign _zz_7818 = ($signed(_zz_7819) * $signed(twiddle_factor_table_26_real));
  assign _zz_7819 = ($signed(data_mid_4_27_imag) - $signed(data_mid_4_27_real));
  assign _zz_7820 = fixTo_835_dout;
  assign _zz_7821 = _zz_7822[35 : 0];
  assign _zz_7822 = _zz_7823;
  assign _zz_7823 = ($signed(_zz_7824) >>> _zz_699);
  assign _zz_7824 = _zz_7825;
  assign _zz_7825 = ($signed(_zz_7827) - $signed(_zz_696));
  assign _zz_7826 = ({9'd0,data_mid_4_11_real} <<< 9);
  assign _zz_7827 = {{9{_zz_7826[26]}}, _zz_7826};
  assign _zz_7828 = fixTo_836_dout;
  assign _zz_7829 = _zz_7830[35 : 0];
  assign _zz_7830 = _zz_7831;
  assign _zz_7831 = ($signed(_zz_7832) >>> _zz_699);
  assign _zz_7832 = _zz_7833;
  assign _zz_7833 = ($signed(_zz_7835) - $signed(_zz_697));
  assign _zz_7834 = ({9'd0,data_mid_4_11_imag} <<< 9);
  assign _zz_7835 = {{9{_zz_7834[26]}}, _zz_7834};
  assign _zz_7836 = fixTo_837_dout;
  assign _zz_7837 = _zz_7838[35 : 0];
  assign _zz_7838 = _zz_7839;
  assign _zz_7839 = ($signed(_zz_7840) >>> _zz_700);
  assign _zz_7840 = _zz_7841;
  assign _zz_7841 = ($signed(_zz_7843) + $signed(_zz_696));
  assign _zz_7842 = ({9'd0,data_mid_4_11_real} <<< 9);
  assign _zz_7843 = {{9{_zz_7842[26]}}, _zz_7842};
  assign _zz_7844 = fixTo_838_dout;
  assign _zz_7845 = _zz_7846[35 : 0];
  assign _zz_7846 = _zz_7847;
  assign _zz_7847 = ($signed(_zz_7848) >>> _zz_700);
  assign _zz_7848 = _zz_7849;
  assign _zz_7849 = ($signed(_zz_7851) + $signed(_zz_697));
  assign _zz_7850 = ({9'd0,data_mid_4_11_imag} <<< 9);
  assign _zz_7851 = {{9{_zz_7850[26]}}, _zz_7850};
  assign _zz_7852 = fixTo_839_dout;
  assign _zz_7853 = ($signed(twiddle_factor_table_27_real) + $signed(twiddle_factor_table_27_imag));
  assign _zz_7854 = ($signed(_zz_703) - $signed(_zz_7855));
  assign _zz_7855 = ($signed(_zz_7856) * $signed(twiddle_factor_table_27_imag));
  assign _zz_7856 = ($signed(data_mid_4_28_real) + $signed(data_mid_4_28_imag));
  assign _zz_7857 = fixTo_840_dout;
  assign _zz_7858 = ($signed(_zz_703) + $signed(_zz_7859));
  assign _zz_7859 = ($signed(_zz_7860) * $signed(twiddle_factor_table_27_real));
  assign _zz_7860 = ($signed(data_mid_4_28_imag) - $signed(data_mid_4_28_real));
  assign _zz_7861 = fixTo_841_dout;
  assign _zz_7862 = _zz_7863[35 : 0];
  assign _zz_7863 = _zz_7864;
  assign _zz_7864 = ($signed(_zz_7865) >>> _zz_704);
  assign _zz_7865 = _zz_7866;
  assign _zz_7866 = ($signed(_zz_7868) - $signed(_zz_701));
  assign _zz_7867 = ({9'd0,data_mid_4_12_real} <<< 9);
  assign _zz_7868 = {{9{_zz_7867[26]}}, _zz_7867};
  assign _zz_7869 = fixTo_842_dout;
  assign _zz_7870 = _zz_7871[35 : 0];
  assign _zz_7871 = _zz_7872;
  assign _zz_7872 = ($signed(_zz_7873) >>> _zz_704);
  assign _zz_7873 = _zz_7874;
  assign _zz_7874 = ($signed(_zz_7876) - $signed(_zz_702));
  assign _zz_7875 = ({9'd0,data_mid_4_12_imag} <<< 9);
  assign _zz_7876 = {{9{_zz_7875[26]}}, _zz_7875};
  assign _zz_7877 = fixTo_843_dout;
  assign _zz_7878 = _zz_7879[35 : 0];
  assign _zz_7879 = _zz_7880;
  assign _zz_7880 = ($signed(_zz_7881) >>> _zz_705);
  assign _zz_7881 = _zz_7882;
  assign _zz_7882 = ($signed(_zz_7884) + $signed(_zz_701));
  assign _zz_7883 = ({9'd0,data_mid_4_12_real} <<< 9);
  assign _zz_7884 = {{9{_zz_7883[26]}}, _zz_7883};
  assign _zz_7885 = fixTo_844_dout;
  assign _zz_7886 = _zz_7887[35 : 0];
  assign _zz_7887 = _zz_7888;
  assign _zz_7888 = ($signed(_zz_7889) >>> _zz_705);
  assign _zz_7889 = _zz_7890;
  assign _zz_7890 = ($signed(_zz_7892) + $signed(_zz_702));
  assign _zz_7891 = ({9'd0,data_mid_4_12_imag} <<< 9);
  assign _zz_7892 = {{9{_zz_7891[26]}}, _zz_7891};
  assign _zz_7893 = fixTo_845_dout;
  assign _zz_7894 = ($signed(twiddle_factor_table_28_real) + $signed(twiddle_factor_table_28_imag));
  assign _zz_7895 = ($signed(_zz_708) - $signed(_zz_7896));
  assign _zz_7896 = ($signed(_zz_7897) * $signed(twiddle_factor_table_28_imag));
  assign _zz_7897 = ($signed(data_mid_4_29_real) + $signed(data_mid_4_29_imag));
  assign _zz_7898 = fixTo_846_dout;
  assign _zz_7899 = ($signed(_zz_708) + $signed(_zz_7900));
  assign _zz_7900 = ($signed(_zz_7901) * $signed(twiddle_factor_table_28_real));
  assign _zz_7901 = ($signed(data_mid_4_29_imag) - $signed(data_mid_4_29_real));
  assign _zz_7902 = fixTo_847_dout;
  assign _zz_7903 = _zz_7904[35 : 0];
  assign _zz_7904 = _zz_7905;
  assign _zz_7905 = ($signed(_zz_7906) >>> _zz_709);
  assign _zz_7906 = _zz_7907;
  assign _zz_7907 = ($signed(_zz_7909) - $signed(_zz_706));
  assign _zz_7908 = ({9'd0,data_mid_4_13_real} <<< 9);
  assign _zz_7909 = {{9{_zz_7908[26]}}, _zz_7908};
  assign _zz_7910 = fixTo_848_dout;
  assign _zz_7911 = _zz_7912[35 : 0];
  assign _zz_7912 = _zz_7913;
  assign _zz_7913 = ($signed(_zz_7914) >>> _zz_709);
  assign _zz_7914 = _zz_7915;
  assign _zz_7915 = ($signed(_zz_7917) - $signed(_zz_707));
  assign _zz_7916 = ({9'd0,data_mid_4_13_imag} <<< 9);
  assign _zz_7917 = {{9{_zz_7916[26]}}, _zz_7916};
  assign _zz_7918 = fixTo_849_dout;
  assign _zz_7919 = _zz_7920[35 : 0];
  assign _zz_7920 = _zz_7921;
  assign _zz_7921 = ($signed(_zz_7922) >>> _zz_710);
  assign _zz_7922 = _zz_7923;
  assign _zz_7923 = ($signed(_zz_7925) + $signed(_zz_706));
  assign _zz_7924 = ({9'd0,data_mid_4_13_real} <<< 9);
  assign _zz_7925 = {{9{_zz_7924[26]}}, _zz_7924};
  assign _zz_7926 = fixTo_850_dout;
  assign _zz_7927 = _zz_7928[35 : 0];
  assign _zz_7928 = _zz_7929;
  assign _zz_7929 = ($signed(_zz_7930) >>> _zz_710);
  assign _zz_7930 = _zz_7931;
  assign _zz_7931 = ($signed(_zz_7933) + $signed(_zz_707));
  assign _zz_7932 = ({9'd0,data_mid_4_13_imag} <<< 9);
  assign _zz_7933 = {{9{_zz_7932[26]}}, _zz_7932};
  assign _zz_7934 = fixTo_851_dout;
  assign _zz_7935 = ($signed(twiddle_factor_table_29_real) + $signed(twiddle_factor_table_29_imag));
  assign _zz_7936 = ($signed(_zz_713) - $signed(_zz_7937));
  assign _zz_7937 = ($signed(_zz_7938) * $signed(twiddle_factor_table_29_imag));
  assign _zz_7938 = ($signed(data_mid_4_30_real) + $signed(data_mid_4_30_imag));
  assign _zz_7939 = fixTo_852_dout;
  assign _zz_7940 = ($signed(_zz_713) + $signed(_zz_7941));
  assign _zz_7941 = ($signed(_zz_7942) * $signed(twiddle_factor_table_29_real));
  assign _zz_7942 = ($signed(data_mid_4_30_imag) - $signed(data_mid_4_30_real));
  assign _zz_7943 = fixTo_853_dout;
  assign _zz_7944 = _zz_7945[35 : 0];
  assign _zz_7945 = _zz_7946;
  assign _zz_7946 = ($signed(_zz_7947) >>> _zz_714);
  assign _zz_7947 = _zz_7948;
  assign _zz_7948 = ($signed(_zz_7950) - $signed(_zz_711));
  assign _zz_7949 = ({9'd0,data_mid_4_14_real} <<< 9);
  assign _zz_7950 = {{9{_zz_7949[26]}}, _zz_7949};
  assign _zz_7951 = fixTo_854_dout;
  assign _zz_7952 = _zz_7953[35 : 0];
  assign _zz_7953 = _zz_7954;
  assign _zz_7954 = ($signed(_zz_7955) >>> _zz_714);
  assign _zz_7955 = _zz_7956;
  assign _zz_7956 = ($signed(_zz_7958) - $signed(_zz_712));
  assign _zz_7957 = ({9'd0,data_mid_4_14_imag} <<< 9);
  assign _zz_7958 = {{9{_zz_7957[26]}}, _zz_7957};
  assign _zz_7959 = fixTo_855_dout;
  assign _zz_7960 = _zz_7961[35 : 0];
  assign _zz_7961 = _zz_7962;
  assign _zz_7962 = ($signed(_zz_7963) >>> _zz_715);
  assign _zz_7963 = _zz_7964;
  assign _zz_7964 = ($signed(_zz_7966) + $signed(_zz_711));
  assign _zz_7965 = ({9'd0,data_mid_4_14_real} <<< 9);
  assign _zz_7966 = {{9{_zz_7965[26]}}, _zz_7965};
  assign _zz_7967 = fixTo_856_dout;
  assign _zz_7968 = _zz_7969[35 : 0];
  assign _zz_7969 = _zz_7970;
  assign _zz_7970 = ($signed(_zz_7971) >>> _zz_715);
  assign _zz_7971 = _zz_7972;
  assign _zz_7972 = ($signed(_zz_7974) + $signed(_zz_712));
  assign _zz_7973 = ({9'd0,data_mid_4_14_imag} <<< 9);
  assign _zz_7974 = {{9{_zz_7973[26]}}, _zz_7973};
  assign _zz_7975 = fixTo_857_dout;
  assign _zz_7976 = ($signed(twiddle_factor_table_30_real) + $signed(twiddle_factor_table_30_imag));
  assign _zz_7977 = ($signed(_zz_718) - $signed(_zz_7978));
  assign _zz_7978 = ($signed(_zz_7979) * $signed(twiddle_factor_table_30_imag));
  assign _zz_7979 = ($signed(data_mid_4_31_real) + $signed(data_mid_4_31_imag));
  assign _zz_7980 = fixTo_858_dout;
  assign _zz_7981 = ($signed(_zz_718) + $signed(_zz_7982));
  assign _zz_7982 = ($signed(_zz_7983) * $signed(twiddle_factor_table_30_real));
  assign _zz_7983 = ($signed(data_mid_4_31_imag) - $signed(data_mid_4_31_real));
  assign _zz_7984 = fixTo_859_dout;
  assign _zz_7985 = _zz_7986[35 : 0];
  assign _zz_7986 = _zz_7987;
  assign _zz_7987 = ($signed(_zz_7988) >>> _zz_719);
  assign _zz_7988 = _zz_7989;
  assign _zz_7989 = ($signed(_zz_7991) - $signed(_zz_716));
  assign _zz_7990 = ({9'd0,data_mid_4_15_real} <<< 9);
  assign _zz_7991 = {{9{_zz_7990[26]}}, _zz_7990};
  assign _zz_7992 = fixTo_860_dout;
  assign _zz_7993 = _zz_7994[35 : 0];
  assign _zz_7994 = _zz_7995;
  assign _zz_7995 = ($signed(_zz_7996) >>> _zz_719);
  assign _zz_7996 = _zz_7997;
  assign _zz_7997 = ($signed(_zz_7999) - $signed(_zz_717));
  assign _zz_7998 = ({9'd0,data_mid_4_15_imag} <<< 9);
  assign _zz_7999 = {{9{_zz_7998[26]}}, _zz_7998};
  assign _zz_8000 = fixTo_861_dout;
  assign _zz_8001 = _zz_8002[35 : 0];
  assign _zz_8002 = _zz_8003;
  assign _zz_8003 = ($signed(_zz_8004) >>> _zz_720);
  assign _zz_8004 = _zz_8005;
  assign _zz_8005 = ($signed(_zz_8007) + $signed(_zz_716));
  assign _zz_8006 = ({9'd0,data_mid_4_15_real} <<< 9);
  assign _zz_8007 = {{9{_zz_8006[26]}}, _zz_8006};
  assign _zz_8008 = fixTo_862_dout;
  assign _zz_8009 = _zz_8010[35 : 0];
  assign _zz_8010 = _zz_8011;
  assign _zz_8011 = ($signed(_zz_8012) >>> _zz_720);
  assign _zz_8012 = _zz_8013;
  assign _zz_8013 = ($signed(_zz_8015) + $signed(_zz_717));
  assign _zz_8014 = ({9'd0,data_mid_4_15_imag} <<< 9);
  assign _zz_8015 = {{9{_zz_8014[26]}}, _zz_8014};
  assign _zz_8016 = fixTo_863_dout;
  assign _zz_8017 = ($signed(twiddle_factor_table_15_real) + $signed(twiddle_factor_table_15_imag));
  assign _zz_8018 = ($signed(_zz_723) - $signed(_zz_8019));
  assign _zz_8019 = ($signed(_zz_8020) * $signed(twiddle_factor_table_15_imag));
  assign _zz_8020 = ($signed(data_mid_4_48_real) + $signed(data_mid_4_48_imag));
  assign _zz_8021 = fixTo_864_dout;
  assign _zz_8022 = ($signed(_zz_723) + $signed(_zz_8023));
  assign _zz_8023 = ($signed(_zz_8024) * $signed(twiddle_factor_table_15_real));
  assign _zz_8024 = ($signed(data_mid_4_48_imag) - $signed(data_mid_4_48_real));
  assign _zz_8025 = fixTo_865_dout;
  assign _zz_8026 = _zz_8027[35 : 0];
  assign _zz_8027 = _zz_8028;
  assign _zz_8028 = ($signed(_zz_8029) >>> _zz_724);
  assign _zz_8029 = _zz_8030;
  assign _zz_8030 = ($signed(_zz_8032) - $signed(_zz_721));
  assign _zz_8031 = ({9'd0,data_mid_4_32_real} <<< 9);
  assign _zz_8032 = {{9{_zz_8031[26]}}, _zz_8031};
  assign _zz_8033 = fixTo_866_dout;
  assign _zz_8034 = _zz_8035[35 : 0];
  assign _zz_8035 = _zz_8036;
  assign _zz_8036 = ($signed(_zz_8037) >>> _zz_724);
  assign _zz_8037 = _zz_8038;
  assign _zz_8038 = ($signed(_zz_8040) - $signed(_zz_722));
  assign _zz_8039 = ({9'd0,data_mid_4_32_imag} <<< 9);
  assign _zz_8040 = {{9{_zz_8039[26]}}, _zz_8039};
  assign _zz_8041 = fixTo_867_dout;
  assign _zz_8042 = _zz_8043[35 : 0];
  assign _zz_8043 = _zz_8044;
  assign _zz_8044 = ($signed(_zz_8045) >>> _zz_725);
  assign _zz_8045 = _zz_8046;
  assign _zz_8046 = ($signed(_zz_8048) + $signed(_zz_721));
  assign _zz_8047 = ({9'd0,data_mid_4_32_real} <<< 9);
  assign _zz_8048 = {{9{_zz_8047[26]}}, _zz_8047};
  assign _zz_8049 = fixTo_868_dout;
  assign _zz_8050 = _zz_8051[35 : 0];
  assign _zz_8051 = _zz_8052;
  assign _zz_8052 = ($signed(_zz_8053) >>> _zz_725);
  assign _zz_8053 = _zz_8054;
  assign _zz_8054 = ($signed(_zz_8056) + $signed(_zz_722));
  assign _zz_8055 = ({9'd0,data_mid_4_32_imag} <<< 9);
  assign _zz_8056 = {{9{_zz_8055[26]}}, _zz_8055};
  assign _zz_8057 = fixTo_869_dout;
  assign _zz_8058 = ($signed(twiddle_factor_table_16_real) + $signed(twiddle_factor_table_16_imag));
  assign _zz_8059 = ($signed(_zz_728) - $signed(_zz_8060));
  assign _zz_8060 = ($signed(_zz_8061) * $signed(twiddle_factor_table_16_imag));
  assign _zz_8061 = ($signed(data_mid_4_49_real) + $signed(data_mid_4_49_imag));
  assign _zz_8062 = fixTo_870_dout;
  assign _zz_8063 = ($signed(_zz_728) + $signed(_zz_8064));
  assign _zz_8064 = ($signed(_zz_8065) * $signed(twiddle_factor_table_16_real));
  assign _zz_8065 = ($signed(data_mid_4_49_imag) - $signed(data_mid_4_49_real));
  assign _zz_8066 = fixTo_871_dout;
  assign _zz_8067 = _zz_8068[35 : 0];
  assign _zz_8068 = _zz_8069;
  assign _zz_8069 = ($signed(_zz_8070) >>> _zz_729);
  assign _zz_8070 = _zz_8071;
  assign _zz_8071 = ($signed(_zz_8073) - $signed(_zz_726));
  assign _zz_8072 = ({9'd0,data_mid_4_33_real} <<< 9);
  assign _zz_8073 = {{9{_zz_8072[26]}}, _zz_8072};
  assign _zz_8074 = fixTo_872_dout;
  assign _zz_8075 = _zz_8076[35 : 0];
  assign _zz_8076 = _zz_8077;
  assign _zz_8077 = ($signed(_zz_8078) >>> _zz_729);
  assign _zz_8078 = _zz_8079;
  assign _zz_8079 = ($signed(_zz_8081) - $signed(_zz_727));
  assign _zz_8080 = ({9'd0,data_mid_4_33_imag} <<< 9);
  assign _zz_8081 = {{9{_zz_8080[26]}}, _zz_8080};
  assign _zz_8082 = fixTo_873_dout;
  assign _zz_8083 = _zz_8084[35 : 0];
  assign _zz_8084 = _zz_8085;
  assign _zz_8085 = ($signed(_zz_8086) >>> _zz_730);
  assign _zz_8086 = _zz_8087;
  assign _zz_8087 = ($signed(_zz_8089) + $signed(_zz_726));
  assign _zz_8088 = ({9'd0,data_mid_4_33_real} <<< 9);
  assign _zz_8089 = {{9{_zz_8088[26]}}, _zz_8088};
  assign _zz_8090 = fixTo_874_dout;
  assign _zz_8091 = _zz_8092[35 : 0];
  assign _zz_8092 = _zz_8093;
  assign _zz_8093 = ($signed(_zz_8094) >>> _zz_730);
  assign _zz_8094 = _zz_8095;
  assign _zz_8095 = ($signed(_zz_8097) + $signed(_zz_727));
  assign _zz_8096 = ({9'd0,data_mid_4_33_imag} <<< 9);
  assign _zz_8097 = {{9{_zz_8096[26]}}, _zz_8096};
  assign _zz_8098 = fixTo_875_dout;
  assign _zz_8099 = ($signed(twiddle_factor_table_17_real) + $signed(twiddle_factor_table_17_imag));
  assign _zz_8100 = ($signed(_zz_733) - $signed(_zz_8101));
  assign _zz_8101 = ($signed(_zz_8102) * $signed(twiddle_factor_table_17_imag));
  assign _zz_8102 = ($signed(data_mid_4_50_real) + $signed(data_mid_4_50_imag));
  assign _zz_8103 = fixTo_876_dout;
  assign _zz_8104 = ($signed(_zz_733) + $signed(_zz_8105));
  assign _zz_8105 = ($signed(_zz_8106) * $signed(twiddle_factor_table_17_real));
  assign _zz_8106 = ($signed(data_mid_4_50_imag) - $signed(data_mid_4_50_real));
  assign _zz_8107 = fixTo_877_dout;
  assign _zz_8108 = _zz_8109[35 : 0];
  assign _zz_8109 = _zz_8110;
  assign _zz_8110 = ($signed(_zz_8111) >>> _zz_734);
  assign _zz_8111 = _zz_8112;
  assign _zz_8112 = ($signed(_zz_8114) - $signed(_zz_731));
  assign _zz_8113 = ({9'd0,data_mid_4_34_real} <<< 9);
  assign _zz_8114 = {{9{_zz_8113[26]}}, _zz_8113};
  assign _zz_8115 = fixTo_878_dout;
  assign _zz_8116 = _zz_8117[35 : 0];
  assign _zz_8117 = _zz_8118;
  assign _zz_8118 = ($signed(_zz_8119) >>> _zz_734);
  assign _zz_8119 = _zz_8120;
  assign _zz_8120 = ($signed(_zz_8122) - $signed(_zz_732));
  assign _zz_8121 = ({9'd0,data_mid_4_34_imag} <<< 9);
  assign _zz_8122 = {{9{_zz_8121[26]}}, _zz_8121};
  assign _zz_8123 = fixTo_879_dout;
  assign _zz_8124 = _zz_8125[35 : 0];
  assign _zz_8125 = _zz_8126;
  assign _zz_8126 = ($signed(_zz_8127) >>> _zz_735);
  assign _zz_8127 = _zz_8128;
  assign _zz_8128 = ($signed(_zz_8130) + $signed(_zz_731));
  assign _zz_8129 = ({9'd0,data_mid_4_34_real} <<< 9);
  assign _zz_8130 = {{9{_zz_8129[26]}}, _zz_8129};
  assign _zz_8131 = fixTo_880_dout;
  assign _zz_8132 = _zz_8133[35 : 0];
  assign _zz_8133 = _zz_8134;
  assign _zz_8134 = ($signed(_zz_8135) >>> _zz_735);
  assign _zz_8135 = _zz_8136;
  assign _zz_8136 = ($signed(_zz_8138) + $signed(_zz_732));
  assign _zz_8137 = ({9'd0,data_mid_4_34_imag} <<< 9);
  assign _zz_8138 = {{9{_zz_8137[26]}}, _zz_8137};
  assign _zz_8139 = fixTo_881_dout;
  assign _zz_8140 = ($signed(twiddle_factor_table_18_real) + $signed(twiddle_factor_table_18_imag));
  assign _zz_8141 = ($signed(_zz_738) - $signed(_zz_8142));
  assign _zz_8142 = ($signed(_zz_8143) * $signed(twiddle_factor_table_18_imag));
  assign _zz_8143 = ($signed(data_mid_4_51_real) + $signed(data_mid_4_51_imag));
  assign _zz_8144 = fixTo_882_dout;
  assign _zz_8145 = ($signed(_zz_738) + $signed(_zz_8146));
  assign _zz_8146 = ($signed(_zz_8147) * $signed(twiddle_factor_table_18_real));
  assign _zz_8147 = ($signed(data_mid_4_51_imag) - $signed(data_mid_4_51_real));
  assign _zz_8148 = fixTo_883_dout;
  assign _zz_8149 = _zz_8150[35 : 0];
  assign _zz_8150 = _zz_8151;
  assign _zz_8151 = ($signed(_zz_8152) >>> _zz_739);
  assign _zz_8152 = _zz_8153;
  assign _zz_8153 = ($signed(_zz_8155) - $signed(_zz_736));
  assign _zz_8154 = ({9'd0,data_mid_4_35_real} <<< 9);
  assign _zz_8155 = {{9{_zz_8154[26]}}, _zz_8154};
  assign _zz_8156 = fixTo_884_dout;
  assign _zz_8157 = _zz_8158[35 : 0];
  assign _zz_8158 = _zz_8159;
  assign _zz_8159 = ($signed(_zz_8160) >>> _zz_739);
  assign _zz_8160 = _zz_8161;
  assign _zz_8161 = ($signed(_zz_8163) - $signed(_zz_737));
  assign _zz_8162 = ({9'd0,data_mid_4_35_imag} <<< 9);
  assign _zz_8163 = {{9{_zz_8162[26]}}, _zz_8162};
  assign _zz_8164 = fixTo_885_dout;
  assign _zz_8165 = _zz_8166[35 : 0];
  assign _zz_8166 = _zz_8167;
  assign _zz_8167 = ($signed(_zz_8168) >>> _zz_740);
  assign _zz_8168 = _zz_8169;
  assign _zz_8169 = ($signed(_zz_8171) + $signed(_zz_736));
  assign _zz_8170 = ({9'd0,data_mid_4_35_real} <<< 9);
  assign _zz_8171 = {{9{_zz_8170[26]}}, _zz_8170};
  assign _zz_8172 = fixTo_886_dout;
  assign _zz_8173 = _zz_8174[35 : 0];
  assign _zz_8174 = _zz_8175;
  assign _zz_8175 = ($signed(_zz_8176) >>> _zz_740);
  assign _zz_8176 = _zz_8177;
  assign _zz_8177 = ($signed(_zz_8179) + $signed(_zz_737));
  assign _zz_8178 = ({9'd0,data_mid_4_35_imag} <<< 9);
  assign _zz_8179 = {{9{_zz_8178[26]}}, _zz_8178};
  assign _zz_8180 = fixTo_887_dout;
  assign _zz_8181 = ($signed(twiddle_factor_table_19_real) + $signed(twiddle_factor_table_19_imag));
  assign _zz_8182 = ($signed(_zz_743) - $signed(_zz_8183));
  assign _zz_8183 = ($signed(_zz_8184) * $signed(twiddle_factor_table_19_imag));
  assign _zz_8184 = ($signed(data_mid_4_52_real) + $signed(data_mid_4_52_imag));
  assign _zz_8185 = fixTo_888_dout;
  assign _zz_8186 = ($signed(_zz_743) + $signed(_zz_8187));
  assign _zz_8187 = ($signed(_zz_8188) * $signed(twiddle_factor_table_19_real));
  assign _zz_8188 = ($signed(data_mid_4_52_imag) - $signed(data_mid_4_52_real));
  assign _zz_8189 = fixTo_889_dout;
  assign _zz_8190 = _zz_8191[35 : 0];
  assign _zz_8191 = _zz_8192;
  assign _zz_8192 = ($signed(_zz_8193) >>> _zz_744);
  assign _zz_8193 = _zz_8194;
  assign _zz_8194 = ($signed(_zz_8196) - $signed(_zz_741));
  assign _zz_8195 = ({9'd0,data_mid_4_36_real} <<< 9);
  assign _zz_8196 = {{9{_zz_8195[26]}}, _zz_8195};
  assign _zz_8197 = fixTo_890_dout;
  assign _zz_8198 = _zz_8199[35 : 0];
  assign _zz_8199 = _zz_8200;
  assign _zz_8200 = ($signed(_zz_8201) >>> _zz_744);
  assign _zz_8201 = _zz_8202;
  assign _zz_8202 = ($signed(_zz_8204) - $signed(_zz_742));
  assign _zz_8203 = ({9'd0,data_mid_4_36_imag} <<< 9);
  assign _zz_8204 = {{9{_zz_8203[26]}}, _zz_8203};
  assign _zz_8205 = fixTo_891_dout;
  assign _zz_8206 = _zz_8207[35 : 0];
  assign _zz_8207 = _zz_8208;
  assign _zz_8208 = ($signed(_zz_8209) >>> _zz_745);
  assign _zz_8209 = _zz_8210;
  assign _zz_8210 = ($signed(_zz_8212) + $signed(_zz_741));
  assign _zz_8211 = ({9'd0,data_mid_4_36_real} <<< 9);
  assign _zz_8212 = {{9{_zz_8211[26]}}, _zz_8211};
  assign _zz_8213 = fixTo_892_dout;
  assign _zz_8214 = _zz_8215[35 : 0];
  assign _zz_8215 = _zz_8216;
  assign _zz_8216 = ($signed(_zz_8217) >>> _zz_745);
  assign _zz_8217 = _zz_8218;
  assign _zz_8218 = ($signed(_zz_8220) + $signed(_zz_742));
  assign _zz_8219 = ({9'd0,data_mid_4_36_imag} <<< 9);
  assign _zz_8220 = {{9{_zz_8219[26]}}, _zz_8219};
  assign _zz_8221 = fixTo_893_dout;
  assign _zz_8222 = ($signed(twiddle_factor_table_20_real) + $signed(twiddle_factor_table_20_imag));
  assign _zz_8223 = ($signed(_zz_748) - $signed(_zz_8224));
  assign _zz_8224 = ($signed(_zz_8225) * $signed(twiddle_factor_table_20_imag));
  assign _zz_8225 = ($signed(data_mid_4_53_real) + $signed(data_mid_4_53_imag));
  assign _zz_8226 = fixTo_894_dout;
  assign _zz_8227 = ($signed(_zz_748) + $signed(_zz_8228));
  assign _zz_8228 = ($signed(_zz_8229) * $signed(twiddle_factor_table_20_real));
  assign _zz_8229 = ($signed(data_mid_4_53_imag) - $signed(data_mid_4_53_real));
  assign _zz_8230 = fixTo_895_dout;
  assign _zz_8231 = _zz_8232[35 : 0];
  assign _zz_8232 = _zz_8233;
  assign _zz_8233 = ($signed(_zz_8234) >>> _zz_749);
  assign _zz_8234 = _zz_8235;
  assign _zz_8235 = ($signed(_zz_8237) - $signed(_zz_746));
  assign _zz_8236 = ({9'd0,data_mid_4_37_real} <<< 9);
  assign _zz_8237 = {{9{_zz_8236[26]}}, _zz_8236};
  assign _zz_8238 = fixTo_896_dout;
  assign _zz_8239 = _zz_8240[35 : 0];
  assign _zz_8240 = _zz_8241;
  assign _zz_8241 = ($signed(_zz_8242) >>> _zz_749);
  assign _zz_8242 = _zz_8243;
  assign _zz_8243 = ($signed(_zz_8245) - $signed(_zz_747));
  assign _zz_8244 = ({9'd0,data_mid_4_37_imag} <<< 9);
  assign _zz_8245 = {{9{_zz_8244[26]}}, _zz_8244};
  assign _zz_8246 = fixTo_897_dout;
  assign _zz_8247 = _zz_8248[35 : 0];
  assign _zz_8248 = _zz_8249;
  assign _zz_8249 = ($signed(_zz_8250) >>> _zz_750);
  assign _zz_8250 = _zz_8251;
  assign _zz_8251 = ($signed(_zz_8253) + $signed(_zz_746));
  assign _zz_8252 = ({9'd0,data_mid_4_37_real} <<< 9);
  assign _zz_8253 = {{9{_zz_8252[26]}}, _zz_8252};
  assign _zz_8254 = fixTo_898_dout;
  assign _zz_8255 = _zz_8256[35 : 0];
  assign _zz_8256 = _zz_8257;
  assign _zz_8257 = ($signed(_zz_8258) >>> _zz_750);
  assign _zz_8258 = _zz_8259;
  assign _zz_8259 = ($signed(_zz_8261) + $signed(_zz_747));
  assign _zz_8260 = ({9'd0,data_mid_4_37_imag} <<< 9);
  assign _zz_8261 = {{9{_zz_8260[26]}}, _zz_8260};
  assign _zz_8262 = fixTo_899_dout;
  assign _zz_8263 = ($signed(twiddle_factor_table_21_real) + $signed(twiddle_factor_table_21_imag));
  assign _zz_8264 = ($signed(_zz_753) - $signed(_zz_8265));
  assign _zz_8265 = ($signed(_zz_8266) * $signed(twiddle_factor_table_21_imag));
  assign _zz_8266 = ($signed(data_mid_4_54_real) + $signed(data_mid_4_54_imag));
  assign _zz_8267 = fixTo_900_dout;
  assign _zz_8268 = ($signed(_zz_753) + $signed(_zz_8269));
  assign _zz_8269 = ($signed(_zz_8270) * $signed(twiddle_factor_table_21_real));
  assign _zz_8270 = ($signed(data_mid_4_54_imag) - $signed(data_mid_4_54_real));
  assign _zz_8271 = fixTo_901_dout;
  assign _zz_8272 = _zz_8273[35 : 0];
  assign _zz_8273 = _zz_8274;
  assign _zz_8274 = ($signed(_zz_8275) >>> _zz_754);
  assign _zz_8275 = _zz_8276;
  assign _zz_8276 = ($signed(_zz_8278) - $signed(_zz_751));
  assign _zz_8277 = ({9'd0,data_mid_4_38_real} <<< 9);
  assign _zz_8278 = {{9{_zz_8277[26]}}, _zz_8277};
  assign _zz_8279 = fixTo_902_dout;
  assign _zz_8280 = _zz_8281[35 : 0];
  assign _zz_8281 = _zz_8282;
  assign _zz_8282 = ($signed(_zz_8283) >>> _zz_754);
  assign _zz_8283 = _zz_8284;
  assign _zz_8284 = ($signed(_zz_8286) - $signed(_zz_752));
  assign _zz_8285 = ({9'd0,data_mid_4_38_imag} <<< 9);
  assign _zz_8286 = {{9{_zz_8285[26]}}, _zz_8285};
  assign _zz_8287 = fixTo_903_dout;
  assign _zz_8288 = _zz_8289[35 : 0];
  assign _zz_8289 = _zz_8290;
  assign _zz_8290 = ($signed(_zz_8291) >>> _zz_755);
  assign _zz_8291 = _zz_8292;
  assign _zz_8292 = ($signed(_zz_8294) + $signed(_zz_751));
  assign _zz_8293 = ({9'd0,data_mid_4_38_real} <<< 9);
  assign _zz_8294 = {{9{_zz_8293[26]}}, _zz_8293};
  assign _zz_8295 = fixTo_904_dout;
  assign _zz_8296 = _zz_8297[35 : 0];
  assign _zz_8297 = _zz_8298;
  assign _zz_8298 = ($signed(_zz_8299) >>> _zz_755);
  assign _zz_8299 = _zz_8300;
  assign _zz_8300 = ($signed(_zz_8302) + $signed(_zz_752));
  assign _zz_8301 = ({9'd0,data_mid_4_38_imag} <<< 9);
  assign _zz_8302 = {{9{_zz_8301[26]}}, _zz_8301};
  assign _zz_8303 = fixTo_905_dout;
  assign _zz_8304 = ($signed(twiddle_factor_table_22_real) + $signed(twiddle_factor_table_22_imag));
  assign _zz_8305 = ($signed(_zz_758) - $signed(_zz_8306));
  assign _zz_8306 = ($signed(_zz_8307) * $signed(twiddle_factor_table_22_imag));
  assign _zz_8307 = ($signed(data_mid_4_55_real) + $signed(data_mid_4_55_imag));
  assign _zz_8308 = fixTo_906_dout;
  assign _zz_8309 = ($signed(_zz_758) + $signed(_zz_8310));
  assign _zz_8310 = ($signed(_zz_8311) * $signed(twiddle_factor_table_22_real));
  assign _zz_8311 = ($signed(data_mid_4_55_imag) - $signed(data_mid_4_55_real));
  assign _zz_8312 = fixTo_907_dout;
  assign _zz_8313 = _zz_8314[35 : 0];
  assign _zz_8314 = _zz_8315;
  assign _zz_8315 = ($signed(_zz_8316) >>> _zz_759);
  assign _zz_8316 = _zz_8317;
  assign _zz_8317 = ($signed(_zz_8319) - $signed(_zz_756));
  assign _zz_8318 = ({9'd0,data_mid_4_39_real} <<< 9);
  assign _zz_8319 = {{9{_zz_8318[26]}}, _zz_8318};
  assign _zz_8320 = fixTo_908_dout;
  assign _zz_8321 = _zz_8322[35 : 0];
  assign _zz_8322 = _zz_8323;
  assign _zz_8323 = ($signed(_zz_8324) >>> _zz_759);
  assign _zz_8324 = _zz_8325;
  assign _zz_8325 = ($signed(_zz_8327) - $signed(_zz_757));
  assign _zz_8326 = ({9'd0,data_mid_4_39_imag} <<< 9);
  assign _zz_8327 = {{9{_zz_8326[26]}}, _zz_8326};
  assign _zz_8328 = fixTo_909_dout;
  assign _zz_8329 = _zz_8330[35 : 0];
  assign _zz_8330 = _zz_8331;
  assign _zz_8331 = ($signed(_zz_8332) >>> _zz_760);
  assign _zz_8332 = _zz_8333;
  assign _zz_8333 = ($signed(_zz_8335) + $signed(_zz_756));
  assign _zz_8334 = ({9'd0,data_mid_4_39_real} <<< 9);
  assign _zz_8335 = {{9{_zz_8334[26]}}, _zz_8334};
  assign _zz_8336 = fixTo_910_dout;
  assign _zz_8337 = _zz_8338[35 : 0];
  assign _zz_8338 = _zz_8339;
  assign _zz_8339 = ($signed(_zz_8340) >>> _zz_760);
  assign _zz_8340 = _zz_8341;
  assign _zz_8341 = ($signed(_zz_8343) + $signed(_zz_757));
  assign _zz_8342 = ({9'd0,data_mid_4_39_imag} <<< 9);
  assign _zz_8343 = {{9{_zz_8342[26]}}, _zz_8342};
  assign _zz_8344 = fixTo_911_dout;
  assign _zz_8345 = ($signed(twiddle_factor_table_23_real) + $signed(twiddle_factor_table_23_imag));
  assign _zz_8346 = ($signed(_zz_763) - $signed(_zz_8347));
  assign _zz_8347 = ($signed(_zz_8348) * $signed(twiddle_factor_table_23_imag));
  assign _zz_8348 = ($signed(data_mid_4_56_real) + $signed(data_mid_4_56_imag));
  assign _zz_8349 = fixTo_912_dout;
  assign _zz_8350 = ($signed(_zz_763) + $signed(_zz_8351));
  assign _zz_8351 = ($signed(_zz_8352) * $signed(twiddle_factor_table_23_real));
  assign _zz_8352 = ($signed(data_mid_4_56_imag) - $signed(data_mid_4_56_real));
  assign _zz_8353 = fixTo_913_dout;
  assign _zz_8354 = _zz_8355[35 : 0];
  assign _zz_8355 = _zz_8356;
  assign _zz_8356 = ($signed(_zz_8357) >>> _zz_764);
  assign _zz_8357 = _zz_8358;
  assign _zz_8358 = ($signed(_zz_8360) - $signed(_zz_761));
  assign _zz_8359 = ({9'd0,data_mid_4_40_real} <<< 9);
  assign _zz_8360 = {{9{_zz_8359[26]}}, _zz_8359};
  assign _zz_8361 = fixTo_914_dout;
  assign _zz_8362 = _zz_8363[35 : 0];
  assign _zz_8363 = _zz_8364;
  assign _zz_8364 = ($signed(_zz_8365) >>> _zz_764);
  assign _zz_8365 = _zz_8366;
  assign _zz_8366 = ($signed(_zz_8368) - $signed(_zz_762));
  assign _zz_8367 = ({9'd0,data_mid_4_40_imag} <<< 9);
  assign _zz_8368 = {{9{_zz_8367[26]}}, _zz_8367};
  assign _zz_8369 = fixTo_915_dout;
  assign _zz_8370 = _zz_8371[35 : 0];
  assign _zz_8371 = _zz_8372;
  assign _zz_8372 = ($signed(_zz_8373) >>> _zz_765);
  assign _zz_8373 = _zz_8374;
  assign _zz_8374 = ($signed(_zz_8376) + $signed(_zz_761));
  assign _zz_8375 = ({9'd0,data_mid_4_40_real} <<< 9);
  assign _zz_8376 = {{9{_zz_8375[26]}}, _zz_8375};
  assign _zz_8377 = fixTo_916_dout;
  assign _zz_8378 = _zz_8379[35 : 0];
  assign _zz_8379 = _zz_8380;
  assign _zz_8380 = ($signed(_zz_8381) >>> _zz_765);
  assign _zz_8381 = _zz_8382;
  assign _zz_8382 = ($signed(_zz_8384) + $signed(_zz_762));
  assign _zz_8383 = ({9'd0,data_mid_4_40_imag} <<< 9);
  assign _zz_8384 = {{9{_zz_8383[26]}}, _zz_8383};
  assign _zz_8385 = fixTo_917_dout;
  assign _zz_8386 = ($signed(twiddle_factor_table_24_real) + $signed(twiddle_factor_table_24_imag));
  assign _zz_8387 = ($signed(_zz_768) - $signed(_zz_8388));
  assign _zz_8388 = ($signed(_zz_8389) * $signed(twiddle_factor_table_24_imag));
  assign _zz_8389 = ($signed(data_mid_4_57_real) + $signed(data_mid_4_57_imag));
  assign _zz_8390 = fixTo_918_dout;
  assign _zz_8391 = ($signed(_zz_768) + $signed(_zz_8392));
  assign _zz_8392 = ($signed(_zz_8393) * $signed(twiddle_factor_table_24_real));
  assign _zz_8393 = ($signed(data_mid_4_57_imag) - $signed(data_mid_4_57_real));
  assign _zz_8394 = fixTo_919_dout;
  assign _zz_8395 = _zz_8396[35 : 0];
  assign _zz_8396 = _zz_8397;
  assign _zz_8397 = ($signed(_zz_8398) >>> _zz_769);
  assign _zz_8398 = _zz_8399;
  assign _zz_8399 = ($signed(_zz_8401) - $signed(_zz_766));
  assign _zz_8400 = ({9'd0,data_mid_4_41_real} <<< 9);
  assign _zz_8401 = {{9{_zz_8400[26]}}, _zz_8400};
  assign _zz_8402 = fixTo_920_dout;
  assign _zz_8403 = _zz_8404[35 : 0];
  assign _zz_8404 = _zz_8405;
  assign _zz_8405 = ($signed(_zz_8406) >>> _zz_769);
  assign _zz_8406 = _zz_8407;
  assign _zz_8407 = ($signed(_zz_8409) - $signed(_zz_767));
  assign _zz_8408 = ({9'd0,data_mid_4_41_imag} <<< 9);
  assign _zz_8409 = {{9{_zz_8408[26]}}, _zz_8408};
  assign _zz_8410 = fixTo_921_dout;
  assign _zz_8411 = _zz_8412[35 : 0];
  assign _zz_8412 = _zz_8413;
  assign _zz_8413 = ($signed(_zz_8414) >>> _zz_770);
  assign _zz_8414 = _zz_8415;
  assign _zz_8415 = ($signed(_zz_8417) + $signed(_zz_766));
  assign _zz_8416 = ({9'd0,data_mid_4_41_real} <<< 9);
  assign _zz_8417 = {{9{_zz_8416[26]}}, _zz_8416};
  assign _zz_8418 = fixTo_922_dout;
  assign _zz_8419 = _zz_8420[35 : 0];
  assign _zz_8420 = _zz_8421;
  assign _zz_8421 = ($signed(_zz_8422) >>> _zz_770);
  assign _zz_8422 = _zz_8423;
  assign _zz_8423 = ($signed(_zz_8425) + $signed(_zz_767));
  assign _zz_8424 = ({9'd0,data_mid_4_41_imag} <<< 9);
  assign _zz_8425 = {{9{_zz_8424[26]}}, _zz_8424};
  assign _zz_8426 = fixTo_923_dout;
  assign _zz_8427 = ($signed(twiddle_factor_table_25_real) + $signed(twiddle_factor_table_25_imag));
  assign _zz_8428 = ($signed(_zz_773) - $signed(_zz_8429));
  assign _zz_8429 = ($signed(_zz_8430) * $signed(twiddle_factor_table_25_imag));
  assign _zz_8430 = ($signed(data_mid_4_58_real) + $signed(data_mid_4_58_imag));
  assign _zz_8431 = fixTo_924_dout;
  assign _zz_8432 = ($signed(_zz_773) + $signed(_zz_8433));
  assign _zz_8433 = ($signed(_zz_8434) * $signed(twiddle_factor_table_25_real));
  assign _zz_8434 = ($signed(data_mid_4_58_imag) - $signed(data_mid_4_58_real));
  assign _zz_8435 = fixTo_925_dout;
  assign _zz_8436 = _zz_8437[35 : 0];
  assign _zz_8437 = _zz_8438;
  assign _zz_8438 = ($signed(_zz_8439) >>> _zz_774);
  assign _zz_8439 = _zz_8440;
  assign _zz_8440 = ($signed(_zz_8442) - $signed(_zz_771));
  assign _zz_8441 = ({9'd0,data_mid_4_42_real} <<< 9);
  assign _zz_8442 = {{9{_zz_8441[26]}}, _zz_8441};
  assign _zz_8443 = fixTo_926_dout;
  assign _zz_8444 = _zz_8445[35 : 0];
  assign _zz_8445 = _zz_8446;
  assign _zz_8446 = ($signed(_zz_8447) >>> _zz_774);
  assign _zz_8447 = _zz_8448;
  assign _zz_8448 = ($signed(_zz_8450) - $signed(_zz_772));
  assign _zz_8449 = ({9'd0,data_mid_4_42_imag} <<< 9);
  assign _zz_8450 = {{9{_zz_8449[26]}}, _zz_8449};
  assign _zz_8451 = fixTo_927_dout;
  assign _zz_8452 = _zz_8453[35 : 0];
  assign _zz_8453 = _zz_8454;
  assign _zz_8454 = ($signed(_zz_8455) >>> _zz_775);
  assign _zz_8455 = _zz_8456;
  assign _zz_8456 = ($signed(_zz_8458) + $signed(_zz_771));
  assign _zz_8457 = ({9'd0,data_mid_4_42_real} <<< 9);
  assign _zz_8458 = {{9{_zz_8457[26]}}, _zz_8457};
  assign _zz_8459 = fixTo_928_dout;
  assign _zz_8460 = _zz_8461[35 : 0];
  assign _zz_8461 = _zz_8462;
  assign _zz_8462 = ($signed(_zz_8463) >>> _zz_775);
  assign _zz_8463 = _zz_8464;
  assign _zz_8464 = ($signed(_zz_8466) + $signed(_zz_772));
  assign _zz_8465 = ({9'd0,data_mid_4_42_imag} <<< 9);
  assign _zz_8466 = {{9{_zz_8465[26]}}, _zz_8465};
  assign _zz_8467 = fixTo_929_dout;
  assign _zz_8468 = ($signed(twiddle_factor_table_26_real) + $signed(twiddle_factor_table_26_imag));
  assign _zz_8469 = ($signed(_zz_778) - $signed(_zz_8470));
  assign _zz_8470 = ($signed(_zz_8471) * $signed(twiddle_factor_table_26_imag));
  assign _zz_8471 = ($signed(data_mid_4_59_real) + $signed(data_mid_4_59_imag));
  assign _zz_8472 = fixTo_930_dout;
  assign _zz_8473 = ($signed(_zz_778) + $signed(_zz_8474));
  assign _zz_8474 = ($signed(_zz_8475) * $signed(twiddle_factor_table_26_real));
  assign _zz_8475 = ($signed(data_mid_4_59_imag) - $signed(data_mid_4_59_real));
  assign _zz_8476 = fixTo_931_dout;
  assign _zz_8477 = _zz_8478[35 : 0];
  assign _zz_8478 = _zz_8479;
  assign _zz_8479 = ($signed(_zz_8480) >>> _zz_779);
  assign _zz_8480 = _zz_8481;
  assign _zz_8481 = ($signed(_zz_8483) - $signed(_zz_776));
  assign _zz_8482 = ({9'd0,data_mid_4_43_real} <<< 9);
  assign _zz_8483 = {{9{_zz_8482[26]}}, _zz_8482};
  assign _zz_8484 = fixTo_932_dout;
  assign _zz_8485 = _zz_8486[35 : 0];
  assign _zz_8486 = _zz_8487;
  assign _zz_8487 = ($signed(_zz_8488) >>> _zz_779);
  assign _zz_8488 = _zz_8489;
  assign _zz_8489 = ($signed(_zz_8491) - $signed(_zz_777));
  assign _zz_8490 = ({9'd0,data_mid_4_43_imag} <<< 9);
  assign _zz_8491 = {{9{_zz_8490[26]}}, _zz_8490};
  assign _zz_8492 = fixTo_933_dout;
  assign _zz_8493 = _zz_8494[35 : 0];
  assign _zz_8494 = _zz_8495;
  assign _zz_8495 = ($signed(_zz_8496) >>> _zz_780);
  assign _zz_8496 = _zz_8497;
  assign _zz_8497 = ($signed(_zz_8499) + $signed(_zz_776));
  assign _zz_8498 = ({9'd0,data_mid_4_43_real} <<< 9);
  assign _zz_8499 = {{9{_zz_8498[26]}}, _zz_8498};
  assign _zz_8500 = fixTo_934_dout;
  assign _zz_8501 = _zz_8502[35 : 0];
  assign _zz_8502 = _zz_8503;
  assign _zz_8503 = ($signed(_zz_8504) >>> _zz_780);
  assign _zz_8504 = _zz_8505;
  assign _zz_8505 = ($signed(_zz_8507) + $signed(_zz_777));
  assign _zz_8506 = ({9'd0,data_mid_4_43_imag} <<< 9);
  assign _zz_8507 = {{9{_zz_8506[26]}}, _zz_8506};
  assign _zz_8508 = fixTo_935_dout;
  assign _zz_8509 = ($signed(twiddle_factor_table_27_real) + $signed(twiddle_factor_table_27_imag));
  assign _zz_8510 = ($signed(_zz_783) - $signed(_zz_8511));
  assign _zz_8511 = ($signed(_zz_8512) * $signed(twiddle_factor_table_27_imag));
  assign _zz_8512 = ($signed(data_mid_4_60_real) + $signed(data_mid_4_60_imag));
  assign _zz_8513 = fixTo_936_dout;
  assign _zz_8514 = ($signed(_zz_783) + $signed(_zz_8515));
  assign _zz_8515 = ($signed(_zz_8516) * $signed(twiddle_factor_table_27_real));
  assign _zz_8516 = ($signed(data_mid_4_60_imag) - $signed(data_mid_4_60_real));
  assign _zz_8517 = fixTo_937_dout;
  assign _zz_8518 = _zz_8519[35 : 0];
  assign _zz_8519 = _zz_8520;
  assign _zz_8520 = ($signed(_zz_8521) >>> _zz_784);
  assign _zz_8521 = _zz_8522;
  assign _zz_8522 = ($signed(_zz_8524) - $signed(_zz_781));
  assign _zz_8523 = ({9'd0,data_mid_4_44_real} <<< 9);
  assign _zz_8524 = {{9{_zz_8523[26]}}, _zz_8523};
  assign _zz_8525 = fixTo_938_dout;
  assign _zz_8526 = _zz_8527[35 : 0];
  assign _zz_8527 = _zz_8528;
  assign _zz_8528 = ($signed(_zz_8529) >>> _zz_784);
  assign _zz_8529 = _zz_8530;
  assign _zz_8530 = ($signed(_zz_8532) - $signed(_zz_782));
  assign _zz_8531 = ({9'd0,data_mid_4_44_imag} <<< 9);
  assign _zz_8532 = {{9{_zz_8531[26]}}, _zz_8531};
  assign _zz_8533 = fixTo_939_dout;
  assign _zz_8534 = _zz_8535[35 : 0];
  assign _zz_8535 = _zz_8536;
  assign _zz_8536 = ($signed(_zz_8537) >>> _zz_785);
  assign _zz_8537 = _zz_8538;
  assign _zz_8538 = ($signed(_zz_8540) + $signed(_zz_781));
  assign _zz_8539 = ({9'd0,data_mid_4_44_real} <<< 9);
  assign _zz_8540 = {{9{_zz_8539[26]}}, _zz_8539};
  assign _zz_8541 = fixTo_940_dout;
  assign _zz_8542 = _zz_8543[35 : 0];
  assign _zz_8543 = _zz_8544;
  assign _zz_8544 = ($signed(_zz_8545) >>> _zz_785);
  assign _zz_8545 = _zz_8546;
  assign _zz_8546 = ($signed(_zz_8548) + $signed(_zz_782));
  assign _zz_8547 = ({9'd0,data_mid_4_44_imag} <<< 9);
  assign _zz_8548 = {{9{_zz_8547[26]}}, _zz_8547};
  assign _zz_8549 = fixTo_941_dout;
  assign _zz_8550 = ($signed(twiddle_factor_table_28_real) + $signed(twiddle_factor_table_28_imag));
  assign _zz_8551 = ($signed(_zz_788) - $signed(_zz_8552));
  assign _zz_8552 = ($signed(_zz_8553) * $signed(twiddle_factor_table_28_imag));
  assign _zz_8553 = ($signed(data_mid_4_61_real) + $signed(data_mid_4_61_imag));
  assign _zz_8554 = fixTo_942_dout;
  assign _zz_8555 = ($signed(_zz_788) + $signed(_zz_8556));
  assign _zz_8556 = ($signed(_zz_8557) * $signed(twiddle_factor_table_28_real));
  assign _zz_8557 = ($signed(data_mid_4_61_imag) - $signed(data_mid_4_61_real));
  assign _zz_8558 = fixTo_943_dout;
  assign _zz_8559 = _zz_8560[35 : 0];
  assign _zz_8560 = _zz_8561;
  assign _zz_8561 = ($signed(_zz_8562) >>> _zz_789);
  assign _zz_8562 = _zz_8563;
  assign _zz_8563 = ($signed(_zz_8565) - $signed(_zz_786));
  assign _zz_8564 = ({9'd0,data_mid_4_45_real} <<< 9);
  assign _zz_8565 = {{9{_zz_8564[26]}}, _zz_8564};
  assign _zz_8566 = fixTo_944_dout;
  assign _zz_8567 = _zz_8568[35 : 0];
  assign _zz_8568 = _zz_8569;
  assign _zz_8569 = ($signed(_zz_8570) >>> _zz_789);
  assign _zz_8570 = _zz_8571;
  assign _zz_8571 = ($signed(_zz_8573) - $signed(_zz_787));
  assign _zz_8572 = ({9'd0,data_mid_4_45_imag} <<< 9);
  assign _zz_8573 = {{9{_zz_8572[26]}}, _zz_8572};
  assign _zz_8574 = fixTo_945_dout;
  assign _zz_8575 = _zz_8576[35 : 0];
  assign _zz_8576 = _zz_8577;
  assign _zz_8577 = ($signed(_zz_8578) >>> _zz_790);
  assign _zz_8578 = _zz_8579;
  assign _zz_8579 = ($signed(_zz_8581) + $signed(_zz_786));
  assign _zz_8580 = ({9'd0,data_mid_4_45_real} <<< 9);
  assign _zz_8581 = {{9{_zz_8580[26]}}, _zz_8580};
  assign _zz_8582 = fixTo_946_dout;
  assign _zz_8583 = _zz_8584[35 : 0];
  assign _zz_8584 = _zz_8585;
  assign _zz_8585 = ($signed(_zz_8586) >>> _zz_790);
  assign _zz_8586 = _zz_8587;
  assign _zz_8587 = ($signed(_zz_8589) + $signed(_zz_787));
  assign _zz_8588 = ({9'd0,data_mid_4_45_imag} <<< 9);
  assign _zz_8589 = {{9{_zz_8588[26]}}, _zz_8588};
  assign _zz_8590 = fixTo_947_dout;
  assign _zz_8591 = ($signed(twiddle_factor_table_29_real) + $signed(twiddle_factor_table_29_imag));
  assign _zz_8592 = ($signed(_zz_793) - $signed(_zz_8593));
  assign _zz_8593 = ($signed(_zz_8594) * $signed(twiddle_factor_table_29_imag));
  assign _zz_8594 = ($signed(data_mid_4_62_real) + $signed(data_mid_4_62_imag));
  assign _zz_8595 = fixTo_948_dout;
  assign _zz_8596 = ($signed(_zz_793) + $signed(_zz_8597));
  assign _zz_8597 = ($signed(_zz_8598) * $signed(twiddle_factor_table_29_real));
  assign _zz_8598 = ($signed(data_mid_4_62_imag) - $signed(data_mid_4_62_real));
  assign _zz_8599 = fixTo_949_dout;
  assign _zz_8600 = _zz_8601[35 : 0];
  assign _zz_8601 = _zz_8602;
  assign _zz_8602 = ($signed(_zz_8603) >>> _zz_794);
  assign _zz_8603 = _zz_8604;
  assign _zz_8604 = ($signed(_zz_8606) - $signed(_zz_791));
  assign _zz_8605 = ({9'd0,data_mid_4_46_real} <<< 9);
  assign _zz_8606 = {{9{_zz_8605[26]}}, _zz_8605};
  assign _zz_8607 = fixTo_950_dout;
  assign _zz_8608 = _zz_8609[35 : 0];
  assign _zz_8609 = _zz_8610;
  assign _zz_8610 = ($signed(_zz_8611) >>> _zz_794);
  assign _zz_8611 = _zz_8612;
  assign _zz_8612 = ($signed(_zz_8614) - $signed(_zz_792));
  assign _zz_8613 = ({9'd0,data_mid_4_46_imag} <<< 9);
  assign _zz_8614 = {{9{_zz_8613[26]}}, _zz_8613};
  assign _zz_8615 = fixTo_951_dout;
  assign _zz_8616 = _zz_8617[35 : 0];
  assign _zz_8617 = _zz_8618;
  assign _zz_8618 = ($signed(_zz_8619) >>> _zz_795);
  assign _zz_8619 = _zz_8620;
  assign _zz_8620 = ($signed(_zz_8622) + $signed(_zz_791));
  assign _zz_8621 = ({9'd0,data_mid_4_46_real} <<< 9);
  assign _zz_8622 = {{9{_zz_8621[26]}}, _zz_8621};
  assign _zz_8623 = fixTo_952_dout;
  assign _zz_8624 = _zz_8625[35 : 0];
  assign _zz_8625 = _zz_8626;
  assign _zz_8626 = ($signed(_zz_8627) >>> _zz_795);
  assign _zz_8627 = _zz_8628;
  assign _zz_8628 = ($signed(_zz_8630) + $signed(_zz_792));
  assign _zz_8629 = ({9'd0,data_mid_4_46_imag} <<< 9);
  assign _zz_8630 = {{9{_zz_8629[26]}}, _zz_8629};
  assign _zz_8631 = fixTo_953_dout;
  assign _zz_8632 = ($signed(twiddle_factor_table_30_real) + $signed(twiddle_factor_table_30_imag));
  assign _zz_8633 = ($signed(_zz_798) - $signed(_zz_8634));
  assign _zz_8634 = ($signed(_zz_8635) * $signed(twiddle_factor_table_30_imag));
  assign _zz_8635 = ($signed(data_mid_4_63_real) + $signed(data_mid_4_63_imag));
  assign _zz_8636 = fixTo_954_dout;
  assign _zz_8637 = ($signed(_zz_798) + $signed(_zz_8638));
  assign _zz_8638 = ($signed(_zz_8639) * $signed(twiddle_factor_table_30_real));
  assign _zz_8639 = ($signed(data_mid_4_63_imag) - $signed(data_mid_4_63_real));
  assign _zz_8640 = fixTo_955_dout;
  assign _zz_8641 = _zz_8642[35 : 0];
  assign _zz_8642 = _zz_8643;
  assign _zz_8643 = ($signed(_zz_8644) >>> _zz_799);
  assign _zz_8644 = _zz_8645;
  assign _zz_8645 = ($signed(_zz_8647) - $signed(_zz_796));
  assign _zz_8646 = ({9'd0,data_mid_4_47_real} <<< 9);
  assign _zz_8647 = {{9{_zz_8646[26]}}, _zz_8646};
  assign _zz_8648 = fixTo_956_dout;
  assign _zz_8649 = _zz_8650[35 : 0];
  assign _zz_8650 = _zz_8651;
  assign _zz_8651 = ($signed(_zz_8652) >>> _zz_799);
  assign _zz_8652 = _zz_8653;
  assign _zz_8653 = ($signed(_zz_8655) - $signed(_zz_797));
  assign _zz_8654 = ({9'd0,data_mid_4_47_imag} <<< 9);
  assign _zz_8655 = {{9{_zz_8654[26]}}, _zz_8654};
  assign _zz_8656 = fixTo_957_dout;
  assign _zz_8657 = _zz_8658[35 : 0];
  assign _zz_8658 = _zz_8659;
  assign _zz_8659 = ($signed(_zz_8660) >>> _zz_800);
  assign _zz_8660 = _zz_8661;
  assign _zz_8661 = ($signed(_zz_8663) + $signed(_zz_796));
  assign _zz_8662 = ({9'd0,data_mid_4_47_real} <<< 9);
  assign _zz_8663 = {{9{_zz_8662[26]}}, _zz_8662};
  assign _zz_8664 = fixTo_958_dout;
  assign _zz_8665 = _zz_8666[35 : 0];
  assign _zz_8666 = _zz_8667;
  assign _zz_8667 = ($signed(_zz_8668) >>> _zz_800);
  assign _zz_8668 = _zz_8669;
  assign _zz_8669 = ($signed(_zz_8671) + $signed(_zz_797));
  assign _zz_8670 = ({9'd0,data_mid_4_47_imag} <<< 9);
  assign _zz_8671 = {{9{_zz_8670[26]}}, _zz_8670};
  assign _zz_8672 = fixTo_959_dout;
  assign _zz_8673 = ($signed(twiddle_factor_table_31_real) + $signed(twiddle_factor_table_31_imag));
  assign _zz_8674 = ($signed(_zz_803) - $signed(_zz_8675));
  assign _zz_8675 = ($signed(_zz_8676) * $signed(twiddle_factor_table_31_imag));
  assign _zz_8676 = ($signed(data_mid_5_32_real) + $signed(data_mid_5_32_imag));
  assign _zz_8677 = fixTo_960_dout;
  assign _zz_8678 = ($signed(_zz_803) + $signed(_zz_8679));
  assign _zz_8679 = ($signed(_zz_8680) * $signed(twiddle_factor_table_31_real));
  assign _zz_8680 = ($signed(data_mid_5_32_imag) - $signed(data_mid_5_32_real));
  assign _zz_8681 = fixTo_961_dout;
  assign _zz_8682 = _zz_8683[35 : 0];
  assign _zz_8683 = _zz_8684;
  assign _zz_8684 = ($signed(_zz_8685) >>> _zz_804);
  assign _zz_8685 = _zz_8686;
  assign _zz_8686 = ($signed(_zz_8688) - $signed(_zz_801));
  assign _zz_8687 = ({9'd0,data_mid_5_0_real} <<< 9);
  assign _zz_8688 = {{9{_zz_8687[26]}}, _zz_8687};
  assign _zz_8689 = fixTo_962_dout;
  assign _zz_8690 = _zz_8691[35 : 0];
  assign _zz_8691 = _zz_8692;
  assign _zz_8692 = ($signed(_zz_8693) >>> _zz_804);
  assign _zz_8693 = _zz_8694;
  assign _zz_8694 = ($signed(_zz_8696) - $signed(_zz_802));
  assign _zz_8695 = ({9'd0,data_mid_5_0_imag} <<< 9);
  assign _zz_8696 = {{9{_zz_8695[26]}}, _zz_8695};
  assign _zz_8697 = fixTo_963_dout;
  assign _zz_8698 = _zz_8699[35 : 0];
  assign _zz_8699 = _zz_8700;
  assign _zz_8700 = ($signed(_zz_8701) >>> _zz_805);
  assign _zz_8701 = _zz_8702;
  assign _zz_8702 = ($signed(_zz_8704) + $signed(_zz_801));
  assign _zz_8703 = ({9'd0,data_mid_5_0_real} <<< 9);
  assign _zz_8704 = {{9{_zz_8703[26]}}, _zz_8703};
  assign _zz_8705 = fixTo_964_dout;
  assign _zz_8706 = _zz_8707[35 : 0];
  assign _zz_8707 = _zz_8708;
  assign _zz_8708 = ($signed(_zz_8709) >>> _zz_805);
  assign _zz_8709 = _zz_8710;
  assign _zz_8710 = ($signed(_zz_8712) + $signed(_zz_802));
  assign _zz_8711 = ({9'd0,data_mid_5_0_imag} <<< 9);
  assign _zz_8712 = {{9{_zz_8711[26]}}, _zz_8711};
  assign _zz_8713 = fixTo_965_dout;
  assign _zz_8714 = ($signed(twiddle_factor_table_32_real) + $signed(twiddle_factor_table_32_imag));
  assign _zz_8715 = ($signed(_zz_808) - $signed(_zz_8716));
  assign _zz_8716 = ($signed(_zz_8717) * $signed(twiddle_factor_table_32_imag));
  assign _zz_8717 = ($signed(data_mid_5_33_real) + $signed(data_mid_5_33_imag));
  assign _zz_8718 = fixTo_966_dout;
  assign _zz_8719 = ($signed(_zz_808) + $signed(_zz_8720));
  assign _zz_8720 = ($signed(_zz_8721) * $signed(twiddle_factor_table_32_real));
  assign _zz_8721 = ($signed(data_mid_5_33_imag) - $signed(data_mid_5_33_real));
  assign _zz_8722 = fixTo_967_dout;
  assign _zz_8723 = _zz_8724[35 : 0];
  assign _zz_8724 = _zz_8725;
  assign _zz_8725 = ($signed(_zz_8726) >>> _zz_809);
  assign _zz_8726 = _zz_8727;
  assign _zz_8727 = ($signed(_zz_8729) - $signed(_zz_806));
  assign _zz_8728 = ({9'd0,data_mid_5_1_real} <<< 9);
  assign _zz_8729 = {{9{_zz_8728[26]}}, _zz_8728};
  assign _zz_8730 = fixTo_968_dout;
  assign _zz_8731 = _zz_8732[35 : 0];
  assign _zz_8732 = _zz_8733;
  assign _zz_8733 = ($signed(_zz_8734) >>> _zz_809);
  assign _zz_8734 = _zz_8735;
  assign _zz_8735 = ($signed(_zz_8737) - $signed(_zz_807));
  assign _zz_8736 = ({9'd0,data_mid_5_1_imag} <<< 9);
  assign _zz_8737 = {{9{_zz_8736[26]}}, _zz_8736};
  assign _zz_8738 = fixTo_969_dout;
  assign _zz_8739 = _zz_8740[35 : 0];
  assign _zz_8740 = _zz_8741;
  assign _zz_8741 = ($signed(_zz_8742) >>> _zz_810);
  assign _zz_8742 = _zz_8743;
  assign _zz_8743 = ($signed(_zz_8745) + $signed(_zz_806));
  assign _zz_8744 = ({9'd0,data_mid_5_1_real} <<< 9);
  assign _zz_8745 = {{9{_zz_8744[26]}}, _zz_8744};
  assign _zz_8746 = fixTo_970_dout;
  assign _zz_8747 = _zz_8748[35 : 0];
  assign _zz_8748 = _zz_8749;
  assign _zz_8749 = ($signed(_zz_8750) >>> _zz_810);
  assign _zz_8750 = _zz_8751;
  assign _zz_8751 = ($signed(_zz_8753) + $signed(_zz_807));
  assign _zz_8752 = ({9'd0,data_mid_5_1_imag} <<< 9);
  assign _zz_8753 = {{9{_zz_8752[26]}}, _zz_8752};
  assign _zz_8754 = fixTo_971_dout;
  assign _zz_8755 = ($signed(twiddle_factor_table_33_real) + $signed(twiddle_factor_table_33_imag));
  assign _zz_8756 = ($signed(_zz_813) - $signed(_zz_8757));
  assign _zz_8757 = ($signed(_zz_8758) * $signed(twiddle_factor_table_33_imag));
  assign _zz_8758 = ($signed(data_mid_5_34_real) + $signed(data_mid_5_34_imag));
  assign _zz_8759 = fixTo_972_dout;
  assign _zz_8760 = ($signed(_zz_813) + $signed(_zz_8761));
  assign _zz_8761 = ($signed(_zz_8762) * $signed(twiddle_factor_table_33_real));
  assign _zz_8762 = ($signed(data_mid_5_34_imag) - $signed(data_mid_5_34_real));
  assign _zz_8763 = fixTo_973_dout;
  assign _zz_8764 = _zz_8765[35 : 0];
  assign _zz_8765 = _zz_8766;
  assign _zz_8766 = ($signed(_zz_8767) >>> _zz_814);
  assign _zz_8767 = _zz_8768;
  assign _zz_8768 = ($signed(_zz_8770) - $signed(_zz_811));
  assign _zz_8769 = ({9'd0,data_mid_5_2_real} <<< 9);
  assign _zz_8770 = {{9{_zz_8769[26]}}, _zz_8769};
  assign _zz_8771 = fixTo_974_dout;
  assign _zz_8772 = _zz_8773[35 : 0];
  assign _zz_8773 = _zz_8774;
  assign _zz_8774 = ($signed(_zz_8775) >>> _zz_814);
  assign _zz_8775 = _zz_8776;
  assign _zz_8776 = ($signed(_zz_8778) - $signed(_zz_812));
  assign _zz_8777 = ({9'd0,data_mid_5_2_imag} <<< 9);
  assign _zz_8778 = {{9{_zz_8777[26]}}, _zz_8777};
  assign _zz_8779 = fixTo_975_dout;
  assign _zz_8780 = _zz_8781[35 : 0];
  assign _zz_8781 = _zz_8782;
  assign _zz_8782 = ($signed(_zz_8783) >>> _zz_815);
  assign _zz_8783 = _zz_8784;
  assign _zz_8784 = ($signed(_zz_8786) + $signed(_zz_811));
  assign _zz_8785 = ({9'd0,data_mid_5_2_real} <<< 9);
  assign _zz_8786 = {{9{_zz_8785[26]}}, _zz_8785};
  assign _zz_8787 = fixTo_976_dout;
  assign _zz_8788 = _zz_8789[35 : 0];
  assign _zz_8789 = _zz_8790;
  assign _zz_8790 = ($signed(_zz_8791) >>> _zz_815);
  assign _zz_8791 = _zz_8792;
  assign _zz_8792 = ($signed(_zz_8794) + $signed(_zz_812));
  assign _zz_8793 = ({9'd0,data_mid_5_2_imag} <<< 9);
  assign _zz_8794 = {{9{_zz_8793[26]}}, _zz_8793};
  assign _zz_8795 = fixTo_977_dout;
  assign _zz_8796 = ($signed(twiddle_factor_table_34_real) + $signed(twiddle_factor_table_34_imag));
  assign _zz_8797 = ($signed(_zz_818) - $signed(_zz_8798));
  assign _zz_8798 = ($signed(_zz_8799) * $signed(twiddle_factor_table_34_imag));
  assign _zz_8799 = ($signed(data_mid_5_35_real) + $signed(data_mid_5_35_imag));
  assign _zz_8800 = fixTo_978_dout;
  assign _zz_8801 = ($signed(_zz_818) + $signed(_zz_8802));
  assign _zz_8802 = ($signed(_zz_8803) * $signed(twiddle_factor_table_34_real));
  assign _zz_8803 = ($signed(data_mid_5_35_imag) - $signed(data_mid_5_35_real));
  assign _zz_8804 = fixTo_979_dout;
  assign _zz_8805 = _zz_8806[35 : 0];
  assign _zz_8806 = _zz_8807;
  assign _zz_8807 = ($signed(_zz_8808) >>> _zz_819);
  assign _zz_8808 = _zz_8809;
  assign _zz_8809 = ($signed(_zz_8811) - $signed(_zz_816));
  assign _zz_8810 = ({9'd0,data_mid_5_3_real} <<< 9);
  assign _zz_8811 = {{9{_zz_8810[26]}}, _zz_8810};
  assign _zz_8812 = fixTo_980_dout;
  assign _zz_8813 = _zz_8814[35 : 0];
  assign _zz_8814 = _zz_8815;
  assign _zz_8815 = ($signed(_zz_8816) >>> _zz_819);
  assign _zz_8816 = _zz_8817;
  assign _zz_8817 = ($signed(_zz_8819) - $signed(_zz_817));
  assign _zz_8818 = ({9'd0,data_mid_5_3_imag} <<< 9);
  assign _zz_8819 = {{9{_zz_8818[26]}}, _zz_8818};
  assign _zz_8820 = fixTo_981_dout;
  assign _zz_8821 = _zz_8822[35 : 0];
  assign _zz_8822 = _zz_8823;
  assign _zz_8823 = ($signed(_zz_8824) >>> _zz_820);
  assign _zz_8824 = _zz_8825;
  assign _zz_8825 = ($signed(_zz_8827) + $signed(_zz_816));
  assign _zz_8826 = ({9'd0,data_mid_5_3_real} <<< 9);
  assign _zz_8827 = {{9{_zz_8826[26]}}, _zz_8826};
  assign _zz_8828 = fixTo_982_dout;
  assign _zz_8829 = _zz_8830[35 : 0];
  assign _zz_8830 = _zz_8831;
  assign _zz_8831 = ($signed(_zz_8832) >>> _zz_820);
  assign _zz_8832 = _zz_8833;
  assign _zz_8833 = ($signed(_zz_8835) + $signed(_zz_817));
  assign _zz_8834 = ({9'd0,data_mid_5_3_imag} <<< 9);
  assign _zz_8835 = {{9{_zz_8834[26]}}, _zz_8834};
  assign _zz_8836 = fixTo_983_dout;
  assign _zz_8837 = ($signed(twiddle_factor_table_35_real) + $signed(twiddle_factor_table_35_imag));
  assign _zz_8838 = ($signed(_zz_823) - $signed(_zz_8839));
  assign _zz_8839 = ($signed(_zz_8840) * $signed(twiddle_factor_table_35_imag));
  assign _zz_8840 = ($signed(data_mid_5_36_real) + $signed(data_mid_5_36_imag));
  assign _zz_8841 = fixTo_984_dout;
  assign _zz_8842 = ($signed(_zz_823) + $signed(_zz_8843));
  assign _zz_8843 = ($signed(_zz_8844) * $signed(twiddle_factor_table_35_real));
  assign _zz_8844 = ($signed(data_mid_5_36_imag) - $signed(data_mid_5_36_real));
  assign _zz_8845 = fixTo_985_dout;
  assign _zz_8846 = _zz_8847[35 : 0];
  assign _zz_8847 = _zz_8848;
  assign _zz_8848 = ($signed(_zz_8849) >>> _zz_824);
  assign _zz_8849 = _zz_8850;
  assign _zz_8850 = ($signed(_zz_8852) - $signed(_zz_821));
  assign _zz_8851 = ({9'd0,data_mid_5_4_real} <<< 9);
  assign _zz_8852 = {{9{_zz_8851[26]}}, _zz_8851};
  assign _zz_8853 = fixTo_986_dout;
  assign _zz_8854 = _zz_8855[35 : 0];
  assign _zz_8855 = _zz_8856;
  assign _zz_8856 = ($signed(_zz_8857) >>> _zz_824);
  assign _zz_8857 = _zz_8858;
  assign _zz_8858 = ($signed(_zz_8860) - $signed(_zz_822));
  assign _zz_8859 = ({9'd0,data_mid_5_4_imag} <<< 9);
  assign _zz_8860 = {{9{_zz_8859[26]}}, _zz_8859};
  assign _zz_8861 = fixTo_987_dout;
  assign _zz_8862 = _zz_8863[35 : 0];
  assign _zz_8863 = _zz_8864;
  assign _zz_8864 = ($signed(_zz_8865) >>> _zz_825);
  assign _zz_8865 = _zz_8866;
  assign _zz_8866 = ($signed(_zz_8868) + $signed(_zz_821));
  assign _zz_8867 = ({9'd0,data_mid_5_4_real} <<< 9);
  assign _zz_8868 = {{9{_zz_8867[26]}}, _zz_8867};
  assign _zz_8869 = fixTo_988_dout;
  assign _zz_8870 = _zz_8871[35 : 0];
  assign _zz_8871 = _zz_8872;
  assign _zz_8872 = ($signed(_zz_8873) >>> _zz_825);
  assign _zz_8873 = _zz_8874;
  assign _zz_8874 = ($signed(_zz_8876) + $signed(_zz_822));
  assign _zz_8875 = ({9'd0,data_mid_5_4_imag} <<< 9);
  assign _zz_8876 = {{9{_zz_8875[26]}}, _zz_8875};
  assign _zz_8877 = fixTo_989_dout;
  assign _zz_8878 = ($signed(twiddle_factor_table_36_real) + $signed(twiddle_factor_table_36_imag));
  assign _zz_8879 = ($signed(_zz_828) - $signed(_zz_8880));
  assign _zz_8880 = ($signed(_zz_8881) * $signed(twiddle_factor_table_36_imag));
  assign _zz_8881 = ($signed(data_mid_5_37_real) + $signed(data_mid_5_37_imag));
  assign _zz_8882 = fixTo_990_dout;
  assign _zz_8883 = ($signed(_zz_828) + $signed(_zz_8884));
  assign _zz_8884 = ($signed(_zz_8885) * $signed(twiddle_factor_table_36_real));
  assign _zz_8885 = ($signed(data_mid_5_37_imag) - $signed(data_mid_5_37_real));
  assign _zz_8886 = fixTo_991_dout;
  assign _zz_8887 = _zz_8888[35 : 0];
  assign _zz_8888 = _zz_8889;
  assign _zz_8889 = ($signed(_zz_8890) >>> _zz_829);
  assign _zz_8890 = _zz_8891;
  assign _zz_8891 = ($signed(_zz_8893) - $signed(_zz_826));
  assign _zz_8892 = ({9'd0,data_mid_5_5_real} <<< 9);
  assign _zz_8893 = {{9{_zz_8892[26]}}, _zz_8892};
  assign _zz_8894 = fixTo_992_dout;
  assign _zz_8895 = _zz_8896[35 : 0];
  assign _zz_8896 = _zz_8897;
  assign _zz_8897 = ($signed(_zz_8898) >>> _zz_829);
  assign _zz_8898 = _zz_8899;
  assign _zz_8899 = ($signed(_zz_8901) - $signed(_zz_827));
  assign _zz_8900 = ({9'd0,data_mid_5_5_imag} <<< 9);
  assign _zz_8901 = {{9{_zz_8900[26]}}, _zz_8900};
  assign _zz_8902 = fixTo_993_dout;
  assign _zz_8903 = _zz_8904[35 : 0];
  assign _zz_8904 = _zz_8905;
  assign _zz_8905 = ($signed(_zz_8906) >>> _zz_830);
  assign _zz_8906 = _zz_8907;
  assign _zz_8907 = ($signed(_zz_8909) + $signed(_zz_826));
  assign _zz_8908 = ({9'd0,data_mid_5_5_real} <<< 9);
  assign _zz_8909 = {{9{_zz_8908[26]}}, _zz_8908};
  assign _zz_8910 = fixTo_994_dout;
  assign _zz_8911 = _zz_8912[35 : 0];
  assign _zz_8912 = _zz_8913;
  assign _zz_8913 = ($signed(_zz_8914) >>> _zz_830);
  assign _zz_8914 = _zz_8915;
  assign _zz_8915 = ($signed(_zz_8917) + $signed(_zz_827));
  assign _zz_8916 = ({9'd0,data_mid_5_5_imag} <<< 9);
  assign _zz_8917 = {{9{_zz_8916[26]}}, _zz_8916};
  assign _zz_8918 = fixTo_995_dout;
  assign _zz_8919 = ($signed(twiddle_factor_table_37_real) + $signed(twiddle_factor_table_37_imag));
  assign _zz_8920 = ($signed(_zz_833) - $signed(_zz_8921));
  assign _zz_8921 = ($signed(_zz_8922) * $signed(twiddle_factor_table_37_imag));
  assign _zz_8922 = ($signed(data_mid_5_38_real) + $signed(data_mid_5_38_imag));
  assign _zz_8923 = fixTo_996_dout;
  assign _zz_8924 = ($signed(_zz_833) + $signed(_zz_8925));
  assign _zz_8925 = ($signed(_zz_8926) * $signed(twiddle_factor_table_37_real));
  assign _zz_8926 = ($signed(data_mid_5_38_imag) - $signed(data_mid_5_38_real));
  assign _zz_8927 = fixTo_997_dout;
  assign _zz_8928 = _zz_8929[35 : 0];
  assign _zz_8929 = _zz_8930;
  assign _zz_8930 = ($signed(_zz_8931) >>> _zz_834);
  assign _zz_8931 = _zz_8932;
  assign _zz_8932 = ($signed(_zz_8934) - $signed(_zz_831));
  assign _zz_8933 = ({9'd0,data_mid_5_6_real} <<< 9);
  assign _zz_8934 = {{9{_zz_8933[26]}}, _zz_8933};
  assign _zz_8935 = fixTo_998_dout;
  assign _zz_8936 = _zz_8937[35 : 0];
  assign _zz_8937 = _zz_8938;
  assign _zz_8938 = ($signed(_zz_8939) >>> _zz_834);
  assign _zz_8939 = _zz_8940;
  assign _zz_8940 = ($signed(_zz_8942) - $signed(_zz_832));
  assign _zz_8941 = ({9'd0,data_mid_5_6_imag} <<< 9);
  assign _zz_8942 = {{9{_zz_8941[26]}}, _zz_8941};
  assign _zz_8943 = fixTo_999_dout;
  assign _zz_8944 = _zz_8945[35 : 0];
  assign _zz_8945 = _zz_8946;
  assign _zz_8946 = ($signed(_zz_8947) >>> _zz_835);
  assign _zz_8947 = _zz_8948;
  assign _zz_8948 = ($signed(_zz_8950) + $signed(_zz_831));
  assign _zz_8949 = ({9'd0,data_mid_5_6_real} <<< 9);
  assign _zz_8950 = {{9{_zz_8949[26]}}, _zz_8949};
  assign _zz_8951 = fixTo_1000_dout;
  assign _zz_8952 = _zz_8953[35 : 0];
  assign _zz_8953 = _zz_8954;
  assign _zz_8954 = ($signed(_zz_8955) >>> _zz_835);
  assign _zz_8955 = _zz_8956;
  assign _zz_8956 = ($signed(_zz_8958) + $signed(_zz_832));
  assign _zz_8957 = ({9'd0,data_mid_5_6_imag} <<< 9);
  assign _zz_8958 = {{9{_zz_8957[26]}}, _zz_8957};
  assign _zz_8959 = fixTo_1001_dout;
  assign _zz_8960 = ($signed(twiddle_factor_table_38_real) + $signed(twiddle_factor_table_38_imag));
  assign _zz_8961 = ($signed(_zz_838) - $signed(_zz_8962));
  assign _zz_8962 = ($signed(_zz_8963) * $signed(twiddle_factor_table_38_imag));
  assign _zz_8963 = ($signed(data_mid_5_39_real) + $signed(data_mid_5_39_imag));
  assign _zz_8964 = fixTo_1002_dout;
  assign _zz_8965 = ($signed(_zz_838) + $signed(_zz_8966));
  assign _zz_8966 = ($signed(_zz_8967) * $signed(twiddle_factor_table_38_real));
  assign _zz_8967 = ($signed(data_mid_5_39_imag) - $signed(data_mid_5_39_real));
  assign _zz_8968 = fixTo_1003_dout;
  assign _zz_8969 = _zz_8970[35 : 0];
  assign _zz_8970 = _zz_8971;
  assign _zz_8971 = ($signed(_zz_8972) >>> _zz_839);
  assign _zz_8972 = _zz_8973;
  assign _zz_8973 = ($signed(_zz_8975) - $signed(_zz_836));
  assign _zz_8974 = ({9'd0,data_mid_5_7_real} <<< 9);
  assign _zz_8975 = {{9{_zz_8974[26]}}, _zz_8974};
  assign _zz_8976 = fixTo_1004_dout;
  assign _zz_8977 = _zz_8978[35 : 0];
  assign _zz_8978 = _zz_8979;
  assign _zz_8979 = ($signed(_zz_8980) >>> _zz_839);
  assign _zz_8980 = _zz_8981;
  assign _zz_8981 = ($signed(_zz_8983) - $signed(_zz_837));
  assign _zz_8982 = ({9'd0,data_mid_5_7_imag} <<< 9);
  assign _zz_8983 = {{9{_zz_8982[26]}}, _zz_8982};
  assign _zz_8984 = fixTo_1005_dout;
  assign _zz_8985 = _zz_8986[35 : 0];
  assign _zz_8986 = _zz_8987;
  assign _zz_8987 = ($signed(_zz_8988) >>> _zz_840);
  assign _zz_8988 = _zz_8989;
  assign _zz_8989 = ($signed(_zz_8991) + $signed(_zz_836));
  assign _zz_8990 = ({9'd0,data_mid_5_7_real} <<< 9);
  assign _zz_8991 = {{9{_zz_8990[26]}}, _zz_8990};
  assign _zz_8992 = fixTo_1006_dout;
  assign _zz_8993 = _zz_8994[35 : 0];
  assign _zz_8994 = _zz_8995;
  assign _zz_8995 = ($signed(_zz_8996) >>> _zz_840);
  assign _zz_8996 = _zz_8997;
  assign _zz_8997 = ($signed(_zz_8999) + $signed(_zz_837));
  assign _zz_8998 = ({9'd0,data_mid_5_7_imag} <<< 9);
  assign _zz_8999 = {{9{_zz_8998[26]}}, _zz_8998};
  assign _zz_9000 = fixTo_1007_dout;
  assign _zz_9001 = ($signed(twiddle_factor_table_39_real) + $signed(twiddle_factor_table_39_imag));
  assign _zz_9002 = ($signed(_zz_843) - $signed(_zz_9003));
  assign _zz_9003 = ($signed(_zz_9004) * $signed(twiddle_factor_table_39_imag));
  assign _zz_9004 = ($signed(data_mid_5_40_real) + $signed(data_mid_5_40_imag));
  assign _zz_9005 = fixTo_1008_dout;
  assign _zz_9006 = ($signed(_zz_843) + $signed(_zz_9007));
  assign _zz_9007 = ($signed(_zz_9008) * $signed(twiddle_factor_table_39_real));
  assign _zz_9008 = ($signed(data_mid_5_40_imag) - $signed(data_mid_5_40_real));
  assign _zz_9009 = fixTo_1009_dout;
  assign _zz_9010 = _zz_9011[35 : 0];
  assign _zz_9011 = _zz_9012;
  assign _zz_9012 = ($signed(_zz_9013) >>> _zz_844);
  assign _zz_9013 = _zz_9014;
  assign _zz_9014 = ($signed(_zz_9016) - $signed(_zz_841));
  assign _zz_9015 = ({9'd0,data_mid_5_8_real} <<< 9);
  assign _zz_9016 = {{9{_zz_9015[26]}}, _zz_9015};
  assign _zz_9017 = fixTo_1010_dout;
  assign _zz_9018 = _zz_9019[35 : 0];
  assign _zz_9019 = _zz_9020;
  assign _zz_9020 = ($signed(_zz_9021) >>> _zz_844);
  assign _zz_9021 = _zz_9022;
  assign _zz_9022 = ($signed(_zz_9024) - $signed(_zz_842));
  assign _zz_9023 = ({9'd0,data_mid_5_8_imag} <<< 9);
  assign _zz_9024 = {{9{_zz_9023[26]}}, _zz_9023};
  assign _zz_9025 = fixTo_1011_dout;
  assign _zz_9026 = _zz_9027[35 : 0];
  assign _zz_9027 = _zz_9028;
  assign _zz_9028 = ($signed(_zz_9029) >>> _zz_845);
  assign _zz_9029 = _zz_9030;
  assign _zz_9030 = ($signed(_zz_9032) + $signed(_zz_841));
  assign _zz_9031 = ({9'd0,data_mid_5_8_real} <<< 9);
  assign _zz_9032 = {{9{_zz_9031[26]}}, _zz_9031};
  assign _zz_9033 = fixTo_1012_dout;
  assign _zz_9034 = _zz_9035[35 : 0];
  assign _zz_9035 = _zz_9036;
  assign _zz_9036 = ($signed(_zz_9037) >>> _zz_845);
  assign _zz_9037 = _zz_9038;
  assign _zz_9038 = ($signed(_zz_9040) + $signed(_zz_842));
  assign _zz_9039 = ({9'd0,data_mid_5_8_imag} <<< 9);
  assign _zz_9040 = {{9{_zz_9039[26]}}, _zz_9039};
  assign _zz_9041 = fixTo_1013_dout;
  assign _zz_9042 = ($signed(twiddle_factor_table_40_real) + $signed(twiddle_factor_table_40_imag));
  assign _zz_9043 = ($signed(_zz_848) - $signed(_zz_9044));
  assign _zz_9044 = ($signed(_zz_9045) * $signed(twiddle_factor_table_40_imag));
  assign _zz_9045 = ($signed(data_mid_5_41_real) + $signed(data_mid_5_41_imag));
  assign _zz_9046 = fixTo_1014_dout;
  assign _zz_9047 = ($signed(_zz_848) + $signed(_zz_9048));
  assign _zz_9048 = ($signed(_zz_9049) * $signed(twiddle_factor_table_40_real));
  assign _zz_9049 = ($signed(data_mid_5_41_imag) - $signed(data_mid_5_41_real));
  assign _zz_9050 = fixTo_1015_dout;
  assign _zz_9051 = _zz_9052[35 : 0];
  assign _zz_9052 = _zz_9053;
  assign _zz_9053 = ($signed(_zz_9054) >>> _zz_849);
  assign _zz_9054 = _zz_9055;
  assign _zz_9055 = ($signed(_zz_9057) - $signed(_zz_846));
  assign _zz_9056 = ({9'd0,data_mid_5_9_real} <<< 9);
  assign _zz_9057 = {{9{_zz_9056[26]}}, _zz_9056};
  assign _zz_9058 = fixTo_1016_dout;
  assign _zz_9059 = _zz_9060[35 : 0];
  assign _zz_9060 = _zz_9061;
  assign _zz_9061 = ($signed(_zz_9062) >>> _zz_849);
  assign _zz_9062 = _zz_9063;
  assign _zz_9063 = ($signed(_zz_9065) - $signed(_zz_847));
  assign _zz_9064 = ({9'd0,data_mid_5_9_imag} <<< 9);
  assign _zz_9065 = {{9{_zz_9064[26]}}, _zz_9064};
  assign _zz_9066 = fixTo_1017_dout;
  assign _zz_9067 = _zz_9068[35 : 0];
  assign _zz_9068 = _zz_9069;
  assign _zz_9069 = ($signed(_zz_9070) >>> _zz_850);
  assign _zz_9070 = _zz_9071;
  assign _zz_9071 = ($signed(_zz_9073) + $signed(_zz_846));
  assign _zz_9072 = ({9'd0,data_mid_5_9_real} <<< 9);
  assign _zz_9073 = {{9{_zz_9072[26]}}, _zz_9072};
  assign _zz_9074 = fixTo_1018_dout;
  assign _zz_9075 = _zz_9076[35 : 0];
  assign _zz_9076 = _zz_9077;
  assign _zz_9077 = ($signed(_zz_9078) >>> _zz_850);
  assign _zz_9078 = _zz_9079;
  assign _zz_9079 = ($signed(_zz_9081) + $signed(_zz_847));
  assign _zz_9080 = ({9'd0,data_mid_5_9_imag} <<< 9);
  assign _zz_9081 = {{9{_zz_9080[26]}}, _zz_9080};
  assign _zz_9082 = fixTo_1019_dout;
  assign _zz_9083 = ($signed(twiddle_factor_table_41_real) + $signed(twiddle_factor_table_41_imag));
  assign _zz_9084 = ($signed(_zz_853) - $signed(_zz_9085));
  assign _zz_9085 = ($signed(_zz_9086) * $signed(twiddle_factor_table_41_imag));
  assign _zz_9086 = ($signed(data_mid_5_42_real) + $signed(data_mid_5_42_imag));
  assign _zz_9087 = fixTo_1020_dout;
  assign _zz_9088 = ($signed(_zz_853) + $signed(_zz_9089));
  assign _zz_9089 = ($signed(_zz_9090) * $signed(twiddle_factor_table_41_real));
  assign _zz_9090 = ($signed(data_mid_5_42_imag) - $signed(data_mid_5_42_real));
  assign _zz_9091 = fixTo_1021_dout;
  assign _zz_9092 = _zz_9093[35 : 0];
  assign _zz_9093 = _zz_9094;
  assign _zz_9094 = ($signed(_zz_9095) >>> _zz_854);
  assign _zz_9095 = _zz_9096;
  assign _zz_9096 = ($signed(_zz_9098) - $signed(_zz_851));
  assign _zz_9097 = ({9'd0,data_mid_5_10_real} <<< 9);
  assign _zz_9098 = {{9{_zz_9097[26]}}, _zz_9097};
  assign _zz_9099 = fixTo_1022_dout;
  assign _zz_9100 = _zz_9101[35 : 0];
  assign _zz_9101 = _zz_9102;
  assign _zz_9102 = ($signed(_zz_9103) >>> _zz_854);
  assign _zz_9103 = _zz_9104;
  assign _zz_9104 = ($signed(_zz_9106) - $signed(_zz_852));
  assign _zz_9105 = ({9'd0,data_mid_5_10_imag} <<< 9);
  assign _zz_9106 = {{9{_zz_9105[26]}}, _zz_9105};
  assign _zz_9107 = fixTo_1023_dout;
  assign _zz_9108 = _zz_9109[35 : 0];
  assign _zz_9109 = _zz_9110;
  assign _zz_9110 = ($signed(_zz_9111) >>> _zz_855);
  assign _zz_9111 = _zz_9112;
  assign _zz_9112 = ($signed(_zz_9114) + $signed(_zz_851));
  assign _zz_9113 = ({9'd0,data_mid_5_10_real} <<< 9);
  assign _zz_9114 = {{9{_zz_9113[26]}}, _zz_9113};
  assign _zz_9115 = fixTo_1024_dout;
  assign _zz_9116 = _zz_9117[35 : 0];
  assign _zz_9117 = _zz_9118;
  assign _zz_9118 = ($signed(_zz_9119) >>> _zz_855);
  assign _zz_9119 = _zz_9120;
  assign _zz_9120 = ($signed(_zz_9122) + $signed(_zz_852));
  assign _zz_9121 = ({9'd0,data_mid_5_10_imag} <<< 9);
  assign _zz_9122 = {{9{_zz_9121[26]}}, _zz_9121};
  assign _zz_9123 = fixTo_1025_dout;
  assign _zz_9124 = ($signed(twiddle_factor_table_42_real) + $signed(twiddle_factor_table_42_imag));
  assign _zz_9125 = ($signed(_zz_858) - $signed(_zz_9126));
  assign _zz_9126 = ($signed(_zz_9127) * $signed(twiddle_factor_table_42_imag));
  assign _zz_9127 = ($signed(data_mid_5_43_real) + $signed(data_mid_5_43_imag));
  assign _zz_9128 = fixTo_1026_dout;
  assign _zz_9129 = ($signed(_zz_858) + $signed(_zz_9130));
  assign _zz_9130 = ($signed(_zz_9131) * $signed(twiddle_factor_table_42_real));
  assign _zz_9131 = ($signed(data_mid_5_43_imag) - $signed(data_mid_5_43_real));
  assign _zz_9132 = fixTo_1027_dout;
  assign _zz_9133 = _zz_9134[35 : 0];
  assign _zz_9134 = _zz_9135;
  assign _zz_9135 = ($signed(_zz_9136) >>> _zz_859);
  assign _zz_9136 = _zz_9137;
  assign _zz_9137 = ($signed(_zz_9139) - $signed(_zz_856));
  assign _zz_9138 = ({9'd0,data_mid_5_11_real} <<< 9);
  assign _zz_9139 = {{9{_zz_9138[26]}}, _zz_9138};
  assign _zz_9140 = fixTo_1028_dout;
  assign _zz_9141 = _zz_9142[35 : 0];
  assign _zz_9142 = _zz_9143;
  assign _zz_9143 = ($signed(_zz_9144) >>> _zz_859);
  assign _zz_9144 = _zz_9145;
  assign _zz_9145 = ($signed(_zz_9147) - $signed(_zz_857));
  assign _zz_9146 = ({9'd0,data_mid_5_11_imag} <<< 9);
  assign _zz_9147 = {{9{_zz_9146[26]}}, _zz_9146};
  assign _zz_9148 = fixTo_1029_dout;
  assign _zz_9149 = _zz_9150[35 : 0];
  assign _zz_9150 = _zz_9151;
  assign _zz_9151 = ($signed(_zz_9152) >>> _zz_860);
  assign _zz_9152 = _zz_9153;
  assign _zz_9153 = ($signed(_zz_9155) + $signed(_zz_856));
  assign _zz_9154 = ({9'd0,data_mid_5_11_real} <<< 9);
  assign _zz_9155 = {{9{_zz_9154[26]}}, _zz_9154};
  assign _zz_9156 = fixTo_1030_dout;
  assign _zz_9157 = _zz_9158[35 : 0];
  assign _zz_9158 = _zz_9159;
  assign _zz_9159 = ($signed(_zz_9160) >>> _zz_860);
  assign _zz_9160 = _zz_9161;
  assign _zz_9161 = ($signed(_zz_9163) + $signed(_zz_857));
  assign _zz_9162 = ({9'd0,data_mid_5_11_imag} <<< 9);
  assign _zz_9163 = {{9{_zz_9162[26]}}, _zz_9162};
  assign _zz_9164 = fixTo_1031_dout;
  assign _zz_9165 = ($signed(twiddle_factor_table_43_real) + $signed(twiddle_factor_table_43_imag));
  assign _zz_9166 = ($signed(_zz_863) - $signed(_zz_9167));
  assign _zz_9167 = ($signed(_zz_9168) * $signed(twiddle_factor_table_43_imag));
  assign _zz_9168 = ($signed(data_mid_5_44_real) + $signed(data_mid_5_44_imag));
  assign _zz_9169 = fixTo_1032_dout;
  assign _zz_9170 = ($signed(_zz_863) + $signed(_zz_9171));
  assign _zz_9171 = ($signed(_zz_9172) * $signed(twiddle_factor_table_43_real));
  assign _zz_9172 = ($signed(data_mid_5_44_imag) - $signed(data_mid_5_44_real));
  assign _zz_9173 = fixTo_1033_dout;
  assign _zz_9174 = _zz_9175[35 : 0];
  assign _zz_9175 = _zz_9176;
  assign _zz_9176 = ($signed(_zz_9177) >>> _zz_864);
  assign _zz_9177 = _zz_9178;
  assign _zz_9178 = ($signed(_zz_9180) - $signed(_zz_861));
  assign _zz_9179 = ({9'd0,data_mid_5_12_real} <<< 9);
  assign _zz_9180 = {{9{_zz_9179[26]}}, _zz_9179};
  assign _zz_9181 = fixTo_1034_dout;
  assign _zz_9182 = _zz_9183[35 : 0];
  assign _zz_9183 = _zz_9184;
  assign _zz_9184 = ($signed(_zz_9185) >>> _zz_864);
  assign _zz_9185 = _zz_9186;
  assign _zz_9186 = ($signed(_zz_9188) - $signed(_zz_862));
  assign _zz_9187 = ({9'd0,data_mid_5_12_imag} <<< 9);
  assign _zz_9188 = {{9{_zz_9187[26]}}, _zz_9187};
  assign _zz_9189 = fixTo_1035_dout;
  assign _zz_9190 = _zz_9191[35 : 0];
  assign _zz_9191 = _zz_9192;
  assign _zz_9192 = ($signed(_zz_9193) >>> _zz_865);
  assign _zz_9193 = _zz_9194;
  assign _zz_9194 = ($signed(_zz_9196) + $signed(_zz_861));
  assign _zz_9195 = ({9'd0,data_mid_5_12_real} <<< 9);
  assign _zz_9196 = {{9{_zz_9195[26]}}, _zz_9195};
  assign _zz_9197 = fixTo_1036_dout;
  assign _zz_9198 = _zz_9199[35 : 0];
  assign _zz_9199 = _zz_9200;
  assign _zz_9200 = ($signed(_zz_9201) >>> _zz_865);
  assign _zz_9201 = _zz_9202;
  assign _zz_9202 = ($signed(_zz_9204) + $signed(_zz_862));
  assign _zz_9203 = ({9'd0,data_mid_5_12_imag} <<< 9);
  assign _zz_9204 = {{9{_zz_9203[26]}}, _zz_9203};
  assign _zz_9205 = fixTo_1037_dout;
  assign _zz_9206 = ($signed(twiddle_factor_table_44_real) + $signed(twiddle_factor_table_44_imag));
  assign _zz_9207 = ($signed(_zz_868) - $signed(_zz_9208));
  assign _zz_9208 = ($signed(_zz_9209) * $signed(twiddle_factor_table_44_imag));
  assign _zz_9209 = ($signed(data_mid_5_45_real) + $signed(data_mid_5_45_imag));
  assign _zz_9210 = fixTo_1038_dout;
  assign _zz_9211 = ($signed(_zz_868) + $signed(_zz_9212));
  assign _zz_9212 = ($signed(_zz_9213) * $signed(twiddle_factor_table_44_real));
  assign _zz_9213 = ($signed(data_mid_5_45_imag) - $signed(data_mid_5_45_real));
  assign _zz_9214 = fixTo_1039_dout;
  assign _zz_9215 = _zz_9216[35 : 0];
  assign _zz_9216 = _zz_9217;
  assign _zz_9217 = ($signed(_zz_9218) >>> _zz_869);
  assign _zz_9218 = _zz_9219;
  assign _zz_9219 = ($signed(_zz_9221) - $signed(_zz_866));
  assign _zz_9220 = ({9'd0,data_mid_5_13_real} <<< 9);
  assign _zz_9221 = {{9{_zz_9220[26]}}, _zz_9220};
  assign _zz_9222 = fixTo_1040_dout;
  assign _zz_9223 = _zz_9224[35 : 0];
  assign _zz_9224 = _zz_9225;
  assign _zz_9225 = ($signed(_zz_9226) >>> _zz_869);
  assign _zz_9226 = _zz_9227;
  assign _zz_9227 = ($signed(_zz_9229) - $signed(_zz_867));
  assign _zz_9228 = ({9'd0,data_mid_5_13_imag} <<< 9);
  assign _zz_9229 = {{9{_zz_9228[26]}}, _zz_9228};
  assign _zz_9230 = fixTo_1041_dout;
  assign _zz_9231 = _zz_9232[35 : 0];
  assign _zz_9232 = _zz_9233;
  assign _zz_9233 = ($signed(_zz_9234) >>> _zz_870);
  assign _zz_9234 = _zz_9235;
  assign _zz_9235 = ($signed(_zz_9237) + $signed(_zz_866));
  assign _zz_9236 = ({9'd0,data_mid_5_13_real} <<< 9);
  assign _zz_9237 = {{9{_zz_9236[26]}}, _zz_9236};
  assign _zz_9238 = fixTo_1042_dout;
  assign _zz_9239 = _zz_9240[35 : 0];
  assign _zz_9240 = _zz_9241;
  assign _zz_9241 = ($signed(_zz_9242) >>> _zz_870);
  assign _zz_9242 = _zz_9243;
  assign _zz_9243 = ($signed(_zz_9245) + $signed(_zz_867));
  assign _zz_9244 = ({9'd0,data_mid_5_13_imag} <<< 9);
  assign _zz_9245 = {{9{_zz_9244[26]}}, _zz_9244};
  assign _zz_9246 = fixTo_1043_dout;
  assign _zz_9247 = ($signed(twiddle_factor_table_45_real) + $signed(twiddle_factor_table_45_imag));
  assign _zz_9248 = ($signed(_zz_873) - $signed(_zz_9249));
  assign _zz_9249 = ($signed(_zz_9250) * $signed(twiddle_factor_table_45_imag));
  assign _zz_9250 = ($signed(data_mid_5_46_real) + $signed(data_mid_5_46_imag));
  assign _zz_9251 = fixTo_1044_dout;
  assign _zz_9252 = ($signed(_zz_873) + $signed(_zz_9253));
  assign _zz_9253 = ($signed(_zz_9254) * $signed(twiddle_factor_table_45_real));
  assign _zz_9254 = ($signed(data_mid_5_46_imag) - $signed(data_mid_5_46_real));
  assign _zz_9255 = fixTo_1045_dout;
  assign _zz_9256 = _zz_9257[35 : 0];
  assign _zz_9257 = _zz_9258;
  assign _zz_9258 = ($signed(_zz_9259) >>> _zz_874);
  assign _zz_9259 = _zz_9260;
  assign _zz_9260 = ($signed(_zz_9262) - $signed(_zz_871));
  assign _zz_9261 = ({9'd0,data_mid_5_14_real} <<< 9);
  assign _zz_9262 = {{9{_zz_9261[26]}}, _zz_9261};
  assign _zz_9263 = fixTo_1046_dout;
  assign _zz_9264 = _zz_9265[35 : 0];
  assign _zz_9265 = _zz_9266;
  assign _zz_9266 = ($signed(_zz_9267) >>> _zz_874);
  assign _zz_9267 = _zz_9268;
  assign _zz_9268 = ($signed(_zz_9270) - $signed(_zz_872));
  assign _zz_9269 = ({9'd0,data_mid_5_14_imag} <<< 9);
  assign _zz_9270 = {{9{_zz_9269[26]}}, _zz_9269};
  assign _zz_9271 = fixTo_1047_dout;
  assign _zz_9272 = _zz_9273[35 : 0];
  assign _zz_9273 = _zz_9274;
  assign _zz_9274 = ($signed(_zz_9275) >>> _zz_875);
  assign _zz_9275 = _zz_9276;
  assign _zz_9276 = ($signed(_zz_9278) + $signed(_zz_871));
  assign _zz_9277 = ({9'd0,data_mid_5_14_real} <<< 9);
  assign _zz_9278 = {{9{_zz_9277[26]}}, _zz_9277};
  assign _zz_9279 = fixTo_1048_dout;
  assign _zz_9280 = _zz_9281[35 : 0];
  assign _zz_9281 = _zz_9282;
  assign _zz_9282 = ($signed(_zz_9283) >>> _zz_875);
  assign _zz_9283 = _zz_9284;
  assign _zz_9284 = ($signed(_zz_9286) + $signed(_zz_872));
  assign _zz_9285 = ({9'd0,data_mid_5_14_imag} <<< 9);
  assign _zz_9286 = {{9{_zz_9285[26]}}, _zz_9285};
  assign _zz_9287 = fixTo_1049_dout;
  assign _zz_9288 = ($signed(twiddle_factor_table_46_real) + $signed(twiddle_factor_table_46_imag));
  assign _zz_9289 = ($signed(_zz_878) - $signed(_zz_9290));
  assign _zz_9290 = ($signed(_zz_9291) * $signed(twiddle_factor_table_46_imag));
  assign _zz_9291 = ($signed(data_mid_5_47_real) + $signed(data_mid_5_47_imag));
  assign _zz_9292 = fixTo_1050_dout;
  assign _zz_9293 = ($signed(_zz_878) + $signed(_zz_9294));
  assign _zz_9294 = ($signed(_zz_9295) * $signed(twiddle_factor_table_46_real));
  assign _zz_9295 = ($signed(data_mid_5_47_imag) - $signed(data_mid_5_47_real));
  assign _zz_9296 = fixTo_1051_dout;
  assign _zz_9297 = _zz_9298[35 : 0];
  assign _zz_9298 = _zz_9299;
  assign _zz_9299 = ($signed(_zz_9300) >>> _zz_879);
  assign _zz_9300 = _zz_9301;
  assign _zz_9301 = ($signed(_zz_9303) - $signed(_zz_876));
  assign _zz_9302 = ({9'd0,data_mid_5_15_real} <<< 9);
  assign _zz_9303 = {{9{_zz_9302[26]}}, _zz_9302};
  assign _zz_9304 = fixTo_1052_dout;
  assign _zz_9305 = _zz_9306[35 : 0];
  assign _zz_9306 = _zz_9307;
  assign _zz_9307 = ($signed(_zz_9308) >>> _zz_879);
  assign _zz_9308 = _zz_9309;
  assign _zz_9309 = ($signed(_zz_9311) - $signed(_zz_877));
  assign _zz_9310 = ({9'd0,data_mid_5_15_imag} <<< 9);
  assign _zz_9311 = {{9{_zz_9310[26]}}, _zz_9310};
  assign _zz_9312 = fixTo_1053_dout;
  assign _zz_9313 = _zz_9314[35 : 0];
  assign _zz_9314 = _zz_9315;
  assign _zz_9315 = ($signed(_zz_9316) >>> _zz_880);
  assign _zz_9316 = _zz_9317;
  assign _zz_9317 = ($signed(_zz_9319) + $signed(_zz_876));
  assign _zz_9318 = ({9'd0,data_mid_5_15_real} <<< 9);
  assign _zz_9319 = {{9{_zz_9318[26]}}, _zz_9318};
  assign _zz_9320 = fixTo_1054_dout;
  assign _zz_9321 = _zz_9322[35 : 0];
  assign _zz_9322 = _zz_9323;
  assign _zz_9323 = ($signed(_zz_9324) >>> _zz_880);
  assign _zz_9324 = _zz_9325;
  assign _zz_9325 = ($signed(_zz_9327) + $signed(_zz_877));
  assign _zz_9326 = ({9'd0,data_mid_5_15_imag} <<< 9);
  assign _zz_9327 = {{9{_zz_9326[26]}}, _zz_9326};
  assign _zz_9328 = fixTo_1055_dout;
  assign _zz_9329 = ($signed(twiddle_factor_table_47_real) + $signed(twiddle_factor_table_47_imag));
  assign _zz_9330 = ($signed(_zz_883) - $signed(_zz_9331));
  assign _zz_9331 = ($signed(_zz_9332) * $signed(twiddle_factor_table_47_imag));
  assign _zz_9332 = ($signed(data_mid_5_48_real) + $signed(data_mid_5_48_imag));
  assign _zz_9333 = fixTo_1056_dout;
  assign _zz_9334 = ($signed(_zz_883) + $signed(_zz_9335));
  assign _zz_9335 = ($signed(_zz_9336) * $signed(twiddle_factor_table_47_real));
  assign _zz_9336 = ($signed(data_mid_5_48_imag) - $signed(data_mid_5_48_real));
  assign _zz_9337 = fixTo_1057_dout;
  assign _zz_9338 = _zz_9339[35 : 0];
  assign _zz_9339 = _zz_9340;
  assign _zz_9340 = ($signed(_zz_9341) >>> _zz_884);
  assign _zz_9341 = _zz_9342;
  assign _zz_9342 = ($signed(_zz_9344) - $signed(_zz_881));
  assign _zz_9343 = ({9'd0,data_mid_5_16_real} <<< 9);
  assign _zz_9344 = {{9{_zz_9343[26]}}, _zz_9343};
  assign _zz_9345 = fixTo_1058_dout;
  assign _zz_9346 = _zz_9347[35 : 0];
  assign _zz_9347 = _zz_9348;
  assign _zz_9348 = ($signed(_zz_9349) >>> _zz_884);
  assign _zz_9349 = _zz_9350;
  assign _zz_9350 = ($signed(_zz_9352) - $signed(_zz_882));
  assign _zz_9351 = ({9'd0,data_mid_5_16_imag} <<< 9);
  assign _zz_9352 = {{9{_zz_9351[26]}}, _zz_9351};
  assign _zz_9353 = fixTo_1059_dout;
  assign _zz_9354 = _zz_9355[35 : 0];
  assign _zz_9355 = _zz_9356;
  assign _zz_9356 = ($signed(_zz_9357) >>> _zz_885);
  assign _zz_9357 = _zz_9358;
  assign _zz_9358 = ($signed(_zz_9360) + $signed(_zz_881));
  assign _zz_9359 = ({9'd0,data_mid_5_16_real} <<< 9);
  assign _zz_9360 = {{9{_zz_9359[26]}}, _zz_9359};
  assign _zz_9361 = fixTo_1060_dout;
  assign _zz_9362 = _zz_9363[35 : 0];
  assign _zz_9363 = _zz_9364;
  assign _zz_9364 = ($signed(_zz_9365) >>> _zz_885);
  assign _zz_9365 = _zz_9366;
  assign _zz_9366 = ($signed(_zz_9368) + $signed(_zz_882));
  assign _zz_9367 = ({9'd0,data_mid_5_16_imag} <<< 9);
  assign _zz_9368 = {{9{_zz_9367[26]}}, _zz_9367};
  assign _zz_9369 = fixTo_1061_dout;
  assign _zz_9370 = ($signed(twiddle_factor_table_48_real) + $signed(twiddle_factor_table_48_imag));
  assign _zz_9371 = ($signed(_zz_888) - $signed(_zz_9372));
  assign _zz_9372 = ($signed(_zz_9373) * $signed(twiddle_factor_table_48_imag));
  assign _zz_9373 = ($signed(data_mid_5_49_real) + $signed(data_mid_5_49_imag));
  assign _zz_9374 = fixTo_1062_dout;
  assign _zz_9375 = ($signed(_zz_888) + $signed(_zz_9376));
  assign _zz_9376 = ($signed(_zz_9377) * $signed(twiddle_factor_table_48_real));
  assign _zz_9377 = ($signed(data_mid_5_49_imag) - $signed(data_mid_5_49_real));
  assign _zz_9378 = fixTo_1063_dout;
  assign _zz_9379 = _zz_9380[35 : 0];
  assign _zz_9380 = _zz_9381;
  assign _zz_9381 = ($signed(_zz_9382) >>> _zz_889);
  assign _zz_9382 = _zz_9383;
  assign _zz_9383 = ($signed(_zz_9385) - $signed(_zz_886));
  assign _zz_9384 = ({9'd0,data_mid_5_17_real} <<< 9);
  assign _zz_9385 = {{9{_zz_9384[26]}}, _zz_9384};
  assign _zz_9386 = fixTo_1064_dout;
  assign _zz_9387 = _zz_9388[35 : 0];
  assign _zz_9388 = _zz_9389;
  assign _zz_9389 = ($signed(_zz_9390) >>> _zz_889);
  assign _zz_9390 = _zz_9391;
  assign _zz_9391 = ($signed(_zz_9393) - $signed(_zz_887));
  assign _zz_9392 = ({9'd0,data_mid_5_17_imag} <<< 9);
  assign _zz_9393 = {{9{_zz_9392[26]}}, _zz_9392};
  assign _zz_9394 = fixTo_1065_dout;
  assign _zz_9395 = _zz_9396[35 : 0];
  assign _zz_9396 = _zz_9397;
  assign _zz_9397 = ($signed(_zz_9398) >>> _zz_890);
  assign _zz_9398 = _zz_9399;
  assign _zz_9399 = ($signed(_zz_9401) + $signed(_zz_886));
  assign _zz_9400 = ({9'd0,data_mid_5_17_real} <<< 9);
  assign _zz_9401 = {{9{_zz_9400[26]}}, _zz_9400};
  assign _zz_9402 = fixTo_1066_dout;
  assign _zz_9403 = _zz_9404[35 : 0];
  assign _zz_9404 = _zz_9405;
  assign _zz_9405 = ($signed(_zz_9406) >>> _zz_890);
  assign _zz_9406 = _zz_9407;
  assign _zz_9407 = ($signed(_zz_9409) + $signed(_zz_887));
  assign _zz_9408 = ({9'd0,data_mid_5_17_imag} <<< 9);
  assign _zz_9409 = {{9{_zz_9408[26]}}, _zz_9408};
  assign _zz_9410 = fixTo_1067_dout;
  assign _zz_9411 = ($signed(twiddle_factor_table_49_real) + $signed(twiddle_factor_table_49_imag));
  assign _zz_9412 = ($signed(_zz_893) - $signed(_zz_9413));
  assign _zz_9413 = ($signed(_zz_9414) * $signed(twiddle_factor_table_49_imag));
  assign _zz_9414 = ($signed(data_mid_5_50_real) + $signed(data_mid_5_50_imag));
  assign _zz_9415 = fixTo_1068_dout;
  assign _zz_9416 = ($signed(_zz_893) + $signed(_zz_9417));
  assign _zz_9417 = ($signed(_zz_9418) * $signed(twiddle_factor_table_49_real));
  assign _zz_9418 = ($signed(data_mid_5_50_imag) - $signed(data_mid_5_50_real));
  assign _zz_9419 = fixTo_1069_dout;
  assign _zz_9420 = _zz_9421[35 : 0];
  assign _zz_9421 = _zz_9422;
  assign _zz_9422 = ($signed(_zz_9423) >>> _zz_894);
  assign _zz_9423 = _zz_9424;
  assign _zz_9424 = ($signed(_zz_9426) - $signed(_zz_891));
  assign _zz_9425 = ({9'd0,data_mid_5_18_real} <<< 9);
  assign _zz_9426 = {{9{_zz_9425[26]}}, _zz_9425};
  assign _zz_9427 = fixTo_1070_dout;
  assign _zz_9428 = _zz_9429[35 : 0];
  assign _zz_9429 = _zz_9430;
  assign _zz_9430 = ($signed(_zz_9431) >>> _zz_894);
  assign _zz_9431 = _zz_9432;
  assign _zz_9432 = ($signed(_zz_9434) - $signed(_zz_892));
  assign _zz_9433 = ({9'd0,data_mid_5_18_imag} <<< 9);
  assign _zz_9434 = {{9{_zz_9433[26]}}, _zz_9433};
  assign _zz_9435 = fixTo_1071_dout;
  assign _zz_9436 = _zz_9437[35 : 0];
  assign _zz_9437 = _zz_9438;
  assign _zz_9438 = ($signed(_zz_9439) >>> _zz_895);
  assign _zz_9439 = _zz_9440;
  assign _zz_9440 = ($signed(_zz_9442) + $signed(_zz_891));
  assign _zz_9441 = ({9'd0,data_mid_5_18_real} <<< 9);
  assign _zz_9442 = {{9{_zz_9441[26]}}, _zz_9441};
  assign _zz_9443 = fixTo_1072_dout;
  assign _zz_9444 = _zz_9445[35 : 0];
  assign _zz_9445 = _zz_9446;
  assign _zz_9446 = ($signed(_zz_9447) >>> _zz_895);
  assign _zz_9447 = _zz_9448;
  assign _zz_9448 = ($signed(_zz_9450) + $signed(_zz_892));
  assign _zz_9449 = ({9'd0,data_mid_5_18_imag} <<< 9);
  assign _zz_9450 = {{9{_zz_9449[26]}}, _zz_9449};
  assign _zz_9451 = fixTo_1073_dout;
  assign _zz_9452 = ($signed(twiddle_factor_table_50_real) + $signed(twiddle_factor_table_50_imag));
  assign _zz_9453 = ($signed(_zz_898) - $signed(_zz_9454));
  assign _zz_9454 = ($signed(_zz_9455) * $signed(twiddle_factor_table_50_imag));
  assign _zz_9455 = ($signed(data_mid_5_51_real) + $signed(data_mid_5_51_imag));
  assign _zz_9456 = fixTo_1074_dout;
  assign _zz_9457 = ($signed(_zz_898) + $signed(_zz_9458));
  assign _zz_9458 = ($signed(_zz_9459) * $signed(twiddle_factor_table_50_real));
  assign _zz_9459 = ($signed(data_mid_5_51_imag) - $signed(data_mid_5_51_real));
  assign _zz_9460 = fixTo_1075_dout;
  assign _zz_9461 = _zz_9462[35 : 0];
  assign _zz_9462 = _zz_9463;
  assign _zz_9463 = ($signed(_zz_9464) >>> _zz_899);
  assign _zz_9464 = _zz_9465;
  assign _zz_9465 = ($signed(_zz_9467) - $signed(_zz_896));
  assign _zz_9466 = ({9'd0,data_mid_5_19_real} <<< 9);
  assign _zz_9467 = {{9{_zz_9466[26]}}, _zz_9466};
  assign _zz_9468 = fixTo_1076_dout;
  assign _zz_9469 = _zz_9470[35 : 0];
  assign _zz_9470 = _zz_9471;
  assign _zz_9471 = ($signed(_zz_9472) >>> _zz_899);
  assign _zz_9472 = _zz_9473;
  assign _zz_9473 = ($signed(_zz_9475) - $signed(_zz_897));
  assign _zz_9474 = ({9'd0,data_mid_5_19_imag} <<< 9);
  assign _zz_9475 = {{9{_zz_9474[26]}}, _zz_9474};
  assign _zz_9476 = fixTo_1077_dout;
  assign _zz_9477 = _zz_9478[35 : 0];
  assign _zz_9478 = _zz_9479;
  assign _zz_9479 = ($signed(_zz_9480) >>> _zz_900);
  assign _zz_9480 = _zz_9481;
  assign _zz_9481 = ($signed(_zz_9483) + $signed(_zz_896));
  assign _zz_9482 = ({9'd0,data_mid_5_19_real} <<< 9);
  assign _zz_9483 = {{9{_zz_9482[26]}}, _zz_9482};
  assign _zz_9484 = fixTo_1078_dout;
  assign _zz_9485 = _zz_9486[35 : 0];
  assign _zz_9486 = _zz_9487;
  assign _zz_9487 = ($signed(_zz_9488) >>> _zz_900);
  assign _zz_9488 = _zz_9489;
  assign _zz_9489 = ($signed(_zz_9491) + $signed(_zz_897));
  assign _zz_9490 = ({9'd0,data_mid_5_19_imag} <<< 9);
  assign _zz_9491 = {{9{_zz_9490[26]}}, _zz_9490};
  assign _zz_9492 = fixTo_1079_dout;
  assign _zz_9493 = ($signed(twiddle_factor_table_51_real) + $signed(twiddle_factor_table_51_imag));
  assign _zz_9494 = ($signed(_zz_903) - $signed(_zz_9495));
  assign _zz_9495 = ($signed(_zz_9496) * $signed(twiddle_factor_table_51_imag));
  assign _zz_9496 = ($signed(data_mid_5_52_real) + $signed(data_mid_5_52_imag));
  assign _zz_9497 = fixTo_1080_dout;
  assign _zz_9498 = ($signed(_zz_903) + $signed(_zz_9499));
  assign _zz_9499 = ($signed(_zz_9500) * $signed(twiddle_factor_table_51_real));
  assign _zz_9500 = ($signed(data_mid_5_52_imag) - $signed(data_mid_5_52_real));
  assign _zz_9501 = fixTo_1081_dout;
  assign _zz_9502 = _zz_9503[35 : 0];
  assign _zz_9503 = _zz_9504;
  assign _zz_9504 = ($signed(_zz_9505) >>> _zz_904);
  assign _zz_9505 = _zz_9506;
  assign _zz_9506 = ($signed(_zz_9508) - $signed(_zz_901));
  assign _zz_9507 = ({9'd0,data_mid_5_20_real} <<< 9);
  assign _zz_9508 = {{9{_zz_9507[26]}}, _zz_9507};
  assign _zz_9509 = fixTo_1082_dout;
  assign _zz_9510 = _zz_9511[35 : 0];
  assign _zz_9511 = _zz_9512;
  assign _zz_9512 = ($signed(_zz_9513) >>> _zz_904);
  assign _zz_9513 = _zz_9514;
  assign _zz_9514 = ($signed(_zz_9516) - $signed(_zz_902));
  assign _zz_9515 = ({9'd0,data_mid_5_20_imag} <<< 9);
  assign _zz_9516 = {{9{_zz_9515[26]}}, _zz_9515};
  assign _zz_9517 = fixTo_1083_dout;
  assign _zz_9518 = _zz_9519[35 : 0];
  assign _zz_9519 = _zz_9520;
  assign _zz_9520 = ($signed(_zz_9521) >>> _zz_905);
  assign _zz_9521 = _zz_9522;
  assign _zz_9522 = ($signed(_zz_9524) + $signed(_zz_901));
  assign _zz_9523 = ({9'd0,data_mid_5_20_real} <<< 9);
  assign _zz_9524 = {{9{_zz_9523[26]}}, _zz_9523};
  assign _zz_9525 = fixTo_1084_dout;
  assign _zz_9526 = _zz_9527[35 : 0];
  assign _zz_9527 = _zz_9528;
  assign _zz_9528 = ($signed(_zz_9529) >>> _zz_905);
  assign _zz_9529 = _zz_9530;
  assign _zz_9530 = ($signed(_zz_9532) + $signed(_zz_902));
  assign _zz_9531 = ({9'd0,data_mid_5_20_imag} <<< 9);
  assign _zz_9532 = {{9{_zz_9531[26]}}, _zz_9531};
  assign _zz_9533 = fixTo_1085_dout;
  assign _zz_9534 = ($signed(twiddle_factor_table_52_real) + $signed(twiddle_factor_table_52_imag));
  assign _zz_9535 = ($signed(_zz_908) - $signed(_zz_9536));
  assign _zz_9536 = ($signed(_zz_9537) * $signed(twiddle_factor_table_52_imag));
  assign _zz_9537 = ($signed(data_mid_5_53_real) + $signed(data_mid_5_53_imag));
  assign _zz_9538 = fixTo_1086_dout;
  assign _zz_9539 = ($signed(_zz_908) + $signed(_zz_9540));
  assign _zz_9540 = ($signed(_zz_9541) * $signed(twiddle_factor_table_52_real));
  assign _zz_9541 = ($signed(data_mid_5_53_imag) - $signed(data_mid_5_53_real));
  assign _zz_9542 = fixTo_1087_dout;
  assign _zz_9543 = _zz_9544[35 : 0];
  assign _zz_9544 = _zz_9545;
  assign _zz_9545 = ($signed(_zz_9546) >>> _zz_909);
  assign _zz_9546 = _zz_9547;
  assign _zz_9547 = ($signed(_zz_9549) - $signed(_zz_906));
  assign _zz_9548 = ({9'd0,data_mid_5_21_real} <<< 9);
  assign _zz_9549 = {{9{_zz_9548[26]}}, _zz_9548};
  assign _zz_9550 = fixTo_1088_dout;
  assign _zz_9551 = _zz_9552[35 : 0];
  assign _zz_9552 = _zz_9553;
  assign _zz_9553 = ($signed(_zz_9554) >>> _zz_909);
  assign _zz_9554 = _zz_9555;
  assign _zz_9555 = ($signed(_zz_9557) - $signed(_zz_907));
  assign _zz_9556 = ({9'd0,data_mid_5_21_imag} <<< 9);
  assign _zz_9557 = {{9{_zz_9556[26]}}, _zz_9556};
  assign _zz_9558 = fixTo_1089_dout;
  assign _zz_9559 = _zz_9560[35 : 0];
  assign _zz_9560 = _zz_9561;
  assign _zz_9561 = ($signed(_zz_9562) >>> _zz_910);
  assign _zz_9562 = _zz_9563;
  assign _zz_9563 = ($signed(_zz_9565) + $signed(_zz_906));
  assign _zz_9564 = ({9'd0,data_mid_5_21_real} <<< 9);
  assign _zz_9565 = {{9{_zz_9564[26]}}, _zz_9564};
  assign _zz_9566 = fixTo_1090_dout;
  assign _zz_9567 = _zz_9568[35 : 0];
  assign _zz_9568 = _zz_9569;
  assign _zz_9569 = ($signed(_zz_9570) >>> _zz_910);
  assign _zz_9570 = _zz_9571;
  assign _zz_9571 = ($signed(_zz_9573) + $signed(_zz_907));
  assign _zz_9572 = ({9'd0,data_mid_5_21_imag} <<< 9);
  assign _zz_9573 = {{9{_zz_9572[26]}}, _zz_9572};
  assign _zz_9574 = fixTo_1091_dout;
  assign _zz_9575 = ($signed(twiddle_factor_table_53_real) + $signed(twiddle_factor_table_53_imag));
  assign _zz_9576 = ($signed(_zz_913) - $signed(_zz_9577));
  assign _zz_9577 = ($signed(_zz_9578) * $signed(twiddle_factor_table_53_imag));
  assign _zz_9578 = ($signed(data_mid_5_54_real) + $signed(data_mid_5_54_imag));
  assign _zz_9579 = fixTo_1092_dout;
  assign _zz_9580 = ($signed(_zz_913) + $signed(_zz_9581));
  assign _zz_9581 = ($signed(_zz_9582) * $signed(twiddle_factor_table_53_real));
  assign _zz_9582 = ($signed(data_mid_5_54_imag) - $signed(data_mid_5_54_real));
  assign _zz_9583 = fixTo_1093_dout;
  assign _zz_9584 = _zz_9585[35 : 0];
  assign _zz_9585 = _zz_9586;
  assign _zz_9586 = ($signed(_zz_9587) >>> _zz_914);
  assign _zz_9587 = _zz_9588;
  assign _zz_9588 = ($signed(_zz_9590) - $signed(_zz_911));
  assign _zz_9589 = ({9'd0,data_mid_5_22_real} <<< 9);
  assign _zz_9590 = {{9{_zz_9589[26]}}, _zz_9589};
  assign _zz_9591 = fixTo_1094_dout;
  assign _zz_9592 = _zz_9593[35 : 0];
  assign _zz_9593 = _zz_9594;
  assign _zz_9594 = ($signed(_zz_9595) >>> _zz_914);
  assign _zz_9595 = _zz_9596;
  assign _zz_9596 = ($signed(_zz_9598) - $signed(_zz_912));
  assign _zz_9597 = ({9'd0,data_mid_5_22_imag} <<< 9);
  assign _zz_9598 = {{9{_zz_9597[26]}}, _zz_9597};
  assign _zz_9599 = fixTo_1095_dout;
  assign _zz_9600 = _zz_9601[35 : 0];
  assign _zz_9601 = _zz_9602;
  assign _zz_9602 = ($signed(_zz_9603) >>> _zz_915);
  assign _zz_9603 = _zz_9604;
  assign _zz_9604 = ($signed(_zz_9606) + $signed(_zz_911));
  assign _zz_9605 = ({9'd0,data_mid_5_22_real} <<< 9);
  assign _zz_9606 = {{9{_zz_9605[26]}}, _zz_9605};
  assign _zz_9607 = fixTo_1096_dout;
  assign _zz_9608 = _zz_9609[35 : 0];
  assign _zz_9609 = _zz_9610;
  assign _zz_9610 = ($signed(_zz_9611) >>> _zz_915);
  assign _zz_9611 = _zz_9612;
  assign _zz_9612 = ($signed(_zz_9614) + $signed(_zz_912));
  assign _zz_9613 = ({9'd0,data_mid_5_22_imag} <<< 9);
  assign _zz_9614 = {{9{_zz_9613[26]}}, _zz_9613};
  assign _zz_9615 = fixTo_1097_dout;
  assign _zz_9616 = ($signed(twiddle_factor_table_54_real) + $signed(twiddle_factor_table_54_imag));
  assign _zz_9617 = ($signed(_zz_918) - $signed(_zz_9618));
  assign _zz_9618 = ($signed(_zz_9619) * $signed(twiddle_factor_table_54_imag));
  assign _zz_9619 = ($signed(data_mid_5_55_real) + $signed(data_mid_5_55_imag));
  assign _zz_9620 = fixTo_1098_dout;
  assign _zz_9621 = ($signed(_zz_918) + $signed(_zz_9622));
  assign _zz_9622 = ($signed(_zz_9623) * $signed(twiddle_factor_table_54_real));
  assign _zz_9623 = ($signed(data_mid_5_55_imag) - $signed(data_mid_5_55_real));
  assign _zz_9624 = fixTo_1099_dout;
  assign _zz_9625 = _zz_9626[35 : 0];
  assign _zz_9626 = _zz_9627;
  assign _zz_9627 = ($signed(_zz_9628) >>> _zz_919);
  assign _zz_9628 = _zz_9629;
  assign _zz_9629 = ($signed(_zz_9631) - $signed(_zz_916));
  assign _zz_9630 = ({9'd0,data_mid_5_23_real} <<< 9);
  assign _zz_9631 = {{9{_zz_9630[26]}}, _zz_9630};
  assign _zz_9632 = fixTo_1100_dout;
  assign _zz_9633 = _zz_9634[35 : 0];
  assign _zz_9634 = _zz_9635;
  assign _zz_9635 = ($signed(_zz_9636) >>> _zz_919);
  assign _zz_9636 = _zz_9637;
  assign _zz_9637 = ($signed(_zz_9639) - $signed(_zz_917));
  assign _zz_9638 = ({9'd0,data_mid_5_23_imag} <<< 9);
  assign _zz_9639 = {{9{_zz_9638[26]}}, _zz_9638};
  assign _zz_9640 = fixTo_1101_dout;
  assign _zz_9641 = _zz_9642[35 : 0];
  assign _zz_9642 = _zz_9643;
  assign _zz_9643 = ($signed(_zz_9644) >>> _zz_920);
  assign _zz_9644 = _zz_9645;
  assign _zz_9645 = ($signed(_zz_9647) + $signed(_zz_916));
  assign _zz_9646 = ({9'd0,data_mid_5_23_real} <<< 9);
  assign _zz_9647 = {{9{_zz_9646[26]}}, _zz_9646};
  assign _zz_9648 = fixTo_1102_dout;
  assign _zz_9649 = _zz_9650[35 : 0];
  assign _zz_9650 = _zz_9651;
  assign _zz_9651 = ($signed(_zz_9652) >>> _zz_920);
  assign _zz_9652 = _zz_9653;
  assign _zz_9653 = ($signed(_zz_9655) + $signed(_zz_917));
  assign _zz_9654 = ({9'd0,data_mid_5_23_imag} <<< 9);
  assign _zz_9655 = {{9{_zz_9654[26]}}, _zz_9654};
  assign _zz_9656 = fixTo_1103_dout;
  assign _zz_9657 = ($signed(twiddle_factor_table_55_real) + $signed(twiddle_factor_table_55_imag));
  assign _zz_9658 = ($signed(_zz_923) - $signed(_zz_9659));
  assign _zz_9659 = ($signed(_zz_9660) * $signed(twiddle_factor_table_55_imag));
  assign _zz_9660 = ($signed(data_mid_5_56_real) + $signed(data_mid_5_56_imag));
  assign _zz_9661 = fixTo_1104_dout;
  assign _zz_9662 = ($signed(_zz_923) + $signed(_zz_9663));
  assign _zz_9663 = ($signed(_zz_9664) * $signed(twiddle_factor_table_55_real));
  assign _zz_9664 = ($signed(data_mid_5_56_imag) - $signed(data_mid_5_56_real));
  assign _zz_9665 = fixTo_1105_dout;
  assign _zz_9666 = _zz_9667[35 : 0];
  assign _zz_9667 = _zz_9668;
  assign _zz_9668 = ($signed(_zz_9669) >>> _zz_924);
  assign _zz_9669 = _zz_9670;
  assign _zz_9670 = ($signed(_zz_9672) - $signed(_zz_921));
  assign _zz_9671 = ({9'd0,data_mid_5_24_real} <<< 9);
  assign _zz_9672 = {{9{_zz_9671[26]}}, _zz_9671};
  assign _zz_9673 = fixTo_1106_dout;
  assign _zz_9674 = _zz_9675[35 : 0];
  assign _zz_9675 = _zz_9676;
  assign _zz_9676 = ($signed(_zz_9677) >>> _zz_924);
  assign _zz_9677 = _zz_9678;
  assign _zz_9678 = ($signed(_zz_9680) - $signed(_zz_922));
  assign _zz_9679 = ({9'd0,data_mid_5_24_imag} <<< 9);
  assign _zz_9680 = {{9{_zz_9679[26]}}, _zz_9679};
  assign _zz_9681 = fixTo_1107_dout;
  assign _zz_9682 = _zz_9683[35 : 0];
  assign _zz_9683 = _zz_9684;
  assign _zz_9684 = ($signed(_zz_9685) >>> _zz_925);
  assign _zz_9685 = _zz_9686;
  assign _zz_9686 = ($signed(_zz_9688) + $signed(_zz_921));
  assign _zz_9687 = ({9'd0,data_mid_5_24_real} <<< 9);
  assign _zz_9688 = {{9{_zz_9687[26]}}, _zz_9687};
  assign _zz_9689 = fixTo_1108_dout;
  assign _zz_9690 = _zz_9691[35 : 0];
  assign _zz_9691 = _zz_9692;
  assign _zz_9692 = ($signed(_zz_9693) >>> _zz_925);
  assign _zz_9693 = _zz_9694;
  assign _zz_9694 = ($signed(_zz_9696) + $signed(_zz_922));
  assign _zz_9695 = ({9'd0,data_mid_5_24_imag} <<< 9);
  assign _zz_9696 = {{9{_zz_9695[26]}}, _zz_9695};
  assign _zz_9697 = fixTo_1109_dout;
  assign _zz_9698 = ($signed(twiddle_factor_table_56_real) + $signed(twiddle_factor_table_56_imag));
  assign _zz_9699 = ($signed(_zz_928) - $signed(_zz_9700));
  assign _zz_9700 = ($signed(_zz_9701) * $signed(twiddle_factor_table_56_imag));
  assign _zz_9701 = ($signed(data_mid_5_57_real) + $signed(data_mid_5_57_imag));
  assign _zz_9702 = fixTo_1110_dout;
  assign _zz_9703 = ($signed(_zz_928) + $signed(_zz_9704));
  assign _zz_9704 = ($signed(_zz_9705) * $signed(twiddle_factor_table_56_real));
  assign _zz_9705 = ($signed(data_mid_5_57_imag) - $signed(data_mid_5_57_real));
  assign _zz_9706 = fixTo_1111_dout;
  assign _zz_9707 = _zz_9708[35 : 0];
  assign _zz_9708 = _zz_9709;
  assign _zz_9709 = ($signed(_zz_9710) >>> _zz_929);
  assign _zz_9710 = _zz_9711;
  assign _zz_9711 = ($signed(_zz_9713) - $signed(_zz_926));
  assign _zz_9712 = ({9'd0,data_mid_5_25_real} <<< 9);
  assign _zz_9713 = {{9{_zz_9712[26]}}, _zz_9712};
  assign _zz_9714 = fixTo_1112_dout;
  assign _zz_9715 = _zz_9716[35 : 0];
  assign _zz_9716 = _zz_9717;
  assign _zz_9717 = ($signed(_zz_9718) >>> _zz_929);
  assign _zz_9718 = _zz_9719;
  assign _zz_9719 = ($signed(_zz_9721) - $signed(_zz_927));
  assign _zz_9720 = ({9'd0,data_mid_5_25_imag} <<< 9);
  assign _zz_9721 = {{9{_zz_9720[26]}}, _zz_9720};
  assign _zz_9722 = fixTo_1113_dout;
  assign _zz_9723 = _zz_9724[35 : 0];
  assign _zz_9724 = _zz_9725;
  assign _zz_9725 = ($signed(_zz_9726) >>> _zz_930);
  assign _zz_9726 = _zz_9727;
  assign _zz_9727 = ($signed(_zz_9729) + $signed(_zz_926));
  assign _zz_9728 = ({9'd0,data_mid_5_25_real} <<< 9);
  assign _zz_9729 = {{9{_zz_9728[26]}}, _zz_9728};
  assign _zz_9730 = fixTo_1114_dout;
  assign _zz_9731 = _zz_9732[35 : 0];
  assign _zz_9732 = _zz_9733;
  assign _zz_9733 = ($signed(_zz_9734) >>> _zz_930);
  assign _zz_9734 = _zz_9735;
  assign _zz_9735 = ($signed(_zz_9737) + $signed(_zz_927));
  assign _zz_9736 = ({9'd0,data_mid_5_25_imag} <<< 9);
  assign _zz_9737 = {{9{_zz_9736[26]}}, _zz_9736};
  assign _zz_9738 = fixTo_1115_dout;
  assign _zz_9739 = ($signed(twiddle_factor_table_57_real) + $signed(twiddle_factor_table_57_imag));
  assign _zz_9740 = ($signed(_zz_933) - $signed(_zz_9741));
  assign _zz_9741 = ($signed(_zz_9742) * $signed(twiddle_factor_table_57_imag));
  assign _zz_9742 = ($signed(data_mid_5_58_real) + $signed(data_mid_5_58_imag));
  assign _zz_9743 = fixTo_1116_dout;
  assign _zz_9744 = ($signed(_zz_933) + $signed(_zz_9745));
  assign _zz_9745 = ($signed(_zz_9746) * $signed(twiddle_factor_table_57_real));
  assign _zz_9746 = ($signed(data_mid_5_58_imag) - $signed(data_mid_5_58_real));
  assign _zz_9747 = fixTo_1117_dout;
  assign _zz_9748 = _zz_9749[35 : 0];
  assign _zz_9749 = _zz_9750;
  assign _zz_9750 = ($signed(_zz_9751) >>> _zz_934);
  assign _zz_9751 = _zz_9752;
  assign _zz_9752 = ($signed(_zz_9754) - $signed(_zz_931));
  assign _zz_9753 = ({9'd0,data_mid_5_26_real} <<< 9);
  assign _zz_9754 = {{9{_zz_9753[26]}}, _zz_9753};
  assign _zz_9755 = fixTo_1118_dout;
  assign _zz_9756 = _zz_9757[35 : 0];
  assign _zz_9757 = _zz_9758;
  assign _zz_9758 = ($signed(_zz_9759) >>> _zz_934);
  assign _zz_9759 = _zz_9760;
  assign _zz_9760 = ($signed(_zz_9762) - $signed(_zz_932));
  assign _zz_9761 = ({9'd0,data_mid_5_26_imag} <<< 9);
  assign _zz_9762 = {{9{_zz_9761[26]}}, _zz_9761};
  assign _zz_9763 = fixTo_1119_dout;
  assign _zz_9764 = _zz_9765[35 : 0];
  assign _zz_9765 = _zz_9766;
  assign _zz_9766 = ($signed(_zz_9767) >>> _zz_935);
  assign _zz_9767 = _zz_9768;
  assign _zz_9768 = ($signed(_zz_9770) + $signed(_zz_931));
  assign _zz_9769 = ({9'd0,data_mid_5_26_real} <<< 9);
  assign _zz_9770 = {{9{_zz_9769[26]}}, _zz_9769};
  assign _zz_9771 = fixTo_1120_dout;
  assign _zz_9772 = _zz_9773[35 : 0];
  assign _zz_9773 = _zz_9774;
  assign _zz_9774 = ($signed(_zz_9775) >>> _zz_935);
  assign _zz_9775 = _zz_9776;
  assign _zz_9776 = ($signed(_zz_9778) + $signed(_zz_932));
  assign _zz_9777 = ({9'd0,data_mid_5_26_imag} <<< 9);
  assign _zz_9778 = {{9{_zz_9777[26]}}, _zz_9777};
  assign _zz_9779 = fixTo_1121_dout;
  assign _zz_9780 = ($signed(twiddle_factor_table_58_real) + $signed(twiddle_factor_table_58_imag));
  assign _zz_9781 = ($signed(_zz_938) - $signed(_zz_9782));
  assign _zz_9782 = ($signed(_zz_9783) * $signed(twiddle_factor_table_58_imag));
  assign _zz_9783 = ($signed(data_mid_5_59_real) + $signed(data_mid_5_59_imag));
  assign _zz_9784 = fixTo_1122_dout;
  assign _zz_9785 = ($signed(_zz_938) + $signed(_zz_9786));
  assign _zz_9786 = ($signed(_zz_9787) * $signed(twiddle_factor_table_58_real));
  assign _zz_9787 = ($signed(data_mid_5_59_imag) - $signed(data_mid_5_59_real));
  assign _zz_9788 = fixTo_1123_dout;
  assign _zz_9789 = _zz_9790[35 : 0];
  assign _zz_9790 = _zz_9791;
  assign _zz_9791 = ($signed(_zz_9792) >>> _zz_939);
  assign _zz_9792 = _zz_9793;
  assign _zz_9793 = ($signed(_zz_9795) - $signed(_zz_936));
  assign _zz_9794 = ({9'd0,data_mid_5_27_real} <<< 9);
  assign _zz_9795 = {{9{_zz_9794[26]}}, _zz_9794};
  assign _zz_9796 = fixTo_1124_dout;
  assign _zz_9797 = _zz_9798[35 : 0];
  assign _zz_9798 = _zz_9799;
  assign _zz_9799 = ($signed(_zz_9800) >>> _zz_939);
  assign _zz_9800 = _zz_9801;
  assign _zz_9801 = ($signed(_zz_9803) - $signed(_zz_937));
  assign _zz_9802 = ({9'd0,data_mid_5_27_imag} <<< 9);
  assign _zz_9803 = {{9{_zz_9802[26]}}, _zz_9802};
  assign _zz_9804 = fixTo_1125_dout;
  assign _zz_9805 = _zz_9806[35 : 0];
  assign _zz_9806 = _zz_9807;
  assign _zz_9807 = ($signed(_zz_9808) >>> _zz_940);
  assign _zz_9808 = _zz_9809;
  assign _zz_9809 = ($signed(_zz_9811) + $signed(_zz_936));
  assign _zz_9810 = ({9'd0,data_mid_5_27_real} <<< 9);
  assign _zz_9811 = {{9{_zz_9810[26]}}, _zz_9810};
  assign _zz_9812 = fixTo_1126_dout;
  assign _zz_9813 = _zz_9814[35 : 0];
  assign _zz_9814 = _zz_9815;
  assign _zz_9815 = ($signed(_zz_9816) >>> _zz_940);
  assign _zz_9816 = _zz_9817;
  assign _zz_9817 = ($signed(_zz_9819) + $signed(_zz_937));
  assign _zz_9818 = ({9'd0,data_mid_5_27_imag} <<< 9);
  assign _zz_9819 = {{9{_zz_9818[26]}}, _zz_9818};
  assign _zz_9820 = fixTo_1127_dout;
  assign _zz_9821 = ($signed(twiddle_factor_table_59_real) + $signed(twiddle_factor_table_59_imag));
  assign _zz_9822 = ($signed(_zz_943) - $signed(_zz_9823));
  assign _zz_9823 = ($signed(_zz_9824) * $signed(twiddle_factor_table_59_imag));
  assign _zz_9824 = ($signed(data_mid_5_60_real) + $signed(data_mid_5_60_imag));
  assign _zz_9825 = fixTo_1128_dout;
  assign _zz_9826 = ($signed(_zz_943) + $signed(_zz_9827));
  assign _zz_9827 = ($signed(_zz_9828) * $signed(twiddle_factor_table_59_real));
  assign _zz_9828 = ($signed(data_mid_5_60_imag) - $signed(data_mid_5_60_real));
  assign _zz_9829 = fixTo_1129_dout;
  assign _zz_9830 = _zz_9831[35 : 0];
  assign _zz_9831 = _zz_9832;
  assign _zz_9832 = ($signed(_zz_9833) >>> _zz_944);
  assign _zz_9833 = _zz_9834;
  assign _zz_9834 = ($signed(_zz_9836) - $signed(_zz_941));
  assign _zz_9835 = ({9'd0,data_mid_5_28_real} <<< 9);
  assign _zz_9836 = {{9{_zz_9835[26]}}, _zz_9835};
  assign _zz_9837 = fixTo_1130_dout;
  assign _zz_9838 = _zz_9839[35 : 0];
  assign _zz_9839 = _zz_9840;
  assign _zz_9840 = ($signed(_zz_9841) >>> _zz_944);
  assign _zz_9841 = _zz_9842;
  assign _zz_9842 = ($signed(_zz_9844) - $signed(_zz_942));
  assign _zz_9843 = ({9'd0,data_mid_5_28_imag} <<< 9);
  assign _zz_9844 = {{9{_zz_9843[26]}}, _zz_9843};
  assign _zz_9845 = fixTo_1131_dout;
  assign _zz_9846 = _zz_9847[35 : 0];
  assign _zz_9847 = _zz_9848;
  assign _zz_9848 = ($signed(_zz_9849) >>> _zz_945);
  assign _zz_9849 = _zz_9850;
  assign _zz_9850 = ($signed(_zz_9852) + $signed(_zz_941));
  assign _zz_9851 = ({9'd0,data_mid_5_28_real} <<< 9);
  assign _zz_9852 = {{9{_zz_9851[26]}}, _zz_9851};
  assign _zz_9853 = fixTo_1132_dout;
  assign _zz_9854 = _zz_9855[35 : 0];
  assign _zz_9855 = _zz_9856;
  assign _zz_9856 = ($signed(_zz_9857) >>> _zz_945);
  assign _zz_9857 = _zz_9858;
  assign _zz_9858 = ($signed(_zz_9860) + $signed(_zz_942));
  assign _zz_9859 = ({9'd0,data_mid_5_28_imag} <<< 9);
  assign _zz_9860 = {{9{_zz_9859[26]}}, _zz_9859};
  assign _zz_9861 = fixTo_1133_dout;
  assign _zz_9862 = ($signed(twiddle_factor_table_60_real) + $signed(twiddle_factor_table_60_imag));
  assign _zz_9863 = ($signed(_zz_948) - $signed(_zz_9864));
  assign _zz_9864 = ($signed(_zz_9865) * $signed(twiddle_factor_table_60_imag));
  assign _zz_9865 = ($signed(data_mid_5_61_real) + $signed(data_mid_5_61_imag));
  assign _zz_9866 = fixTo_1134_dout;
  assign _zz_9867 = ($signed(_zz_948) + $signed(_zz_9868));
  assign _zz_9868 = ($signed(_zz_9869) * $signed(twiddle_factor_table_60_real));
  assign _zz_9869 = ($signed(data_mid_5_61_imag) - $signed(data_mid_5_61_real));
  assign _zz_9870 = fixTo_1135_dout;
  assign _zz_9871 = _zz_9872[35 : 0];
  assign _zz_9872 = _zz_9873;
  assign _zz_9873 = ($signed(_zz_9874) >>> _zz_949);
  assign _zz_9874 = _zz_9875;
  assign _zz_9875 = ($signed(_zz_9877) - $signed(_zz_946));
  assign _zz_9876 = ({9'd0,data_mid_5_29_real} <<< 9);
  assign _zz_9877 = {{9{_zz_9876[26]}}, _zz_9876};
  assign _zz_9878 = fixTo_1136_dout;
  assign _zz_9879 = _zz_9880[35 : 0];
  assign _zz_9880 = _zz_9881;
  assign _zz_9881 = ($signed(_zz_9882) >>> _zz_949);
  assign _zz_9882 = _zz_9883;
  assign _zz_9883 = ($signed(_zz_9885) - $signed(_zz_947));
  assign _zz_9884 = ({9'd0,data_mid_5_29_imag} <<< 9);
  assign _zz_9885 = {{9{_zz_9884[26]}}, _zz_9884};
  assign _zz_9886 = fixTo_1137_dout;
  assign _zz_9887 = _zz_9888[35 : 0];
  assign _zz_9888 = _zz_9889;
  assign _zz_9889 = ($signed(_zz_9890) >>> _zz_950);
  assign _zz_9890 = _zz_9891;
  assign _zz_9891 = ($signed(_zz_9893) + $signed(_zz_946));
  assign _zz_9892 = ({9'd0,data_mid_5_29_real} <<< 9);
  assign _zz_9893 = {{9{_zz_9892[26]}}, _zz_9892};
  assign _zz_9894 = fixTo_1138_dout;
  assign _zz_9895 = _zz_9896[35 : 0];
  assign _zz_9896 = _zz_9897;
  assign _zz_9897 = ($signed(_zz_9898) >>> _zz_950);
  assign _zz_9898 = _zz_9899;
  assign _zz_9899 = ($signed(_zz_9901) + $signed(_zz_947));
  assign _zz_9900 = ({9'd0,data_mid_5_29_imag} <<< 9);
  assign _zz_9901 = {{9{_zz_9900[26]}}, _zz_9900};
  assign _zz_9902 = fixTo_1139_dout;
  assign _zz_9903 = ($signed(twiddle_factor_table_61_real) + $signed(twiddle_factor_table_61_imag));
  assign _zz_9904 = ($signed(_zz_953) - $signed(_zz_9905));
  assign _zz_9905 = ($signed(_zz_9906) * $signed(twiddle_factor_table_61_imag));
  assign _zz_9906 = ($signed(data_mid_5_62_real) + $signed(data_mid_5_62_imag));
  assign _zz_9907 = fixTo_1140_dout;
  assign _zz_9908 = ($signed(_zz_953) + $signed(_zz_9909));
  assign _zz_9909 = ($signed(_zz_9910) * $signed(twiddle_factor_table_61_real));
  assign _zz_9910 = ($signed(data_mid_5_62_imag) - $signed(data_mid_5_62_real));
  assign _zz_9911 = fixTo_1141_dout;
  assign _zz_9912 = _zz_9913[35 : 0];
  assign _zz_9913 = _zz_9914;
  assign _zz_9914 = ($signed(_zz_9915) >>> _zz_954);
  assign _zz_9915 = _zz_9916;
  assign _zz_9916 = ($signed(_zz_9918) - $signed(_zz_951));
  assign _zz_9917 = ({9'd0,data_mid_5_30_real} <<< 9);
  assign _zz_9918 = {{9{_zz_9917[26]}}, _zz_9917};
  assign _zz_9919 = fixTo_1142_dout;
  assign _zz_9920 = _zz_9921[35 : 0];
  assign _zz_9921 = _zz_9922;
  assign _zz_9922 = ($signed(_zz_9923) >>> _zz_954);
  assign _zz_9923 = _zz_9924;
  assign _zz_9924 = ($signed(_zz_9926) - $signed(_zz_952));
  assign _zz_9925 = ({9'd0,data_mid_5_30_imag} <<< 9);
  assign _zz_9926 = {{9{_zz_9925[26]}}, _zz_9925};
  assign _zz_9927 = fixTo_1143_dout;
  assign _zz_9928 = _zz_9929[35 : 0];
  assign _zz_9929 = _zz_9930;
  assign _zz_9930 = ($signed(_zz_9931) >>> _zz_955);
  assign _zz_9931 = _zz_9932;
  assign _zz_9932 = ($signed(_zz_9934) + $signed(_zz_951));
  assign _zz_9933 = ({9'd0,data_mid_5_30_real} <<< 9);
  assign _zz_9934 = {{9{_zz_9933[26]}}, _zz_9933};
  assign _zz_9935 = fixTo_1144_dout;
  assign _zz_9936 = _zz_9937[35 : 0];
  assign _zz_9937 = _zz_9938;
  assign _zz_9938 = ($signed(_zz_9939) >>> _zz_955);
  assign _zz_9939 = _zz_9940;
  assign _zz_9940 = ($signed(_zz_9942) + $signed(_zz_952));
  assign _zz_9941 = ({9'd0,data_mid_5_30_imag} <<< 9);
  assign _zz_9942 = {{9{_zz_9941[26]}}, _zz_9941};
  assign _zz_9943 = fixTo_1145_dout;
  assign _zz_9944 = ($signed(twiddle_factor_table_62_real) + $signed(twiddle_factor_table_62_imag));
  assign _zz_9945 = ($signed(_zz_958) - $signed(_zz_9946));
  assign _zz_9946 = ($signed(_zz_9947) * $signed(twiddle_factor_table_62_imag));
  assign _zz_9947 = ($signed(data_mid_5_63_real) + $signed(data_mid_5_63_imag));
  assign _zz_9948 = fixTo_1146_dout;
  assign _zz_9949 = ($signed(_zz_958) + $signed(_zz_9950));
  assign _zz_9950 = ($signed(_zz_9951) * $signed(twiddle_factor_table_62_real));
  assign _zz_9951 = ($signed(data_mid_5_63_imag) - $signed(data_mid_5_63_real));
  assign _zz_9952 = fixTo_1147_dout;
  assign _zz_9953 = _zz_9954[35 : 0];
  assign _zz_9954 = _zz_9955;
  assign _zz_9955 = ($signed(_zz_9956) >>> _zz_959);
  assign _zz_9956 = _zz_9957;
  assign _zz_9957 = ($signed(_zz_9959) - $signed(_zz_956));
  assign _zz_9958 = ({9'd0,data_mid_5_31_real} <<< 9);
  assign _zz_9959 = {{9{_zz_9958[26]}}, _zz_9958};
  assign _zz_9960 = fixTo_1148_dout;
  assign _zz_9961 = _zz_9962[35 : 0];
  assign _zz_9962 = _zz_9963;
  assign _zz_9963 = ($signed(_zz_9964) >>> _zz_959);
  assign _zz_9964 = _zz_9965;
  assign _zz_9965 = ($signed(_zz_9967) - $signed(_zz_957));
  assign _zz_9966 = ({9'd0,data_mid_5_31_imag} <<< 9);
  assign _zz_9967 = {{9{_zz_9966[26]}}, _zz_9966};
  assign _zz_9968 = fixTo_1149_dout;
  assign _zz_9969 = _zz_9970[35 : 0];
  assign _zz_9970 = _zz_9971;
  assign _zz_9971 = ($signed(_zz_9972) >>> _zz_960);
  assign _zz_9972 = _zz_9973;
  assign _zz_9973 = ($signed(_zz_9975) + $signed(_zz_956));
  assign _zz_9974 = ({9'd0,data_mid_5_31_real} <<< 9);
  assign _zz_9975 = {{9{_zz_9974[26]}}, _zz_9974};
  assign _zz_9976 = fixTo_1150_dout;
  assign _zz_9977 = _zz_9978[35 : 0];
  assign _zz_9978 = _zz_9979;
  assign _zz_9979 = ($signed(_zz_9980) >>> _zz_960);
  assign _zz_9980 = _zz_9981;
  assign _zz_9981 = ($signed(_zz_9983) + $signed(_zz_957));
  assign _zz_9982 = ({9'd0,data_mid_5_31_imag} <<< 9);
  assign _zz_9983 = {{9{_zz_9982[26]}}, _zz_9982};
  assign _zz_9984 = fixTo_1151_dout;
  SInt36fixTo35_0_ROUNDTOINF fixTo (
    .din     (_zz_961[35:0]     ), //i
    .dout    (fixTo_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1 (
    .din     (_zz_962[35:0]       ), //i
    .dout    (fixTo_1_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_2 (
    .din     (_zz_963[35:0]       ), //i
    .dout    (fixTo_2_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_3 (
    .din     (_zz_964[35:0]       ), //i
    .dout    (fixTo_3_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_4 (
    .din     (_zz_965[35:0]       ), //i
    .dout    (fixTo_4_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_5 (
    .din     (_zz_966[35:0]       ), //i
    .dout    (fixTo_5_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_6 (
    .din     (_zz_967[35:0]       ), //i
    .dout    (fixTo_6_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_7 (
    .din     (_zz_968[35:0]       ), //i
    .dout    (fixTo_7_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_8 (
    .din     (_zz_969[35:0]       ), //i
    .dout    (fixTo_8_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_9 (
    .din     (_zz_970[35:0]       ), //i
    .dout    (fixTo_9_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_10 (
    .din     (_zz_971[35:0]        ), //i
    .dout    (fixTo_10_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_11 (
    .din     (_zz_972[35:0]        ), //i
    .dout    (fixTo_11_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_12 (
    .din     (_zz_973[35:0]        ), //i
    .dout    (fixTo_12_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_13 (
    .din     (_zz_974[35:0]        ), //i
    .dout    (fixTo_13_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_14 (
    .din     (_zz_975[35:0]        ), //i
    .dout    (fixTo_14_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_15 (
    .din     (_zz_976[35:0]        ), //i
    .dout    (fixTo_15_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_16 (
    .din     (_zz_977[35:0]        ), //i
    .dout    (fixTo_16_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_17 (
    .din     (_zz_978[35:0]        ), //i
    .dout    (fixTo_17_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_18 (
    .din     (_zz_979[35:0]        ), //i
    .dout    (fixTo_18_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_19 (
    .din     (_zz_980[35:0]        ), //i
    .dout    (fixTo_19_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_20 (
    .din     (_zz_981[35:0]        ), //i
    .dout    (fixTo_20_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_21 (
    .din     (_zz_982[35:0]        ), //i
    .dout    (fixTo_21_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_22 (
    .din     (_zz_983[35:0]        ), //i
    .dout    (fixTo_22_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_23 (
    .din     (_zz_984[35:0]        ), //i
    .dout    (fixTo_23_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_24 (
    .din     (_zz_985[35:0]        ), //i
    .dout    (fixTo_24_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_25 (
    .din     (_zz_986[35:0]        ), //i
    .dout    (fixTo_25_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_26 (
    .din     (_zz_987[35:0]        ), //i
    .dout    (fixTo_26_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_27 (
    .din     (_zz_988[35:0]        ), //i
    .dout    (fixTo_27_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_28 (
    .din     (_zz_989[35:0]        ), //i
    .dout    (fixTo_28_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_29 (
    .din     (_zz_990[35:0]        ), //i
    .dout    (fixTo_29_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_30 (
    .din     (_zz_991[35:0]        ), //i
    .dout    (fixTo_30_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_31 (
    .din     (_zz_992[35:0]        ), //i
    .dout    (fixTo_31_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_32 (
    .din     (_zz_993[35:0]        ), //i
    .dout    (fixTo_32_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_33 (
    .din     (_zz_994[35:0]        ), //i
    .dout    (fixTo_33_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_34 (
    .din     (_zz_995[35:0]        ), //i
    .dout    (fixTo_34_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_35 (
    .din     (_zz_996[35:0]        ), //i
    .dout    (fixTo_35_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_36 (
    .din     (_zz_997[35:0]        ), //i
    .dout    (fixTo_36_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_37 (
    .din     (_zz_998[35:0]        ), //i
    .dout    (fixTo_37_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_38 (
    .din     (_zz_999[35:0]        ), //i
    .dout    (fixTo_38_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_39 (
    .din     (_zz_1000[35:0]       ), //i
    .dout    (fixTo_39_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_40 (
    .din     (_zz_1001[35:0]       ), //i
    .dout    (fixTo_40_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_41 (
    .din     (_zz_1002[35:0]       ), //i
    .dout    (fixTo_41_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_42 (
    .din     (_zz_1003[35:0]       ), //i
    .dout    (fixTo_42_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_43 (
    .din     (_zz_1004[35:0]       ), //i
    .dout    (fixTo_43_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_44 (
    .din     (_zz_1005[35:0]       ), //i
    .dout    (fixTo_44_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_45 (
    .din     (_zz_1006[35:0]       ), //i
    .dout    (fixTo_45_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_46 (
    .din     (_zz_1007[35:0]       ), //i
    .dout    (fixTo_46_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_47 (
    .din     (_zz_1008[35:0]       ), //i
    .dout    (fixTo_47_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_48 (
    .din     (_zz_1009[35:0]       ), //i
    .dout    (fixTo_48_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_49 (
    .din     (_zz_1010[35:0]       ), //i
    .dout    (fixTo_49_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_50 (
    .din     (_zz_1011[35:0]       ), //i
    .dout    (fixTo_50_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_51 (
    .din     (_zz_1012[35:0]       ), //i
    .dout    (fixTo_51_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_52 (
    .din     (_zz_1013[35:0]       ), //i
    .dout    (fixTo_52_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_53 (
    .din     (_zz_1014[35:0]       ), //i
    .dout    (fixTo_53_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_54 (
    .din     (_zz_1015[35:0]       ), //i
    .dout    (fixTo_54_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_55 (
    .din     (_zz_1016[35:0]       ), //i
    .dout    (fixTo_55_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_56 (
    .din     (_zz_1017[35:0]       ), //i
    .dout    (fixTo_56_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_57 (
    .din     (_zz_1018[35:0]       ), //i
    .dout    (fixTo_57_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_58 (
    .din     (_zz_1019[35:0]       ), //i
    .dout    (fixTo_58_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_59 (
    .din     (_zz_1020[35:0]       ), //i
    .dout    (fixTo_59_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_60 (
    .din     (_zz_1021[35:0]       ), //i
    .dout    (fixTo_60_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_61 (
    .din     (_zz_1022[35:0]       ), //i
    .dout    (fixTo_61_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_62 (
    .din     (_zz_1023[35:0]       ), //i
    .dout    (fixTo_62_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_63 (
    .din     (_zz_1024[35:0]       ), //i
    .dout    (fixTo_63_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_64 (
    .din     (_zz_1025[35:0]       ), //i
    .dout    (fixTo_64_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_65 (
    .din     (_zz_1026[35:0]       ), //i
    .dout    (fixTo_65_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_66 (
    .din     (_zz_1027[35:0]       ), //i
    .dout    (fixTo_66_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_67 (
    .din     (_zz_1028[35:0]       ), //i
    .dout    (fixTo_67_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_68 (
    .din     (_zz_1029[35:0]       ), //i
    .dout    (fixTo_68_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_69 (
    .din     (_zz_1030[35:0]       ), //i
    .dout    (fixTo_69_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_70 (
    .din     (_zz_1031[35:0]       ), //i
    .dout    (fixTo_70_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_71 (
    .din     (_zz_1032[35:0]       ), //i
    .dout    (fixTo_71_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_72 (
    .din     (_zz_1033[35:0]       ), //i
    .dout    (fixTo_72_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_73 (
    .din     (_zz_1034[35:0]       ), //i
    .dout    (fixTo_73_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_74 (
    .din     (_zz_1035[35:0]       ), //i
    .dout    (fixTo_74_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_75 (
    .din     (_zz_1036[35:0]       ), //i
    .dout    (fixTo_75_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_76 (
    .din     (_zz_1037[35:0]       ), //i
    .dout    (fixTo_76_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_77 (
    .din     (_zz_1038[35:0]       ), //i
    .dout    (fixTo_77_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_78 (
    .din     (_zz_1039[35:0]       ), //i
    .dout    (fixTo_78_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_79 (
    .din     (_zz_1040[35:0]       ), //i
    .dout    (fixTo_79_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_80 (
    .din     (_zz_1041[35:0]       ), //i
    .dout    (fixTo_80_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_81 (
    .din     (_zz_1042[35:0]       ), //i
    .dout    (fixTo_81_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_82 (
    .din     (_zz_1043[35:0]       ), //i
    .dout    (fixTo_82_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_83 (
    .din     (_zz_1044[35:0]       ), //i
    .dout    (fixTo_83_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_84 (
    .din     (_zz_1045[35:0]       ), //i
    .dout    (fixTo_84_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_85 (
    .din     (_zz_1046[35:0]       ), //i
    .dout    (fixTo_85_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_86 (
    .din     (_zz_1047[35:0]       ), //i
    .dout    (fixTo_86_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_87 (
    .din     (_zz_1048[35:0]       ), //i
    .dout    (fixTo_87_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_88 (
    .din     (_zz_1049[35:0]       ), //i
    .dout    (fixTo_88_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_89 (
    .din     (_zz_1050[35:0]       ), //i
    .dout    (fixTo_89_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_90 (
    .din     (_zz_1051[35:0]       ), //i
    .dout    (fixTo_90_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_91 (
    .din     (_zz_1052[35:0]       ), //i
    .dout    (fixTo_91_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_92 (
    .din     (_zz_1053[35:0]       ), //i
    .dout    (fixTo_92_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_93 (
    .din     (_zz_1054[35:0]       ), //i
    .dout    (fixTo_93_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_94 (
    .din     (_zz_1055[35:0]       ), //i
    .dout    (fixTo_94_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_95 (
    .din     (_zz_1056[35:0]       ), //i
    .dout    (fixTo_95_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_96 (
    .din     (_zz_1057[35:0]       ), //i
    .dout    (fixTo_96_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_97 (
    .din     (_zz_1058[35:0]       ), //i
    .dout    (fixTo_97_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_98 (
    .din     (_zz_1059[35:0]       ), //i
    .dout    (fixTo_98_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_99 (
    .din     (_zz_1060[35:0]       ), //i
    .dout    (fixTo_99_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_100 (
    .din     (_zz_1061[35:0]        ), //i
    .dout    (fixTo_100_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_101 (
    .din     (_zz_1062[35:0]        ), //i
    .dout    (fixTo_101_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_102 (
    .din     (_zz_1063[35:0]        ), //i
    .dout    (fixTo_102_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_103 (
    .din     (_zz_1064[35:0]        ), //i
    .dout    (fixTo_103_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_104 (
    .din     (_zz_1065[35:0]        ), //i
    .dout    (fixTo_104_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_105 (
    .din     (_zz_1066[35:0]        ), //i
    .dout    (fixTo_105_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_106 (
    .din     (_zz_1067[35:0]        ), //i
    .dout    (fixTo_106_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_107 (
    .din     (_zz_1068[35:0]        ), //i
    .dout    (fixTo_107_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_108 (
    .din     (_zz_1069[35:0]        ), //i
    .dout    (fixTo_108_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_109 (
    .din     (_zz_1070[35:0]        ), //i
    .dout    (fixTo_109_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_110 (
    .din     (_zz_1071[35:0]        ), //i
    .dout    (fixTo_110_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_111 (
    .din     (_zz_1072[35:0]        ), //i
    .dout    (fixTo_111_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_112 (
    .din     (_zz_1073[35:0]        ), //i
    .dout    (fixTo_112_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_113 (
    .din     (_zz_1074[35:0]        ), //i
    .dout    (fixTo_113_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_114 (
    .din     (_zz_1075[35:0]        ), //i
    .dout    (fixTo_114_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_115 (
    .din     (_zz_1076[35:0]        ), //i
    .dout    (fixTo_115_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_116 (
    .din     (_zz_1077[35:0]        ), //i
    .dout    (fixTo_116_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_117 (
    .din     (_zz_1078[35:0]        ), //i
    .dout    (fixTo_117_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_118 (
    .din     (_zz_1079[35:0]        ), //i
    .dout    (fixTo_118_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_119 (
    .din     (_zz_1080[35:0]        ), //i
    .dout    (fixTo_119_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_120 (
    .din     (_zz_1081[35:0]        ), //i
    .dout    (fixTo_120_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_121 (
    .din     (_zz_1082[35:0]        ), //i
    .dout    (fixTo_121_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_122 (
    .din     (_zz_1083[35:0]        ), //i
    .dout    (fixTo_122_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_123 (
    .din     (_zz_1084[35:0]        ), //i
    .dout    (fixTo_123_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_124 (
    .din     (_zz_1085[35:0]        ), //i
    .dout    (fixTo_124_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_125 (
    .din     (_zz_1086[35:0]        ), //i
    .dout    (fixTo_125_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_126 (
    .din     (_zz_1087[35:0]        ), //i
    .dout    (fixTo_126_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_127 (
    .din     (_zz_1088[35:0]        ), //i
    .dout    (fixTo_127_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_128 (
    .din     (_zz_1089[35:0]        ), //i
    .dout    (fixTo_128_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_129 (
    .din     (_zz_1090[35:0]        ), //i
    .dout    (fixTo_129_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_130 (
    .din     (_zz_1091[35:0]        ), //i
    .dout    (fixTo_130_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_131 (
    .din     (_zz_1092[35:0]        ), //i
    .dout    (fixTo_131_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_132 (
    .din     (_zz_1093[35:0]        ), //i
    .dout    (fixTo_132_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_133 (
    .din     (_zz_1094[35:0]        ), //i
    .dout    (fixTo_133_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_134 (
    .din     (_zz_1095[35:0]        ), //i
    .dout    (fixTo_134_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_135 (
    .din     (_zz_1096[35:0]        ), //i
    .dout    (fixTo_135_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_136 (
    .din     (_zz_1097[35:0]        ), //i
    .dout    (fixTo_136_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_137 (
    .din     (_zz_1098[35:0]        ), //i
    .dout    (fixTo_137_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_138 (
    .din     (_zz_1099[35:0]        ), //i
    .dout    (fixTo_138_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_139 (
    .din     (_zz_1100[35:0]        ), //i
    .dout    (fixTo_139_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_140 (
    .din     (_zz_1101[35:0]        ), //i
    .dout    (fixTo_140_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_141 (
    .din     (_zz_1102[35:0]        ), //i
    .dout    (fixTo_141_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_142 (
    .din     (_zz_1103[35:0]        ), //i
    .dout    (fixTo_142_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_143 (
    .din     (_zz_1104[35:0]        ), //i
    .dout    (fixTo_143_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_144 (
    .din     (_zz_1105[35:0]        ), //i
    .dout    (fixTo_144_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_145 (
    .din     (_zz_1106[35:0]        ), //i
    .dout    (fixTo_145_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_146 (
    .din     (_zz_1107[35:0]        ), //i
    .dout    (fixTo_146_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_147 (
    .din     (_zz_1108[35:0]        ), //i
    .dout    (fixTo_147_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_148 (
    .din     (_zz_1109[35:0]        ), //i
    .dout    (fixTo_148_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_149 (
    .din     (_zz_1110[35:0]        ), //i
    .dout    (fixTo_149_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_150 (
    .din     (_zz_1111[35:0]        ), //i
    .dout    (fixTo_150_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_151 (
    .din     (_zz_1112[35:0]        ), //i
    .dout    (fixTo_151_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_152 (
    .din     (_zz_1113[35:0]        ), //i
    .dout    (fixTo_152_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_153 (
    .din     (_zz_1114[35:0]        ), //i
    .dout    (fixTo_153_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_154 (
    .din     (_zz_1115[35:0]        ), //i
    .dout    (fixTo_154_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_155 (
    .din     (_zz_1116[35:0]        ), //i
    .dout    (fixTo_155_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_156 (
    .din     (_zz_1117[35:0]        ), //i
    .dout    (fixTo_156_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_157 (
    .din     (_zz_1118[35:0]        ), //i
    .dout    (fixTo_157_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_158 (
    .din     (_zz_1119[35:0]        ), //i
    .dout    (fixTo_158_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_159 (
    .din     (_zz_1120[35:0]        ), //i
    .dout    (fixTo_159_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_160 (
    .din     (_zz_1121[35:0]        ), //i
    .dout    (fixTo_160_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_161 (
    .din     (_zz_1122[35:0]        ), //i
    .dout    (fixTo_161_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_162 (
    .din     (_zz_1123[35:0]        ), //i
    .dout    (fixTo_162_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_163 (
    .din     (_zz_1124[35:0]        ), //i
    .dout    (fixTo_163_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_164 (
    .din     (_zz_1125[35:0]        ), //i
    .dout    (fixTo_164_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_165 (
    .din     (_zz_1126[35:0]        ), //i
    .dout    (fixTo_165_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_166 (
    .din     (_zz_1127[35:0]        ), //i
    .dout    (fixTo_166_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_167 (
    .din     (_zz_1128[35:0]        ), //i
    .dout    (fixTo_167_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_168 (
    .din     (_zz_1129[35:0]        ), //i
    .dout    (fixTo_168_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_169 (
    .din     (_zz_1130[35:0]        ), //i
    .dout    (fixTo_169_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_170 (
    .din     (_zz_1131[35:0]        ), //i
    .dout    (fixTo_170_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_171 (
    .din     (_zz_1132[35:0]        ), //i
    .dout    (fixTo_171_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_172 (
    .din     (_zz_1133[35:0]        ), //i
    .dout    (fixTo_172_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_173 (
    .din     (_zz_1134[35:0]        ), //i
    .dout    (fixTo_173_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_174 (
    .din     (_zz_1135[35:0]        ), //i
    .dout    (fixTo_174_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_175 (
    .din     (_zz_1136[35:0]        ), //i
    .dout    (fixTo_175_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_176 (
    .din     (_zz_1137[35:0]        ), //i
    .dout    (fixTo_176_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_177 (
    .din     (_zz_1138[35:0]        ), //i
    .dout    (fixTo_177_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_178 (
    .din     (_zz_1139[35:0]        ), //i
    .dout    (fixTo_178_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_179 (
    .din     (_zz_1140[35:0]        ), //i
    .dout    (fixTo_179_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_180 (
    .din     (_zz_1141[35:0]        ), //i
    .dout    (fixTo_180_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_181 (
    .din     (_zz_1142[35:0]        ), //i
    .dout    (fixTo_181_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_182 (
    .din     (_zz_1143[35:0]        ), //i
    .dout    (fixTo_182_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_183 (
    .din     (_zz_1144[35:0]        ), //i
    .dout    (fixTo_183_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_184 (
    .din     (_zz_1145[35:0]        ), //i
    .dout    (fixTo_184_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_185 (
    .din     (_zz_1146[35:0]        ), //i
    .dout    (fixTo_185_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_186 (
    .din     (_zz_1147[35:0]        ), //i
    .dout    (fixTo_186_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_187 (
    .din     (_zz_1148[35:0]        ), //i
    .dout    (fixTo_187_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_188 (
    .din     (_zz_1149[35:0]        ), //i
    .dout    (fixTo_188_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_189 (
    .din     (_zz_1150[35:0]        ), //i
    .dout    (fixTo_189_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_190 (
    .din     (_zz_1151[35:0]        ), //i
    .dout    (fixTo_190_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_191 (
    .din     (_zz_1152[35:0]        ), //i
    .dout    (fixTo_191_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_192 (
    .din     (_zz_1153[35:0]        ), //i
    .dout    (fixTo_192_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_193 (
    .din     (_zz_1154[35:0]        ), //i
    .dout    (fixTo_193_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_194 (
    .din     (_zz_1155[35:0]        ), //i
    .dout    (fixTo_194_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_195 (
    .din     (_zz_1156[35:0]        ), //i
    .dout    (fixTo_195_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_196 (
    .din     (_zz_1157[35:0]        ), //i
    .dout    (fixTo_196_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_197 (
    .din     (_zz_1158[35:0]        ), //i
    .dout    (fixTo_197_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_198 (
    .din     (_zz_1159[35:0]        ), //i
    .dout    (fixTo_198_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_199 (
    .din     (_zz_1160[35:0]        ), //i
    .dout    (fixTo_199_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_200 (
    .din     (_zz_1161[35:0]        ), //i
    .dout    (fixTo_200_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_201 (
    .din     (_zz_1162[35:0]        ), //i
    .dout    (fixTo_201_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_202 (
    .din     (_zz_1163[35:0]        ), //i
    .dout    (fixTo_202_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_203 (
    .din     (_zz_1164[35:0]        ), //i
    .dout    (fixTo_203_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_204 (
    .din     (_zz_1165[35:0]        ), //i
    .dout    (fixTo_204_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_205 (
    .din     (_zz_1166[35:0]        ), //i
    .dout    (fixTo_205_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_206 (
    .din     (_zz_1167[35:0]        ), //i
    .dout    (fixTo_206_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_207 (
    .din     (_zz_1168[35:0]        ), //i
    .dout    (fixTo_207_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_208 (
    .din     (_zz_1169[35:0]        ), //i
    .dout    (fixTo_208_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_209 (
    .din     (_zz_1170[35:0]        ), //i
    .dout    (fixTo_209_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_210 (
    .din     (_zz_1171[35:0]        ), //i
    .dout    (fixTo_210_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_211 (
    .din     (_zz_1172[35:0]        ), //i
    .dout    (fixTo_211_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_212 (
    .din     (_zz_1173[35:0]        ), //i
    .dout    (fixTo_212_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_213 (
    .din     (_zz_1174[35:0]        ), //i
    .dout    (fixTo_213_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_214 (
    .din     (_zz_1175[35:0]        ), //i
    .dout    (fixTo_214_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_215 (
    .din     (_zz_1176[35:0]        ), //i
    .dout    (fixTo_215_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_216 (
    .din     (_zz_1177[35:0]        ), //i
    .dout    (fixTo_216_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_217 (
    .din     (_zz_1178[35:0]        ), //i
    .dout    (fixTo_217_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_218 (
    .din     (_zz_1179[35:0]        ), //i
    .dout    (fixTo_218_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_219 (
    .din     (_zz_1180[35:0]        ), //i
    .dout    (fixTo_219_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_220 (
    .din     (_zz_1181[35:0]        ), //i
    .dout    (fixTo_220_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_221 (
    .din     (_zz_1182[35:0]        ), //i
    .dout    (fixTo_221_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_222 (
    .din     (_zz_1183[35:0]        ), //i
    .dout    (fixTo_222_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_223 (
    .din     (_zz_1184[35:0]        ), //i
    .dout    (fixTo_223_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_224 (
    .din     (_zz_1185[35:0]        ), //i
    .dout    (fixTo_224_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_225 (
    .din     (_zz_1186[35:0]        ), //i
    .dout    (fixTo_225_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_226 (
    .din     (_zz_1187[35:0]        ), //i
    .dout    (fixTo_226_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_227 (
    .din     (_zz_1188[35:0]        ), //i
    .dout    (fixTo_227_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_228 (
    .din     (_zz_1189[35:0]        ), //i
    .dout    (fixTo_228_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_229 (
    .din     (_zz_1190[35:0]        ), //i
    .dout    (fixTo_229_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_230 (
    .din     (_zz_1191[35:0]        ), //i
    .dout    (fixTo_230_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_231 (
    .din     (_zz_1192[35:0]        ), //i
    .dout    (fixTo_231_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_232 (
    .din     (_zz_1193[35:0]        ), //i
    .dout    (fixTo_232_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_233 (
    .din     (_zz_1194[35:0]        ), //i
    .dout    (fixTo_233_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_234 (
    .din     (_zz_1195[35:0]        ), //i
    .dout    (fixTo_234_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_235 (
    .din     (_zz_1196[35:0]        ), //i
    .dout    (fixTo_235_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_236 (
    .din     (_zz_1197[35:0]        ), //i
    .dout    (fixTo_236_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_237 (
    .din     (_zz_1198[35:0]        ), //i
    .dout    (fixTo_237_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_238 (
    .din     (_zz_1199[35:0]        ), //i
    .dout    (fixTo_238_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_239 (
    .din     (_zz_1200[35:0]        ), //i
    .dout    (fixTo_239_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_240 (
    .din     (_zz_1201[35:0]        ), //i
    .dout    (fixTo_240_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_241 (
    .din     (_zz_1202[35:0]        ), //i
    .dout    (fixTo_241_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_242 (
    .din     (_zz_1203[35:0]        ), //i
    .dout    (fixTo_242_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_243 (
    .din     (_zz_1204[35:0]        ), //i
    .dout    (fixTo_243_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_244 (
    .din     (_zz_1205[35:0]        ), //i
    .dout    (fixTo_244_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_245 (
    .din     (_zz_1206[35:0]        ), //i
    .dout    (fixTo_245_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_246 (
    .din     (_zz_1207[35:0]        ), //i
    .dout    (fixTo_246_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_247 (
    .din     (_zz_1208[35:0]        ), //i
    .dout    (fixTo_247_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_248 (
    .din     (_zz_1209[35:0]        ), //i
    .dout    (fixTo_248_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_249 (
    .din     (_zz_1210[35:0]        ), //i
    .dout    (fixTo_249_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_250 (
    .din     (_zz_1211[35:0]        ), //i
    .dout    (fixTo_250_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_251 (
    .din     (_zz_1212[35:0]        ), //i
    .dout    (fixTo_251_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_252 (
    .din     (_zz_1213[35:0]        ), //i
    .dout    (fixTo_252_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_253 (
    .din     (_zz_1214[35:0]        ), //i
    .dout    (fixTo_253_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_254 (
    .din     (_zz_1215[35:0]        ), //i
    .dout    (fixTo_254_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_255 (
    .din     (_zz_1216[35:0]        ), //i
    .dout    (fixTo_255_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_256 (
    .din     (_zz_1217[35:0]        ), //i
    .dout    (fixTo_256_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_257 (
    .din     (_zz_1218[35:0]        ), //i
    .dout    (fixTo_257_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_258 (
    .din     (_zz_1219[35:0]        ), //i
    .dout    (fixTo_258_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_259 (
    .din     (_zz_1220[35:0]        ), //i
    .dout    (fixTo_259_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_260 (
    .din     (_zz_1221[35:0]        ), //i
    .dout    (fixTo_260_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_261 (
    .din     (_zz_1222[35:0]        ), //i
    .dout    (fixTo_261_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_262 (
    .din     (_zz_1223[35:0]        ), //i
    .dout    (fixTo_262_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_263 (
    .din     (_zz_1224[35:0]        ), //i
    .dout    (fixTo_263_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_264 (
    .din     (_zz_1225[35:0]        ), //i
    .dout    (fixTo_264_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_265 (
    .din     (_zz_1226[35:0]        ), //i
    .dout    (fixTo_265_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_266 (
    .din     (_zz_1227[35:0]        ), //i
    .dout    (fixTo_266_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_267 (
    .din     (_zz_1228[35:0]        ), //i
    .dout    (fixTo_267_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_268 (
    .din     (_zz_1229[35:0]        ), //i
    .dout    (fixTo_268_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_269 (
    .din     (_zz_1230[35:0]        ), //i
    .dout    (fixTo_269_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_270 (
    .din     (_zz_1231[35:0]        ), //i
    .dout    (fixTo_270_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_271 (
    .din     (_zz_1232[35:0]        ), //i
    .dout    (fixTo_271_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_272 (
    .din     (_zz_1233[35:0]        ), //i
    .dout    (fixTo_272_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_273 (
    .din     (_zz_1234[35:0]        ), //i
    .dout    (fixTo_273_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_274 (
    .din     (_zz_1235[35:0]        ), //i
    .dout    (fixTo_274_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_275 (
    .din     (_zz_1236[35:0]        ), //i
    .dout    (fixTo_275_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_276 (
    .din     (_zz_1237[35:0]        ), //i
    .dout    (fixTo_276_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_277 (
    .din     (_zz_1238[35:0]        ), //i
    .dout    (fixTo_277_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_278 (
    .din     (_zz_1239[35:0]        ), //i
    .dout    (fixTo_278_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_279 (
    .din     (_zz_1240[35:0]        ), //i
    .dout    (fixTo_279_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_280 (
    .din     (_zz_1241[35:0]        ), //i
    .dout    (fixTo_280_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_281 (
    .din     (_zz_1242[35:0]        ), //i
    .dout    (fixTo_281_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_282 (
    .din     (_zz_1243[35:0]        ), //i
    .dout    (fixTo_282_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_283 (
    .din     (_zz_1244[35:0]        ), //i
    .dout    (fixTo_283_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_284 (
    .din     (_zz_1245[35:0]        ), //i
    .dout    (fixTo_284_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_285 (
    .din     (_zz_1246[35:0]        ), //i
    .dout    (fixTo_285_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_286 (
    .din     (_zz_1247[35:0]        ), //i
    .dout    (fixTo_286_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_287 (
    .din     (_zz_1248[35:0]        ), //i
    .dout    (fixTo_287_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_288 (
    .din     (_zz_1249[35:0]        ), //i
    .dout    (fixTo_288_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_289 (
    .din     (_zz_1250[35:0]        ), //i
    .dout    (fixTo_289_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_290 (
    .din     (_zz_1251[35:0]        ), //i
    .dout    (fixTo_290_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_291 (
    .din     (_zz_1252[35:0]        ), //i
    .dout    (fixTo_291_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_292 (
    .din     (_zz_1253[35:0]        ), //i
    .dout    (fixTo_292_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_293 (
    .din     (_zz_1254[35:0]        ), //i
    .dout    (fixTo_293_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_294 (
    .din     (_zz_1255[35:0]        ), //i
    .dout    (fixTo_294_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_295 (
    .din     (_zz_1256[35:0]        ), //i
    .dout    (fixTo_295_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_296 (
    .din     (_zz_1257[35:0]        ), //i
    .dout    (fixTo_296_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_297 (
    .din     (_zz_1258[35:0]        ), //i
    .dout    (fixTo_297_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_298 (
    .din     (_zz_1259[35:0]        ), //i
    .dout    (fixTo_298_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_299 (
    .din     (_zz_1260[35:0]        ), //i
    .dout    (fixTo_299_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_300 (
    .din     (_zz_1261[35:0]        ), //i
    .dout    (fixTo_300_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_301 (
    .din     (_zz_1262[35:0]        ), //i
    .dout    (fixTo_301_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_302 (
    .din     (_zz_1263[35:0]        ), //i
    .dout    (fixTo_302_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_303 (
    .din     (_zz_1264[35:0]        ), //i
    .dout    (fixTo_303_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_304 (
    .din     (_zz_1265[35:0]        ), //i
    .dout    (fixTo_304_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_305 (
    .din     (_zz_1266[35:0]        ), //i
    .dout    (fixTo_305_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_306 (
    .din     (_zz_1267[35:0]        ), //i
    .dout    (fixTo_306_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_307 (
    .din     (_zz_1268[35:0]        ), //i
    .dout    (fixTo_307_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_308 (
    .din     (_zz_1269[35:0]        ), //i
    .dout    (fixTo_308_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_309 (
    .din     (_zz_1270[35:0]        ), //i
    .dout    (fixTo_309_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_310 (
    .din     (_zz_1271[35:0]        ), //i
    .dout    (fixTo_310_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_311 (
    .din     (_zz_1272[35:0]        ), //i
    .dout    (fixTo_311_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_312 (
    .din     (_zz_1273[35:0]        ), //i
    .dout    (fixTo_312_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_313 (
    .din     (_zz_1274[35:0]        ), //i
    .dout    (fixTo_313_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_314 (
    .din     (_zz_1275[35:0]        ), //i
    .dout    (fixTo_314_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_315 (
    .din     (_zz_1276[35:0]        ), //i
    .dout    (fixTo_315_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_316 (
    .din     (_zz_1277[35:0]        ), //i
    .dout    (fixTo_316_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_317 (
    .din     (_zz_1278[35:0]        ), //i
    .dout    (fixTo_317_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_318 (
    .din     (_zz_1279[35:0]        ), //i
    .dout    (fixTo_318_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_319 (
    .din     (_zz_1280[35:0]        ), //i
    .dout    (fixTo_319_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_320 (
    .din     (_zz_1281[35:0]        ), //i
    .dout    (fixTo_320_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_321 (
    .din     (_zz_1282[35:0]        ), //i
    .dout    (fixTo_321_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_322 (
    .din     (_zz_1283[35:0]        ), //i
    .dout    (fixTo_322_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_323 (
    .din     (_zz_1284[35:0]        ), //i
    .dout    (fixTo_323_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_324 (
    .din     (_zz_1285[35:0]        ), //i
    .dout    (fixTo_324_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_325 (
    .din     (_zz_1286[35:0]        ), //i
    .dout    (fixTo_325_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_326 (
    .din     (_zz_1287[35:0]        ), //i
    .dout    (fixTo_326_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_327 (
    .din     (_zz_1288[35:0]        ), //i
    .dout    (fixTo_327_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_328 (
    .din     (_zz_1289[35:0]        ), //i
    .dout    (fixTo_328_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_329 (
    .din     (_zz_1290[35:0]        ), //i
    .dout    (fixTo_329_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_330 (
    .din     (_zz_1291[35:0]        ), //i
    .dout    (fixTo_330_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_331 (
    .din     (_zz_1292[35:0]        ), //i
    .dout    (fixTo_331_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_332 (
    .din     (_zz_1293[35:0]        ), //i
    .dout    (fixTo_332_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_333 (
    .din     (_zz_1294[35:0]        ), //i
    .dout    (fixTo_333_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_334 (
    .din     (_zz_1295[35:0]        ), //i
    .dout    (fixTo_334_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_335 (
    .din     (_zz_1296[35:0]        ), //i
    .dout    (fixTo_335_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_336 (
    .din     (_zz_1297[35:0]        ), //i
    .dout    (fixTo_336_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_337 (
    .din     (_zz_1298[35:0]        ), //i
    .dout    (fixTo_337_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_338 (
    .din     (_zz_1299[35:0]        ), //i
    .dout    (fixTo_338_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_339 (
    .din     (_zz_1300[35:0]        ), //i
    .dout    (fixTo_339_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_340 (
    .din     (_zz_1301[35:0]        ), //i
    .dout    (fixTo_340_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_341 (
    .din     (_zz_1302[35:0]        ), //i
    .dout    (fixTo_341_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_342 (
    .din     (_zz_1303[35:0]        ), //i
    .dout    (fixTo_342_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_343 (
    .din     (_zz_1304[35:0]        ), //i
    .dout    (fixTo_343_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_344 (
    .din     (_zz_1305[35:0]        ), //i
    .dout    (fixTo_344_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_345 (
    .din     (_zz_1306[35:0]        ), //i
    .dout    (fixTo_345_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_346 (
    .din     (_zz_1307[35:0]        ), //i
    .dout    (fixTo_346_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_347 (
    .din     (_zz_1308[35:0]        ), //i
    .dout    (fixTo_347_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_348 (
    .din     (_zz_1309[35:0]        ), //i
    .dout    (fixTo_348_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_349 (
    .din     (_zz_1310[35:0]        ), //i
    .dout    (fixTo_349_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_350 (
    .din     (_zz_1311[35:0]        ), //i
    .dout    (fixTo_350_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_351 (
    .din     (_zz_1312[35:0]        ), //i
    .dout    (fixTo_351_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_352 (
    .din     (_zz_1313[35:0]        ), //i
    .dout    (fixTo_352_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_353 (
    .din     (_zz_1314[35:0]        ), //i
    .dout    (fixTo_353_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_354 (
    .din     (_zz_1315[35:0]        ), //i
    .dout    (fixTo_354_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_355 (
    .din     (_zz_1316[35:0]        ), //i
    .dout    (fixTo_355_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_356 (
    .din     (_zz_1317[35:0]        ), //i
    .dout    (fixTo_356_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_357 (
    .din     (_zz_1318[35:0]        ), //i
    .dout    (fixTo_357_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_358 (
    .din     (_zz_1319[35:0]        ), //i
    .dout    (fixTo_358_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_359 (
    .din     (_zz_1320[35:0]        ), //i
    .dout    (fixTo_359_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_360 (
    .din     (_zz_1321[35:0]        ), //i
    .dout    (fixTo_360_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_361 (
    .din     (_zz_1322[35:0]        ), //i
    .dout    (fixTo_361_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_362 (
    .din     (_zz_1323[35:0]        ), //i
    .dout    (fixTo_362_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_363 (
    .din     (_zz_1324[35:0]        ), //i
    .dout    (fixTo_363_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_364 (
    .din     (_zz_1325[35:0]        ), //i
    .dout    (fixTo_364_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_365 (
    .din     (_zz_1326[35:0]        ), //i
    .dout    (fixTo_365_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_366 (
    .din     (_zz_1327[35:0]        ), //i
    .dout    (fixTo_366_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_367 (
    .din     (_zz_1328[35:0]        ), //i
    .dout    (fixTo_367_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_368 (
    .din     (_zz_1329[35:0]        ), //i
    .dout    (fixTo_368_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_369 (
    .din     (_zz_1330[35:0]        ), //i
    .dout    (fixTo_369_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_370 (
    .din     (_zz_1331[35:0]        ), //i
    .dout    (fixTo_370_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_371 (
    .din     (_zz_1332[35:0]        ), //i
    .dout    (fixTo_371_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_372 (
    .din     (_zz_1333[35:0]        ), //i
    .dout    (fixTo_372_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_373 (
    .din     (_zz_1334[35:0]        ), //i
    .dout    (fixTo_373_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_374 (
    .din     (_zz_1335[35:0]        ), //i
    .dout    (fixTo_374_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_375 (
    .din     (_zz_1336[35:0]        ), //i
    .dout    (fixTo_375_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_376 (
    .din     (_zz_1337[35:0]        ), //i
    .dout    (fixTo_376_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_377 (
    .din     (_zz_1338[35:0]        ), //i
    .dout    (fixTo_377_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_378 (
    .din     (_zz_1339[35:0]        ), //i
    .dout    (fixTo_378_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_379 (
    .din     (_zz_1340[35:0]        ), //i
    .dout    (fixTo_379_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_380 (
    .din     (_zz_1341[35:0]        ), //i
    .dout    (fixTo_380_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_381 (
    .din     (_zz_1342[35:0]        ), //i
    .dout    (fixTo_381_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_382 (
    .din     (_zz_1343[35:0]        ), //i
    .dout    (fixTo_382_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_383 (
    .din     (_zz_1344[35:0]        ), //i
    .dout    (fixTo_383_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_384 (
    .din     (_zz_1345[35:0]        ), //i
    .dout    (fixTo_384_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_385 (
    .din     (_zz_1346[35:0]        ), //i
    .dout    (fixTo_385_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_386 (
    .din     (_zz_1347[35:0]        ), //i
    .dout    (fixTo_386_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_387 (
    .din     (_zz_1348[35:0]        ), //i
    .dout    (fixTo_387_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_388 (
    .din     (_zz_1349[35:0]        ), //i
    .dout    (fixTo_388_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_389 (
    .din     (_zz_1350[35:0]        ), //i
    .dout    (fixTo_389_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_390 (
    .din     (_zz_1351[35:0]        ), //i
    .dout    (fixTo_390_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_391 (
    .din     (_zz_1352[35:0]        ), //i
    .dout    (fixTo_391_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_392 (
    .din     (_zz_1353[35:0]        ), //i
    .dout    (fixTo_392_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_393 (
    .din     (_zz_1354[35:0]        ), //i
    .dout    (fixTo_393_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_394 (
    .din     (_zz_1355[35:0]        ), //i
    .dout    (fixTo_394_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_395 (
    .din     (_zz_1356[35:0]        ), //i
    .dout    (fixTo_395_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_396 (
    .din     (_zz_1357[35:0]        ), //i
    .dout    (fixTo_396_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_397 (
    .din     (_zz_1358[35:0]        ), //i
    .dout    (fixTo_397_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_398 (
    .din     (_zz_1359[35:0]        ), //i
    .dout    (fixTo_398_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_399 (
    .din     (_zz_1360[35:0]        ), //i
    .dout    (fixTo_399_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_400 (
    .din     (_zz_1361[35:0]        ), //i
    .dout    (fixTo_400_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_401 (
    .din     (_zz_1362[35:0]        ), //i
    .dout    (fixTo_401_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_402 (
    .din     (_zz_1363[35:0]        ), //i
    .dout    (fixTo_402_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_403 (
    .din     (_zz_1364[35:0]        ), //i
    .dout    (fixTo_403_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_404 (
    .din     (_zz_1365[35:0]        ), //i
    .dout    (fixTo_404_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_405 (
    .din     (_zz_1366[35:0]        ), //i
    .dout    (fixTo_405_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_406 (
    .din     (_zz_1367[35:0]        ), //i
    .dout    (fixTo_406_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_407 (
    .din     (_zz_1368[35:0]        ), //i
    .dout    (fixTo_407_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_408 (
    .din     (_zz_1369[35:0]        ), //i
    .dout    (fixTo_408_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_409 (
    .din     (_zz_1370[35:0]        ), //i
    .dout    (fixTo_409_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_410 (
    .din     (_zz_1371[35:0]        ), //i
    .dout    (fixTo_410_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_411 (
    .din     (_zz_1372[35:0]        ), //i
    .dout    (fixTo_411_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_412 (
    .din     (_zz_1373[35:0]        ), //i
    .dout    (fixTo_412_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_413 (
    .din     (_zz_1374[35:0]        ), //i
    .dout    (fixTo_413_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_414 (
    .din     (_zz_1375[35:0]        ), //i
    .dout    (fixTo_414_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_415 (
    .din     (_zz_1376[35:0]        ), //i
    .dout    (fixTo_415_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_416 (
    .din     (_zz_1377[35:0]        ), //i
    .dout    (fixTo_416_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_417 (
    .din     (_zz_1378[35:0]        ), //i
    .dout    (fixTo_417_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_418 (
    .din     (_zz_1379[35:0]        ), //i
    .dout    (fixTo_418_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_419 (
    .din     (_zz_1380[35:0]        ), //i
    .dout    (fixTo_419_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_420 (
    .din     (_zz_1381[35:0]        ), //i
    .dout    (fixTo_420_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_421 (
    .din     (_zz_1382[35:0]        ), //i
    .dout    (fixTo_421_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_422 (
    .din     (_zz_1383[35:0]        ), //i
    .dout    (fixTo_422_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_423 (
    .din     (_zz_1384[35:0]        ), //i
    .dout    (fixTo_423_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_424 (
    .din     (_zz_1385[35:0]        ), //i
    .dout    (fixTo_424_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_425 (
    .din     (_zz_1386[35:0]        ), //i
    .dout    (fixTo_425_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_426 (
    .din     (_zz_1387[35:0]        ), //i
    .dout    (fixTo_426_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_427 (
    .din     (_zz_1388[35:0]        ), //i
    .dout    (fixTo_427_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_428 (
    .din     (_zz_1389[35:0]        ), //i
    .dout    (fixTo_428_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_429 (
    .din     (_zz_1390[35:0]        ), //i
    .dout    (fixTo_429_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_430 (
    .din     (_zz_1391[35:0]        ), //i
    .dout    (fixTo_430_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_431 (
    .din     (_zz_1392[35:0]        ), //i
    .dout    (fixTo_431_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_432 (
    .din     (_zz_1393[35:0]        ), //i
    .dout    (fixTo_432_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_433 (
    .din     (_zz_1394[35:0]        ), //i
    .dout    (fixTo_433_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_434 (
    .din     (_zz_1395[35:0]        ), //i
    .dout    (fixTo_434_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_435 (
    .din     (_zz_1396[35:0]        ), //i
    .dout    (fixTo_435_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_436 (
    .din     (_zz_1397[35:0]        ), //i
    .dout    (fixTo_436_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_437 (
    .din     (_zz_1398[35:0]        ), //i
    .dout    (fixTo_437_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_438 (
    .din     (_zz_1399[35:0]        ), //i
    .dout    (fixTo_438_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_439 (
    .din     (_zz_1400[35:0]        ), //i
    .dout    (fixTo_439_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_440 (
    .din     (_zz_1401[35:0]        ), //i
    .dout    (fixTo_440_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_441 (
    .din     (_zz_1402[35:0]        ), //i
    .dout    (fixTo_441_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_442 (
    .din     (_zz_1403[35:0]        ), //i
    .dout    (fixTo_442_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_443 (
    .din     (_zz_1404[35:0]        ), //i
    .dout    (fixTo_443_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_444 (
    .din     (_zz_1405[35:0]        ), //i
    .dout    (fixTo_444_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_445 (
    .din     (_zz_1406[35:0]        ), //i
    .dout    (fixTo_445_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_446 (
    .din     (_zz_1407[35:0]        ), //i
    .dout    (fixTo_446_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_447 (
    .din     (_zz_1408[35:0]        ), //i
    .dout    (fixTo_447_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_448 (
    .din     (_zz_1409[35:0]        ), //i
    .dout    (fixTo_448_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_449 (
    .din     (_zz_1410[35:0]        ), //i
    .dout    (fixTo_449_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_450 (
    .din     (_zz_1411[35:0]        ), //i
    .dout    (fixTo_450_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_451 (
    .din     (_zz_1412[35:0]        ), //i
    .dout    (fixTo_451_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_452 (
    .din     (_zz_1413[35:0]        ), //i
    .dout    (fixTo_452_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_453 (
    .din     (_zz_1414[35:0]        ), //i
    .dout    (fixTo_453_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_454 (
    .din     (_zz_1415[35:0]        ), //i
    .dout    (fixTo_454_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_455 (
    .din     (_zz_1416[35:0]        ), //i
    .dout    (fixTo_455_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_456 (
    .din     (_zz_1417[35:0]        ), //i
    .dout    (fixTo_456_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_457 (
    .din     (_zz_1418[35:0]        ), //i
    .dout    (fixTo_457_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_458 (
    .din     (_zz_1419[35:0]        ), //i
    .dout    (fixTo_458_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_459 (
    .din     (_zz_1420[35:0]        ), //i
    .dout    (fixTo_459_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_460 (
    .din     (_zz_1421[35:0]        ), //i
    .dout    (fixTo_460_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_461 (
    .din     (_zz_1422[35:0]        ), //i
    .dout    (fixTo_461_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_462 (
    .din     (_zz_1423[35:0]        ), //i
    .dout    (fixTo_462_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_463 (
    .din     (_zz_1424[35:0]        ), //i
    .dout    (fixTo_463_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_464 (
    .din     (_zz_1425[35:0]        ), //i
    .dout    (fixTo_464_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_465 (
    .din     (_zz_1426[35:0]        ), //i
    .dout    (fixTo_465_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_466 (
    .din     (_zz_1427[35:0]        ), //i
    .dout    (fixTo_466_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_467 (
    .din     (_zz_1428[35:0]        ), //i
    .dout    (fixTo_467_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_468 (
    .din     (_zz_1429[35:0]        ), //i
    .dout    (fixTo_468_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_469 (
    .din     (_zz_1430[35:0]        ), //i
    .dout    (fixTo_469_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_470 (
    .din     (_zz_1431[35:0]        ), //i
    .dout    (fixTo_470_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_471 (
    .din     (_zz_1432[35:0]        ), //i
    .dout    (fixTo_471_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_472 (
    .din     (_zz_1433[35:0]        ), //i
    .dout    (fixTo_472_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_473 (
    .din     (_zz_1434[35:0]        ), //i
    .dout    (fixTo_473_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_474 (
    .din     (_zz_1435[35:0]        ), //i
    .dout    (fixTo_474_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_475 (
    .din     (_zz_1436[35:0]        ), //i
    .dout    (fixTo_475_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_476 (
    .din     (_zz_1437[35:0]        ), //i
    .dout    (fixTo_476_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_477 (
    .din     (_zz_1438[35:0]        ), //i
    .dout    (fixTo_477_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_478 (
    .din     (_zz_1439[35:0]        ), //i
    .dout    (fixTo_478_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_479 (
    .din     (_zz_1440[35:0]        ), //i
    .dout    (fixTo_479_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_480 (
    .din     (_zz_1441[35:0]        ), //i
    .dout    (fixTo_480_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_481 (
    .din     (_zz_1442[35:0]        ), //i
    .dout    (fixTo_481_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_482 (
    .din     (_zz_1443[35:0]        ), //i
    .dout    (fixTo_482_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_483 (
    .din     (_zz_1444[35:0]        ), //i
    .dout    (fixTo_483_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_484 (
    .din     (_zz_1445[35:0]        ), //i
    .dout    (fixTo_484_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_485 (
    .din     (_zz_1446[35:0]        ), //i
    .dout    (fixTo_485_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_486 (
    .din     (_zz_1447[35:0]        ), //i
    .dout    (fixTo_486_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_487 (
    .din     (_zz_1448[35:0]        ), //i
    .dout    (fixTo_487_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_488 (
    .din     (_zz_1449[35:0]        ), //i
    .dout    (fixTo_488_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_489 (
    .din     (_zz_1450[35:0]        ), //i
    .dout    (fixTo_489_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_490 (
    .din     (_zz_1451[35:0]        ), //i
    .dout    (fixTo_490_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_491 (
    .din     (_zz_1452[35:0]        ), //i
    .dout    (fixTo_491_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_492 (
    .din     (_zz_1453[35:0]        ), //i
    .dout    (fixTo_492_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_493 (
    .din     (_zz_1454[35:0]        ), //i
    .dout    (fixTo_493_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_494 (
    .din     (_zz_1455[35:0]        ), //i
    .dout    (fixTo_494_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_495 (
    .din     (_zz_1456[35:0]        ), //i
    .dout    (fixTo_495_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_496 (
    .din     (_zz_1457[35:0]        ), //i
    .dout    (fixTo_496_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_497 (
    .din     (_zz_1458[35:0]        ), //i
    .dout    (fixTo_497_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_498 (
    .din     (_zz_1459[35:0]        ), //i
    .dout    (fixTo_498_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_499 (
    .din     (_zz_1460[35:0]        ), //i
    .dout    (fixTo_499_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_500 (
    .din     (_zz_1461[35:0]        ), //i
    .dout    (fixTo_500_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_501 (
    .din     (_zz_1462[35:0]        ), //i
    .dout    (fixTo_501_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_502 (
    .din     (_zz_1463[35:0]        ), //i
    .dout    (fixTo_502_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_503 (
    .din     (_zz_1464[35:0]        ), //i
    .dout    (fixTo_503_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_504 (
    .din     (_zz_1465[35:0]        ), //i
    .dout    (fixTo_504_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_505 (
    .din     (_zz_1466[35:0]        ), //i
    .dout    (fixTo_505_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_506 (
    .din     (_zz_1467[35:0]        ), //i
    .dout    (fixTo_506_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_507 (
    .din     (_zz_1468[35:0]        ), //i
    .dout    (fixTo_507_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_508 (
    .din     (_zz_1469[35:0]        ), //i
    .dout    (fixTo_508_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_509 (
    .din     (_zz_1470[35:0]        ), //i
    .dout    (fixTo_509_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_510 (
    .din     (_zz_1471[35:0]        ), //i
    .dout    (fixTo_510_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_511 (
    .din     (_zz_1472[35:0]        ), //i
    .dout    (fixTo_511_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_512 (
    .din     (_zz_1473[35:0]        ), //i
    .dout    (fixTo_512_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_513 (
    .din     (_zz_1474[35:0]        ), //i
    .dout    (fixTo_513_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_514 (
    .din     (_zz_1475[35:0]        ), //i
    .dout    (fixTo_514_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_515 (
    .din     (_zz_1476[35:0]        ), //i
    .dout    (fixTo_515_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_516 (
    .din     (_zz_1477[35:0]        ), //i
    .dout    (fixTo_516_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_517 (
    .din     (_zz_1478[35:0]        ), //i
    .dout    (fixTo_517_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_518 (
    .din     (_zz_1479[35:0]        ), //i
    .dout    (fixTo_518_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_519 (
    .din     (_zz_1480[35:0]        ), //i
    .dout    (fixTo_519_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_520 (
    .din     (_zz_1481[35:0]        ), //i
    .dout    (fixTo_520_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_521 (
    .din     (_zz_1482[35:0]        ), //i
    .dout    (fixTo_521_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_522 (
    .din     (_zz_1483[35:0]        ), //i
    .dout    (fixTo_522_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_523 (
    .din     (_zz_1484[35:0]        ), //i
    .dout    (fixTo_523_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_524 (
    .din     (_zz_1485[35:0]        ), //i
    .dout    (fixTo_524_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_525 (
    .din     (_zz_1486[35:0]        ), //i
    .dout    (fixTo_525_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_526 (
    .din     (_zz_1487[35:0]        ), //i
    .dout    (fixTo_526_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_527 (
    .din     (_zz_1488[35:0]        ), //i
    .dout    (fixTo_527_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_528 (
    .din     (_zz_1489[35:0]        ), //i
    .dout    (fixTo_528_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_529 (
    .din     (_zz_1490[35:0]        ), //i
    .dout    (fixTo_529_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_530 (
    .din     (_zz_1491[35:0]        ), //i
    .dout    (fixTo_530_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_531 (
    .din     (_zz_1492[35:0]        ), //i
    .dout    (fixTo_531_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_532 (
    .din     (_zz_1493[35:0]        ), //i
    .dout    (fixTo_532_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_533 (
    .din     (_zz_1494[35:0]        ), //i
    .dout    (fixTo_533_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_534 (
    .din     (_zz_1495[35:0]        ), //i
    .dout    (fixTo_534_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_535 (
    .din     (_zz_1496[35:0]        ), //i
    .dout    (fixTo_535_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_536 (
    .din     (_zz_1497[35:0]        ), //i
    .dout    (fixTo_536_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_537 (
    .din     (_zz_1498[35:0]        ), //i
    .dout    (fixTo_537_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_538 (
    .din     (_zz_1499[35:0]        ), //i
    .dout    (fixTo_538_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_539 (
    .din     (_zz_1500[35:0]        ), //i
    .dout    (fixTo_539_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_540 (
    .din     (_zz_1501[35:0]        ), //i
    .dout    (fixTo_540_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_541 (
    .din     (_zz_1502[35:0]        ), //i
    .dout    (fixTo_541_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_542 (
    .din     (_zz_1503[35:0]        ), //i
    .dout    (fixTo_542_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_543 (
    .din     (_zz_1504[35:0]        ), //i
    .dout    (fixTo_543_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_544 (
    .din     (_zz_1505[35:0]        ), //i
    .dout    (fixTo_544_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_545 (
    .din     (_zz_1506[35:0]        ), //i
    .dout    (fixTo_545_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_546 (
    .din     (_zz_1507[35:0]        ), //i
    .dout    (fixTo_546_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_547 (
    .din     (_zz_1508[35:0]        ), //i
    .dout    (fixTo_547_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_548 (
    .din     (_zz_1509[35:0]        ), //i
    .dout    (fixTo_548_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_549 (
    .din     (_zz_1510[35:0]        ), //i
    .dout    (fixTo_549_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_550 (
    .din     (_zz_1511[35:0]        ), //i
    .dout    (fixTo_550_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_551 (
    .din     (_zz_1512[35:0]        ), //i
    .dout    (fixTo_551_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_552 (
    .din     (_zz_1513[35:0]        ), //i
    .dout    (fixTo_552_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_553 (
    .din     (_zz_1514[35:0]        ), //i
    .dout    (fixTo_553_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_554 (
    .din     (_zz_1515[35:0]        ), //i
    .dout    (fixTo_554_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_555 (
    .din     (_zz_1516[35:0]        ), //i
    .dout    (fixTo_555_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_556 (
    .din     (_zz_1517[35:0]        ), //i
    .dout    (fixTo_556_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_557 (
    .din     (_zz_1518[35:0]        ), //i
    .dout    (fixTo_557_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_558 (
    .din     (_zz_1519[35:0]        ), //i
    .dout    (fixTo_558_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_559 (
    .din     (_zz_1520[35:0]        ), //i
    .dout    (fixTo_559_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_560 (
    .din     (_zz_1521[35:0]        ), //i
    .dout    (fixTo_560_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_561 (
    .din     (_zz_1522[35:0]        ), //i
    .dout    (fixTo_561_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_562 (
    .din     (_zz_1523[35:0]        ), //i
    .dout    (fixTo_562_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_563 (
    .din     (_zz_1524[35:0]        ), //i
    .dout    (fixTo_563_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_564 (
    .din     (_zz_1525[35:0]        ), //i
    .dout    (fixTo_564_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_565 (
    .din     (_zz_1526[35:0]        ), //i
    .dout    (fixTo_565_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_566 (
    .din     (_zz_1527[35:0]        ), //i
    .dout    (fixTo_566_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_567 (
    .din     (_zz_1528[35:0]        ), //i
    .dout    (fixTo_567_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_568 (
    .din     (_zz_1529[35:0]        ), //i
    .dout    (fixTo_568_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_569 (
    .din     (_zz_1530[35:0]        ), //i
    .dout    (fixTo_569_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_570 (
    .din     (_zz_1531[35:0]        ), //i
    .dout    (fixTo_570_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_571 (
    .din     (_zz_1532[35:0]        ), //i
    .dout    (fixTo_571_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_572 (
    .din     (_zz_1533[35:0]        ), //i
    .dout    (fixTo_572_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_573 (
    .din     (_zz_1534[35:0]        ), //i
    .dout    (fixTo_573_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_574 (
    .din     (_zz_1535[35:0]        ), //i
    .dout    (fixTo_574_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_575 (
    .din     (_zz_1536[35:0]        ), //i
    .dout    (fixTo_575_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_576 (
    .din     (_zz_1537[35:0]        ), //i
    .dout    (fixTo_576_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_577 (
    .din     (_zz_1538[35:0]        ), //i
    .dout    (fixTo_577_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_578 (
    .din     (_zz_1539[35:0]        ), //i
    .dout    (fixTo_578_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_579 (
    .din     (_zz_1540[35:0]        ), //i
    .dout    (fixTo_579_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_580 (
    .din     (_zz_1541[35:0]        ), //i
    .dout    (fixTo_580_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_581 (
    .din     (_zz_1542[35:0]        ), //i
    .dout    (fixTo_581_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_582 (
    .din     (_zz_1543[35:0]        ), //i
    .dout    (fixTo_582_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_583 (
    .din     (_zz_1544[35:0]        ), //i
    .dout    (fixTo_583_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_584 (
    .din     (_zz_1545[35:0]        ), //i
    .dout    (fixTo_584_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_585 (
    .din     (_zz_1546[35:0]        ), //i
    .dout    (fixTo_585_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_586 (
    .din     (_zz_1547[35:0]        ), //i
    .dout    (fixTo_586_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_587 (
    .din     (_zz_1548[35:0]        ), //i
    .dout    (fixTo_587_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_588 (
    .din     (_zz_1549[35:0]        ), //i
    .dout    (fixTo_588_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_589 (
    .din     (_zz_1550[35:0]        ), //i
    .dout    (fixTo_589_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_590 (
    .din     (_zz_1551[35:0]        ), //i
    .dout    (fixTo_590_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_591 (
    .din     (_zz_1552[35:0]        ), //i
    .dout    (fixTo_591_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_592 (
    .din     (_zz_1553[35:0]        ), //i
    .dout    (fixTo_592_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_593 (
    .din     (_zz_1554[35:0]        ), //i
    .dout    (fixTo_593_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_594 (
    .din     (_zz_1555[35:0]        ), //i
    .dout    (fixTo_594_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_595 (
    .din     (_zz_1556[35:0]        ), //i
    .dout    (fixTo_595_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_596 (
    .din     (_zz_1557[35:0]        ), //i
    .dout    (fixTo_596_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_597 (
    .din     (_zz_1558[35:0]        ), //i
    .dout    (fixTo_597_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_598 (
    .din     (_zz_1559[35:0]        ), //i
    .dout    (fixTo_598_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_599 (
    .din     (_zz_1560[35:0]        ), //i
    .dout    (fixTo_599_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_600 (
    .din     (_zz_1561[35:0]        ), //i
    .dout    (fixTo_600_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_601 (
    .din     (_zz_1562[35:0]        ), //i
    .dout    (fixTo_601_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_602 (
    .din     (_zz_1563[35:0]        ), //i
    .dout    (fixTo_602_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_603 (
    .din     (_zz_1564[35:0]        ), //i
    .dout    (fixTo_603_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_604 (
    .din     (_zz_1565[35:0]        ), //i
    .dout    (fixTo_604_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_605 (
    .din     (_zz_1566[35:0]        ), //i
    .dout    (fixTo_605_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_606 (
    .din     (_zz_1567[35:0]        ), //i
    .dout    (fixTo_606_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_607 (
    .din     (_zz_1568[35:0]        ), //i
    .dout    (fixTo_607_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_608 (
    .din     (_zz_1569[35:0]        ), //i
    .dout    (fixTo_608_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_609 (
    .din     (_zz_1570[35:0]        ), //i
    .dout    (fixTo_609_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_610 (
    .din     (_zz_1571[35:0]        ), //i
    .dout    (fixTo_610_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_611 (
    .din     (_zz_1572[35:0]        ), //i
    .dout    (fixTo_611_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_612 (
    .din     (_zz_1573[35:0]        ), //i
    .dout    (fixTo_612_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_613 (
    .din     (_zz_1574[35:0]        ), //i
    .dout    (fixTo_613_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_614 (
    .din     (_zz_1575[35:0]        ), //i
    .dout    (fixTo_614_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_615 (
    .din     (_zz_1576[35:0]        ), //i
    .dout    (fixTo_615_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_616 (
    .din     (_zz_1577[35:0]        ), //i
    .dout    (fixTo_616_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_617 (
    .din     (_zz_1578[35:0]        ), //i
    .dout    (fixTo_617_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_618 (
    .din     (_zz_1579[35:0]        ), //i
    .dout    (fixTo_618_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_619 (
    .din     (_zz_1580[35:0]        ), //i
    .dout    (fixTo_619_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_620 (
    .din     (_zz_1581[35:0]        ), //i
    .dout    (fixTo_620_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_621 (
    .din     (_zz_1582[35:0]        ), //i
    .dout    (fixTo_621_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_622 (
    .din     (_zz_1583[35:0]        ), //i
    .dout    (fixTo_622_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_623 (
    .din     (_zz_1584[35:0]        ), //i
    .dout    (fixTo_623_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_624 (
    .din     (_zz_1585[35:0]        ), //i
    .dout    (fixTo_624_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_625 (
    .din     (_zz_1586[35:0]        ), //i
    .dout    (fixTo_625_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_626 (
    .din     (_zz_1587[35:0]        ), //i
    .dout    (fixTo_626_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_627 (
    .din     (_zz_1588[35:0]        ), //i
    .dout    (fixTo_627_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_628 (
    .din     (_zz_1589[35:0]        ), //i
    .dout    (fixTo_628_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_629 (
    .din     (_zz_1590[35:0]        ), //i
    .dout    (fixTo_629_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_630 (
    .din     (_zz_1591[35:0]        ), //i
    .dout    (fixTo_630_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_631 (
    .din     (_zz_1592[35:0]        ), //i
    .dout    (fixTo_631_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_632 (
    .din     (_zz_1593[35:0]        ), //i
    .dout    (fixTo_632_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_633 (
    .din     (_zz_1594[35:0]        ), //i
    .dout    (fixTo_633_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_634 (
    .din     (_zz_1595[35:0]        ), //i
    .dout    (fixTo_634_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_635 (
    .din     (_zz_1596[35:0]        ), //i
    .dout    (fixTo_635_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_636 (
    .din     (_zz_1597[35:0]        ), //i
    .dout    (fixTo_636_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_637 (
    .din     (_zz_1598[35:0]        ), //i
    .dout    (fixTo_637_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_638 (
    .din     (_zz_1599[35:0]        ), //i
    .dout    (fixTo_638_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_639 (
    .din     (_zz_1600[35:0]        ), //i
    .dout    (fixTo_639_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_640 (
    .din     (_zz_1601[35:0]        ), //i
    .dout    (fixTo_640_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_641 (
    .din     (_zz_1602[35:0]        ), //i
    .dout    (fixTo_641_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_642 (
    .din     (_zz_1603[35:0]        ), //i
    .dout    (fixTo_642_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_643 (
    .din     (_zz_1604[35:0]        ), //i
    .dout    (fixTo_643_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_644 (
    .din     (_zz_1605[35:0]        ), //i
    .dout    (fixTo_644_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_645 (
    .din     (_zz_1606[35:0]        ), //i
    .dout    (fixTo_645_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_646 (
    .din     (_zz_1607[35:0]        ), //i
    .dout    (fixTo_646_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_647 (
    .din     (_zz_1608[35:0]        ), //i
    .dout    (fixTo_647_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_648 (
    .din     (_zz_1609[35:0]        ), //i
    .dout    (fixTo_648_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_649 (
    .din     (_zz_1610[35:0]        ), //i
    .dout    (fixTo_649_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_650 (
    .din     (_zz_1611[35:0]        ), //i
    .dout    (fixTo_650_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_651 (
    .din     (_zz_1612[35:0]        ), //i
    .dout    (fixTo_651_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_652 (
    .din     (_zz_1613[35:0]        ), //i
    .dout    (fixTo_652_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_653 (
    .din     (_zz_1614[35:0]        ), //i
    .dout    (fixTo_653_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_654 (
    .din     (_zz_1615[35:0]        ), //i
    .dout    (fixTo_654_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_655 (
    .din     (_zz_1616[35:0]        ), //i
    .dout    (fixTo_655_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_656 (
    .din     (_zz_1617[35:0]        ), //i
    .dout    (fixTo_656_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_657 (
    .din     (_zz_1618[35:0]        ), //i
    .dout    (fixTo_657_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_658 (
    .din     (_zz_1619[35:0]        ), //i
    .dout    (fixTo_658_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_659 (
    .din     (_zz_1620[35:0]        ), //i
    .dout    (fixTo_659_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_660 (
    .din     (_zz_1621[35:0]        ), //i
    .dout    (fixTo_660_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_661 (
    .din     (_zz_1622[35:0]        ), //i
    .dout    (fixTo_661_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_662 (
    .din     (_zz_1623[35:0]        ), //i
    .dout    (fixTo_662_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_663 (
    .din     (_zz_1624[35:0]        ), //i
    .dout    (fixTo_663_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_664 (
    .din     (_zz_1625[35:0]        ), //i
    .dout    (fixTo_664_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_665 (
    .din     (_zz_1626[35:0]        ), //i
    .dout    (fixTo_665_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_666 (
    .din     (_zz_1627[35:0]        ), //i
    .dout    (fixTo_666_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_667 (
    .din     (_zz_1628[35:0]        ), //i
    .dout    (fixTo_667_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_668 (
    .din     (_zz_1629[35:0]        ), //i
    .dout    (fixTo_668_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_669 (
    .din     (_zz_1630[35:0]        ), //i
    .dout    (fixTo_669_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_670 (
    .din     (_zz_1631[35:0]        ), //i
    .dout    (fixTo_670_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_671 (
    .din     (_zz_1632[35:0]        ), //i
    .dout    (fixTo_671_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_672 (
    .din     (_zz_1633[35:0]        ), //i
    .dout    (fixTo_672_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_673 (
    .din     (_zz_1634[35:0]        ), //i
    .dout    (fixTo_673_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_674 (
    .din     (_zz_1635[35:0]        ), //i
    .dout    (fixTo_674_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_675 (
    .din     (_zz_1636[35:0]        ), //i
    .dout    (fixTo_675_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_676 (
    .din     (_zz_1637[35:0]        ), //i
    .dout    (fixTo_676_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_677 (
    .din     (_zz_1638[35:0]        ), //i
    .dout    (fixTo_677_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_678 (
    .din     (_zz_1639[35:0]        ), //i
    .dout    (fixTo_678_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_679 (
    .din     (_zz_1640[35:0]        ), //i
    .dout    (fixTo_679_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_680 (
    .din     (_zz_1641[35:0]        ), //i
    .dout    (fixTo_680_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_681 (
    .din     (_zz_1642[35:0]        ), //i
    .dout    (fixTo_681_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_682 (
    .din     (_zz_1643[35:0]        ), //i
    .dout    (fixTo_682_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_683 (
    .din     (_zz_1644[35:0]        ), //i
    .dout    (fixTo_683_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_684 (
    .din     (_zz_1645[35:0]        ), //i
    .dout    (fixTo_684_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_685 (
    .din     (_zz_1646[35:0]        ), //i
    .dout    (fixTo_685_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_686 (
    .din     (_zz_1647[35:0]        ), //i
    .dout    (fixTo_686_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_687 (
    .din     (_zz_1648[35:0]        ), //i
    .dout    (fixTo_687_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_688 (
    .din     (_zz_1649[35:0]        ), //i
    .dout    (fixTo_688_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_689 (
    .din     (_zz_1650[35:0]        ), //i
    .dout    (fixTo_689_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_690 (
    .din     (_zz_1651[35:0]        ), //i
    .dout    (fixTo_690_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_691 (
    .din     (_zz_1652[35:0]        ), //i
    .dout    (fixTo_691_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_692 (
    .din     (_zz_1653[35:0]        ), //i
    .dout    (fixTo_692_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_693 (
    .din     (_zz_1654[35:0]        ), //i
    .dout    (fixTo_693_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_694 (
    .din     (_zz_1655[35:0]        ), //i
    .dout    (fixTo_694_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_695 (
    .din     (_zz_1656[35:0]        ), //i
    .dout    (fixTo_695_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_696 (
    .din     (_zz_1657[35:0]        ), //i
    .dout    (fixTo_696_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_697 (
    .din     (_zz_1658[35:0]        ), //i
    .dout    (fixTo_697_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_698 (
    .din     (_zz_1659[35:0]        ), //i
    .dout    (fixTo_698_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_699 (
    .din     (_zz_1660[35:0]        ), //i
    .dout    (fixTo_699_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_700 (
    .din     (_zz_1661[35:0]        ), //i
    .dout    (fixTo_700_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_701 (
    .din     (_zz_1662[35:0]        ), //i
    .dout    (fixTo_701_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_702 (
    .din     (_zz_1663[35:0]        ), //i
    .dout    (fixTo_702_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_703 (
    .din     (_zz_1664[35:0]        ), //i
    .dout    (fixTo_703_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_704 (
    .din     (_zz_1665[35:0]        ), //i
    .dout    (fixTo_704_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_705 (
    .din     (_zz_1666[35:0]        ), //i
    .dout    (fixTo_705_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_706 (
    .din     (_zz_1667[35:0]        ), //i
    .dout    (fixTo_706_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_707 (
    .din     (_zz_1668[35:0]        ), //i
    .dout    (fixTo_707_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_708 (
    .din     (_zz_1669[35:0]        ), //i
    .dout    (fixTo_708_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_709 (
    .din     (_zz_1670[35:0]        ), //i
    .dout    (fixTo_709_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_710 (
    .din     (_zz_1671[35:0]        ), //i
    .dout    (fixTo_710_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_711 (
    .din     (_zz_1672[35:0]        ), //i
    .dout    (fixTo_711_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_712 (
    .din     (_zz_1673[35:0]        ), //i
    .dout    (fixTo_712_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_713 (
    .din     (_zz_1674[35:0]        ), //i
    .dout    (fixTo_713_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_714 (
    .din     (_zz_1675[35:0]        ), //i
    .dout    (fixTo_714_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_715 (
    .din     (_zz_1676[35:0]        ), //i
    .dout    (fixTo_715_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_716 (
    .din     (_zz_1677[35:0]        ), //i
    .dout    (fixTo_716_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_717 (
    .din     (_zz_1678[35:0]        ), //i
    .dout    (fixTo_717_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_718 (
    .din     (_zz_1679[35:0]        ), //i
    .dout    (fixTo_718_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_719 (
    .din     (_zz_1680[35:0]        ), //i
    .dout    (fixTo_719_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_720 (
    .din     (_zz_1681[35:0]        ), //i
    .dout    (fixTo_720_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_721 (
    .din     (_zz_1682[35:0]        ), //i
    .dout    (fixTo_721_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_722 (
    .din     (_zz_1683[35:0]        ), //i
    .dout    (fixTo_722_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_723 (
    .din     (_zz_1684[35:0]        ), //i
    .dout    (fixTo_723_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_724 (
    .din     (_zz_1685[35:0]        ), //i
    .dout    (fixTo_724_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_725 (
    .din     (_zz_1686[35:0]        ), //i
    .dout    (fixTo_725_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_726 (
    .din     (_zz_1687[35:0]        ), //i
    .dout    (fixTo_726_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_727 (
    .din     (_zz_1688[35:0]        ), //i
    .dout    (fixTo_727_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_728 (
    .din     (_zz_1689[35:0]        ), //i
    .dout    (fixTo_728_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_729 (
    .din     (_zz_1690[35:0]        ), //i
    .dout    (fixTo_729_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_730 (
    .din     (_zz_1691[35:0]        ), //i
    .dout    (fixTo_730_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_731 (
    .din     (_zz_1692[35:0]        ), //i
    .dout    (fixTo_731_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_732 (
    .din     (_zz_1693[35:0]        ), //i
    .dout    (fixTo_732_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_733 (
    .din     (_zz_1694[35:0]        ), //i
    .dout    (fixTo_733_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_734 (
    .din     (_zz_1695[35:0]        ), //i
    .dout    (fixTo_734_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_735 (
    .din     (_zz_1696[35:0]        ), //i
    .dout    (fixTo_735_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_736 (
    .din     (_zz_1697[35:0]        ), //i
    .dout    (fixTo_736_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_737 (
    .din     (_zz_1698[35:0]        ), //i
    .dout    (fixTo_737_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_738 (
    .din     (_zz_1699[35:0]        ), //i
    .dout    (fixTo_738_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_739 (
    .din     (_zz_1700[35:0]        ), //i
    .dout    (fixTo_739_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_740 (
    .din     (_zz_1701[35:0]        ), //i
    .dout    (fixTo_740_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_741 (
    .din     (_zz_1702[35:0]        ), //i
    .dout    (fixTo_741_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_742 (
    .din     (_zz_1703[35:0]        ), //i
    .dout    (fixTo_742_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_743 (
    .din     (_zz_1704[35:0]        ), //i
    .dout    (fixTo_743_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_744 (
    .din     (_zz_1705[35:0]        ), //i
    .dout    (fixTo_744_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_745 (
    .din     (_zz_1706[35:0]        ), //i
    .dout    (fixTo_745_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_746 (
    .din     (_zz_1707[35:0]        ), //i
    .dout    (fixTo_746_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_747 (
    .din     (_zz_1708[35:0]        ), //i
    .dout    (fixTo_747_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_748 (
    .din     (_zz_1709[35:0]        ), //i
    .dout    (fixTo_748_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_749 (
    .din     (_zz_1710[35:0]        ), //i
    .dout    (fixTo_749_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_750 (
    .din     (_zz_1711[35:0]        ), //i
    .dout    (fixTo_750_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_751 (
    .din     (_zz_1712[35:0]        ), //i
    .dout    (fixTo_751_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_752 (
    .din     (_zz_1713[35:0]        ), //i
    .dout    (fixTo_752_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_753 (
    .din     (_zz_1714[35:0]        ), //i
    .dout    (fixTo_753_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_754 (
    .din     (_zz_1715[35:0]        ), //i
    .dout    (fixTo_754_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_755 (
    .din     (_zz_1716[35:0]        ), //i
    .dout    (fixTo_755_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_756 (
    .din     (_zz_1717[35:0]        ), //i
    .dout    (fixTo_756_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_757 (
    .din     (_zz_1718[35:0]        ), //i
    .dout    (fixTo_757_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_758 (
    .din     (_zz_1719[35:0]        ), //i
    .dout    (fixTo_758_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_759 (
    .din     (_zz_1720[35:0]        ), //i
    .dout    (fixTo_759_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_760 (
    .din     (_zz_1721[35:0]        ), //i
    .dout    (fixTo_760_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_761 (
    .din     (_zz_1722[35:0]        ), //i
    .dout    (fixTo_761_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_762 (
    .din     (_zz_1723[35:0]        ), //i
    .dout    (fixTo_762_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_763 (
    .din     (_zz_1724[35:0]        ), //i
    .dout    (fixTo_763_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_764 (
    .din     (_zz_1725[35:0]        ), //i
    .dout    (fixTo_764_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_765 (
    .din     (_zz_1726[35:0]        ), //i
    .dout    (fixTo_765_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_766 (
    .din     (_zz_1727[35:0]        ), //i
    .dout    (fixTo_766_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_767 (
    .din     (_zz_1728[35:0]        ), //i
    .dout    (fixTo_767_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_768 (
    .din     (_zz_1729[35:0]        ), //i
    .dout    (fixTo_768_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_769 (
    .din     (_zz_1730[35:0]        ), //i
    .dout    (fixTo_769_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_770 (
    .din     (_zz_1731[35:0]        ), //i
    .dout    (fixTo_770_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_771 (
    .din     (_zz_1732[35:0]        ), //i
    .dout    (fixTo_771_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_772 (
    .din     (_zz_1733[35:0]        ), //i
    .dout    (fixTo_772_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_773 (
    .din     (_zz_1734[35:0]        ), //i
    .dout    (fixTo_773_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_774 (
    .din     (_zz_1735[35:0]        ), //i
    .dout    (fixTo_774_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_775 (
    .din     (_zz_1736[35:0]        ), //i
    .dout    (fixTo_775_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_776 (
    .din     (_zz_1737[35:0]        ), //i
    .dout    (fixTo_776_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_777 (
    .din     (_zz_1738[35:0]        ), //i
    .dout    (fixTo_777_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_778 (
    .din     (_zz_1739[35:0]        ), //i
    .dout    (fixTo_778_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_779 (
    .din     (_zz_1740[35:0]        ), //i
    .dout    (fixTo_779_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_780 (
    .din     (_zz_1741[35:0]        ), //i
    .dout    (fixTo_780_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_781 (
    .din     (_zz_1742[35:0]        ), //i
    .dout    (fixTo_781_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_782 (
    .din     (_zz_1743[35:0]        ), //i
    .dout    (fixTo_782_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_783 (
    .din     (_zz_1744[35:0]        ), //i
    .dout    (fixTo_783_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_784 (
    .din     (_zz_1745[35:0]        ), //i
    .dout    (fixTo_784_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_785 (
    .din     (_zz_1746[35:0]        ), //i
    .dout    (fixTo_785_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_786 (
    .din     (_zz_1747[35:0]        ), //i
    .dout    (fixTo_786_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_787 (
    .din     (_zz_1748[35:0]        ), //i
    .dout    (fixTo_787_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_788 (
    .din     (_zz_1749[35:0]        ), //i
    .dout    (fixTo_788_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_789 (
    .din     (_zz_1750[35:0]        ), //i
    .dout    (fixTo_789_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_790 (
    .din     (_zz_1751[35:0]        ), //i
    .dout    (fixTo_790_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_791 (
    .din     (_zz_1752[35:0]        ), //i
    .dout    (fixTo_791_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_792 (
    .din     (_zz_1753[35:0]        ), //i
    .dout    (fixTo_792_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_793 (
    .din     (_zz_1754[35:0]        ), //i
    .dout    (fixTo_793_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_794 (
    .din     (_zz_1755[35:0]        ), //i
    .dout    (fixTo_794_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_795 (
    .din     (_zz_1756[35:0]        ), //i
    .dout    (fixTo_795_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_796 (
    .din     (_zz_1757[35:0]        ), //i
    .dout    (fixTo_796_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_797 (
    .din     (_zz_1758[35:0]        ), //i
    .dout    (fixTo_797_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_798 (
    .din     (_zz_1759[35:0]        ), //i
    .dout    (fixTo_798_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_799 (
    .din     (_zz_1760[35:0]        ), //i
    .dout    (fixTo_799_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_800 (
    .din     (_zz_1761[35:0]        ), //i
    .dout    (fixTo_800_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_801 (
    .din     (_zz_1762[35:0]        ), //i
    .dout    (fixTo_801_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_802 (
    .din     (_zz_1763[35:0]        ), //i
    .dout    (fixTo_802_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_803 (
    .din     (_zz_1764[35:0]        ), //i
    .dout    (fixTo_803_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_804 (
    .din     (_zz_1765[35:0]        ), //i
    .dout    (fixTo_804_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_805 (
    .din     (_zz_1766[35:0]        ), //i
    .dout    (fixTo_805_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_806 (
    .din     (_zz_1767[35:0]        ), //i
    .dout    (fixTo_806_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_807 (
    .din     (_zz_1768[35:0]        ), //i
    .dout    (fixTo_807_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_808 (
    .din     (_zz_1769[35:0]        ), //i
    .dout    (fixTo_808_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_809 (
    .din     (_zz_1770[35:0]        ), //i
    .dout    (fixTo_809_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_810 (
    .din     (_zz_1771[35:0]        ), //i
    .dout    (fixTo_810_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_811 (
    .din     (_zz_1772[35:0]        ), //i
    .dout    (fixTo_811_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_812 (
    .din     (_zz_1773[35:0]        ), //i
    .dout    (fixTo_812_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_813 (
    .din     (_zz_1774[35:0]        ), //i
    .dout    (fixTo_813_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_814 (
    .din     (_zz_1775[35:0]        ), //i
    .dout    (fixTo_814_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_815 (
    .din     (_zz_1776[35:0]        ), //i
    .dout    (fixTo_815_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_816 (
    .din     (_zz_1777[35:0]        ), //i
    .dout    (fixTo_816_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_817 (
    .din     (_zz_1778[35:0]        ), //i
    .dout    (fixTo_817_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_818 (
    .din     (_zz_1779[35:0]        ), //i
    .dout    (fixTo_818_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_819 (
    .din     (_zz_1780[35:0]        ), //i
    .dout    (fixTo_819_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_820 (
    .din     (_zz_1781[35:0]        ), //i
    .dout    (fixTo_820_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_821 (
    .din     (_zz_1782[35:0]        ), //i
    .dout    (fixTo_821_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_822 (
    .din     (_zz_1783[35:0]        ), //i
    .dout    (fixTo_822_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_823 (
    .din     (_zz_1784[35:0]        ), //i
    .dout    (fixTo_823_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_824 (
    .din     (_zz_1785[35:0]        ), //i
    .dout    (fixTo_824_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_825 (
    .din     (_zz_1786[35:0]        ), //i
    .dout    (fixTo_825_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_826 (
    .din     (_zz_1787[35:0]        ), //i
    .dout    (fixTo_826_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_827 (
    .din     (_zz_1788[35:0]        ), //i
    .dout    (fixTo_827_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_828 (
    .din     (_zz_1789[35:0]        ), //i
    .dout    (fixTo_828_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_829 (
    .din     (_zz_1790[35:0]        ), //i
    .dout    (fixTo_829_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_830 (
    .din     (_zz_1791[35:0]        ), //i
    .dout    (fixTo_830_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_831 (
    .din     (_zz_1792[35:0]        ), //i
    .dout    (fixTo_831_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_832 (
    .din     (_zz_1793[35:0]        ), //i
    .dout    (fixTo_832_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_833 (
    .din     (_zz_1794[35:0]        ), //i
    .dout    (fixTo_833_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_834 (
    .din     (_zz_1795[35:0]        ), //i
    .dout    (fixTo_834_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_835 (
    .din     (_zz_1796[35:0]        ), //i
    .dout    (fixTo_835_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_836 (
    .din     (_zz_1797[35:0]        ), //i
    .dout    (fixTo_836_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_837 (
    .din     (_zz_1798[35:0]        ), //i
    .dout    (fixTo_837_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_838 (
    .din     (_zz_1799[35:0]        ), //i
    .dout    (fixTo_838_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_839 (
    .din     (_zz_1800[35:0]        ), //i
    .dout    (fixTo_839_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_840 (
    .din     (_zz_1801[35:0]        ), //i
    .dout    (fixTo_840_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_841 (
    .din     (_zz_1802[35:0]        ), //i
    .dout    (fixTo_841_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_842 (
    .din     (_zz_1803[35:0]        ), //i
    .dout    (fixTo_842_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_843 (
    .din     (_zz_1804[35:0]        ), //i
    .dout    (fixTo_843_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_844 (
    .din     (_zz_1805[35:0]        ), //i
    .dout    (fixTo_844_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_845 (
    .din     (_zz_1806[35:0]        ), //i
    .dout    (fixTo_845_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_846 (
    .din     (_zz_1807[35:0]        ), //i
    .dout    (fixTo_846_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_847 (
    .din     (_zz_1808[35:0]        ), //i
    .dout    (fixTo_847_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_848 (
    .din     (_zz_1809[35:0]        ), //i
    .dout    (fixTo_848_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_849 (
    .din     (_zz_1810[35:0]        ), //i
    .dout    (fixTo_849_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_850 (
    .din     (_zz_1811[35:0]        ), //i
    .dout    (fixTo_850_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_851 (
    .din     (_zz_1812[35:0]        ), //i
    .dout    (fixTo_851_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_852 (
    .din     (_zz_1813[35:0]        ), //i
    .dout    (fixTo_852_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_853 (
    .din     (_zz_1814[35:0]        ), //i
    .dout    (fixTo_853_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_854 (
    .din     (_zz_1815[35:0]        ), //i
    .dout    (fixTo_854_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_855 (
    .din     (_zz_1816[35:0]        ), //i
    .dout    (fixTo_855_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_856 (
    .din     (_zz_1817[35:0]        ), //i
    .dout    (fixTo_856_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_857 (
    .din     (_zz_1818[35:0]        ), //i
    .dout    (fixTo_857_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_858 (
    .din     (_zz_1819[35:0]        ), //i
    .dout    (fixTo_858_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_859 (
    .din     (_zz_1820[35:0]        ), //i
    .dout    (fixTo_859_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_860 (
    .din     (_zz_1821[35:0]        ), //i
    .dout    (fixTo_860_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_861 (
    .din     (_zz_1822[35:0]        ), //i
    .dout    (fixTo_861_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_862 (
    .din     (_zz_1823[35:0]        ), //i
    .dout    (fixTo_862_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_863 (
    .din     (_zz_1824[35:0]        ), //i
    .dout    (fixTo_863_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_864 (
    .din     (_zz_1825[35:0]        ), //i
    .dout    (fixTo_864_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_865 (
    .din     (_zz_1826[35:0]        ), //i
    .dout    (fixTo_865_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_866 (
    .din     (_zz_1827[35:0]        ), //i
    .dout    (fixTo_866_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_867 (
    .din     (_zz_1828[35:0]        ), //i
    .dout    (fixTo_867_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_868 (
    .din     (_zz_1829[35:0]        ), //i
    .dout    (fixTo_868_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_869 (
    .din     (_zz_1830[35:0]        ), //i
    .dout    (fixTo_869_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_870 (
    .din     (_zz_1831[35:0]        ), //i
    .dout    (fixTo_870_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_871 (
    .din     (_zz_1832[35:0]        ), //i
    .dout    (fixTo_871_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_872 (
    .din     (_zz_1833[35:0]        ), //i
    .dout    (fixTo_872_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_873 (
    .din     (_zz_1834[35:0]        ), //i
    .dout    (fixTo_873_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_874 (
    .din     (_zz_1835[35:0]        ), //i
    .dout    (fixTo_874_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_875 (
    .din     (_zz_1836[35:0]        ), //i
    .dout    (fixTo_875_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_876 (
    .din     (_zz_1837[35:0]        ), //i
    .dout    (fixTo_876_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_877 (
    .din     (_zz_1838[35:0]        ), //i
    .dout    (fixTo_877_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_878 (
    .din     (_zz_1839[35:0]        ), //i
    .dout    (fixTo_878_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_879 (
    .din     (_zz_1840[35:0]        ), //i
    .dout    (fixTo_879_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_880 (
    .din     (_zz_1841[35:0]        ), //i
    .dout    (fixTo_880_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_881 (
    .din     (_zz_1842[35:0]        ), //i
    .dout    (fixTo_881_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_882 (
    .din     (_zz_1843[35:0]        ), //i
    .dout    (fixTo_882_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_883 (
    .din     (_zz_1844[35:0]        ), //i
    .dout    (fixTo_883_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_884 (
    .din     (_zz_1845[35:0]        ), //i
    .dout    (fixTo_884_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_885 (
    .din     (_zz_1846[35:0]        ), //i
    .dout    (fixTo_885_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_886 (
    .din     (_zz_1847[35:0]        ), //i
    .dout    (fixTo_886_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_887 (
    .din     (_zz_1848[35:0]        ), //i
    .dout    (fixTo_887_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_888 (
    .din     (_zz_1849[35:0]        ), //i
    .dout    (fixTo_888_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_889 (
    .din     (_zz_1850[35:0]        ), //i
    .dout    (fixTo_889_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_890 (
    .din     (_zz_1851[35:0]        ), //i
    .dout    (fixTo_890_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_891 (
    .din     (_zz_1852[35:0]        ), //i
    .dout    (fixTo_891_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_892 (
    .din     (_zz_1853[35:0]        ), //i
    .dout    (fixTo_892_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_893 (
    .din     (_zz_1854[35:0]        ), //i
    .dout    (fixTo_893_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_894 (
    .din     (_zz_1855[35:0]        ), //i
    .dout    (fixTo_894_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_895 (
    .din     (_zz_1856[35:0]        ), //i
    .dout    (fixTo_895_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_896 (
    .din     (_zz_1857[35:0]        ), //i
    .dout    (fixTo_896_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_897 (
    .din     (_zz_1858[35:0]        ), //i
    .dout    (fixTo_897_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_898 (
    .din     (_zz_1859[35:0]        ), //i
    .dout    (fixTo_898_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_899 (
    .din     (_zz_1860[35:0]        ), //i
    .dout    (fixTo_899_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_900 (
    .din     (_zz_1861[35:0]        ), //i
    .dout    (fixTo_900_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_901 (
    .din     (_zz_1862[35:0]        ), //i
    .dout    (fixTo_901_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_902 (
    .din     (_zz_1863[35:0]        ), //i
    .dout    (fixTo_902_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_903 (
    .din     (_zz_1864[35:0]        ), //i
    .dout    (fixTo_903_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_904 (
    .din     (_zz_1865[35:0]        ), //i
    .dout    (fixTo_904_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_905 (
    .din     (_zz_1866[35:0]        ), //i
    .dout    (fixTo_905_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_906 (
    .din     (_zz_1867[35:0]        ), //i
    .dout    (fixTo_906_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_907 (
    .din     (_zz_1868[35:0]        ), //i
    .dout    (fixTo_907_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_908 (
    .din     (_zz_1869[35:0]        ), //i
    .dout    (fixTo_908_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_909 (
    .din     (_zz_1870[35:0]        ), //i
    .dout    (fixTo_909_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_910 (
    .din     (_zz_1871[35:0]        ), //i
    .dout    (fixTo_910_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_911 (
    .din     (_zz_1872[35:0]        ), //i
    .dout    (fixTo_911_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_912 (
    .din     (_zz_1873[35:0]        ), //i
    .dout    (fixTo_912_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_913 (
    .din     (_zz_1874[35:0]        ), //i
    .dout    (fixTo_913_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_914 (
    .din     (_zz_1875[35:0]        ), //i
    .dout    (fixTo_914_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_915 (
    .din     (_zz_1876[35:0]        ), //i
    .dout    (fixTo_915_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_916 (
    .din     (_zz_1877[35:0]        ), //i
    .dout    (fixTo_916_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_917 (
    .din     (_zz_1878[35:0]        ), //i
    .dout    (fixTo_917_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_918 (
    .din     (_zz_1879[35:0]        ), //i
    .dout    (fixTo_918_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_919 (
    .din     (_zz_1880[35:0]        ), //i
    .dout    (fixTo_919_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_920 (
    .din     (_zz_1881[35:0]        ), //i
    .dout    (fixTo_920_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_921 (
    .din     (_zz_1882[35:0]        ), //i
    .dout    (fixTo_921_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_922 (
    .din     (_zz_1883[35:0]        ), //i
    .dout    (fixTo_922_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_923 (
    .din     (_zz_1884[35:0]        ), //i
    .dout    (fixTo_923_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_924 (
    .din     (_zz_1885[35:0]        ), //i
    .dout    (fixTo_924_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_925 (
    .din     (_zz_1886[35:0]        ), //i
    .dout    (fixTo_925_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_926 (
    .din     (_zz_1887[35:0]        ), //i
    .dout    (fixTo_926_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_927 (
    .din     (_zz_1888[35:0]        ), //i
    .dout    (fixTo_927_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_928 (
    .din     (_zz_1889[35:0]        ), //i
    .dout    (fixTo_928_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_929 (
    .din     (_zz_1890[35:0]        ), //i
    .dout    (fixTo_929_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_930 (
    .din     (_zz_1891[35:0]        ), //i
    .dout    (fixTo_930_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_931 (
    .din     (_zz_1892[35:0]        ), //i
    .dout    (fixTo_931_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_932 (
    .din     (_zz_1893[35:0]        ), //i
    .dout    (fixTo_932_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_933 (
    .din     (_zz_1894[35:0]        ), //i
    .dout    (fixTo_933_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_934 (
    .din     (_zz_1895[35:0]        ), //i
    .dout    (fixTo_934_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_935 (
    .din     (_zz_1896[35:0]        ), //i
    .dout    (fixTo_935_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_936 (
    .din     (_zz_1897[35:0]        ), //i
    .dout    (fixTo_936_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_937 (
    .din     (_zz_1898[35:0]        ), //i
    .dout    (fixTo_937_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_938 (
    .din     (_zz_1899[35:0]        ), //i
    .dout    (fixTo_938_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_939 (
    .din     (_zz_1900[35:0]        ), //i
    .dout    (fixTo_939_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_940 (
    .din     (_zz_1901[35:0]        ), //i
    .dout    (fixTo_940_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_941 (
    .din     (_zz_1902[35:0]        ), //i
    .dout    (fixTo_941_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_942 (
    .din     (_zz_1903[35:0]        ), //i
    .dout    (fixTo_942_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_943 (
    .din     (_zz_1904[35:0]        ), //i
    .dout    (fixTo_943_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_944 (
    .din     (_zz_1905[35:0]        ), //i
    .dout    (fixTo_944_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_945 (
    .din     (_zz_1906[35:0]        ), //i
    .dout    (fixTo_945_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_946 (
    .din     (_zz_1907[35:0]        ), //i
    .dout    (fixTo_946_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_947 (
    .din     (_zz_1908[35:0]        ), //i
    .dout    (fixTo_947_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_948 (
    .din     (_zz_1909[35:0]        ), //i
    .dout    (fixTo_948_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_949 (
    .din     (_zz_1910[35:0]        ), //i
    .dout    (fixTo_949_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_950 (
    .din     (_zz_1911[35:0]        ), //i
    .dout    (fixTo_950_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_951 (
    .din     (_zz_1912[35:0]        ), //i
    .dout    (fixTo_951_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_952 (
    .din     (_zz_1913[35:0]        ), //i
    .dout    (fixTo_952_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_953 (
    .din     (_zz_1914[35:0]        ), //i
    .dout    (fixTo_953_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_954 (
    .din     (_zz_1915[35:0]        ), //i
    .dout    (fixTo_954_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_955 (
    .din     (_zz_1916[35:0]        ), //i
    .dout    (fixTo_955_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_956 (
    .din     (_zz_1917[35:0]        ), //i
    .dout    (fixTo_956_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_957 (
    .din     (_zz_1918[35:0]        ), //i
    .dout    (fixTo_957_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_958 (
    .din     (_zz_1919[35:0]        ), //i
    .dout    (fixTo_958_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_959 (
    .din     (_zz_1920[35:0]        ), //i
    .dout    (fixTo_959_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_960 (
    .din     (_zz_1921[35:0]        ), //i
    .dout    (fixTo_960_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_961 (
    .din     (_zz_1922[35:0]        ), //i
    .dout    (fixTo_961_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_962 (
    .din     (_zz_1923[35:0]        ), //i
    .dout    (fixTo_962_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_963 (
    .din     (_zz_1924[35:0]        ), //i
    .dout    (fixTo_963_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_964 (
    .din     (_zz_1925[35:0]        ), //i
    .dout    (fixTo_964_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_965 (
    .din     (_zz_1926[35:0]        ), //i
    .dout    (fixTo_965_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_966 (
    .din     (_zz_1927[35:0]        ), //i
    .dout    (fixTo_966_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_967 (
    .din     (_zz_1928[35:0]        ), //i
    .dout    (fixTo_967_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_968 (
    .din     (_zz_1929[35:0]        ), //i
    .dout    (fixTo_968_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_969 (
    .din     (_zz_1930[35:0]        ), //i
    .dout    (fixTo_969_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_970 (
    .din     (_zz_1931[35:0]        ), //i
    .dout    (fixTo_970_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_971 (
    .din     (_zz_1932[35:0]        ), //i
    .dout    (fixTo_971_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_972 (
    .din     (_zz_1933[35:0]        ), //i
    .dout    (fixTo_972_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_973 (
    .din     (_zz_1934[35:0]        ), //i
    .dout    (fixTo_973_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_974 (
    .din     (_zz_1935[35:0]        ), //i
    .dout    (fixTo_974_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_975 (
    .din     (_zz_1936[35:0]        ), //i
    .dout    (fixTo_975_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_976 (
    .din     (_zz_1937[35:0]        ), //i
    .dout    (fixTo_976_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_977 (
    .din     (_zz_1938[35:0]        ), //i
    .dout    (fixTo_977_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_978 (
    .din     (_zz_1939[35:0]        ), //i
    .dout    (fixTo_978_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_979 (
    .din     (_zz_1940[35:0]        ), //i
    .dout    (fixTo_979_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_980 (
    .din     (_zz_1941[35:0]        ), //i
    .dout    (fixTo_980_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_981 (
    .din     (_zz_1942[35:0]        ), //i
    .dout    (fixTo_981_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_982 (
    .din     (_zz_1943[35:0]        ), //i
    .dout    (fixTo_982_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_983 (
    .din     (_zz_1944[35:0]        ), //i
    .dout    (fixTo_983_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_984 (
    .din     (_zz_1945[35:0]        ), //i
    .dout    (fixTo_984_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_985 (
    .din     (_zz_1946[35:0]        ), //i
    .dout    (fixTo_985_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_986 (
    .din     (_zz_1947[35:0]        ), //i
    .dout    (fixTo_986_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_987 (
    .din     (_zz_1948[35:0]        ), //i
    .dout    (fixTo_987_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_988 (
    .din     (_zz_1949[35:0]        ), //i
    .dout    (fixTo_988_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_989 (
    .din     (_zz_1950[35:0]        ), //i
    .dout    (fixTo_989_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_990 (
    .din     (_zz_1951[35:0]        ), //i
    .dout    (fixTo_990_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_991 (
    .din     (_zz_1952[35:0]        ), //i
    .dout    (fixTo_991_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_992 (
    .din     (_zz_1953[35:0]        ), //i
    .dout    (fixTo_992_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_993 (
    .din     (_zz_1954[35:0]        ), //i
    .dout    (fixTo_993_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_994 (
    .din     (_zz_1955[35:0]        ), //i
    .dout    (fixTo_994_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_995 (
    .din     (_zz_1956[35:0]        ), //i
    .dout    (fixTo_995_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_996 (
    .din     (_zz_1957[35:0]        ), //i
    .dout    (fixTo_996_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_997 (
    .din     (_zz_1958[35:0]        ), //i
    .dout    (fixTo_997_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_998 (
    .din     (_zz_1959[35:0]        ), //i
    .dout    (fixTo_998_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_999 (
    .din     (_zz_1960[35:0]        ), //i
    .dout    (fixTo_999_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1000 (
    .din     (_zz_1961[35:0]         ), //i
    .dout    (fixTo_1000_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1001 (
    .din     (_zz_1962[35:0]         ), //i
    .dout    (fixTo_1001_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1002 (
    .din     (_zz_1963[35:0]         ), //i
    .dout    (fixTo_1002_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1003 (
    .din     (_zz_1964[35:0]         ), //i
    .dout    (fixTo_1003_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1004 (
    .din     (_zz_1965[35:0]         ), //i
    .dout    (fixTo_1004_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1005 (
    .din     (_zz_1966[35:0]         ), //i
    .dout    (fixTo_1005_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1006 (
    .din     (_zz_1967[35:0]         ), //i
    .dout    (fixTo_1006_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1007 (
    .din     (_zz_1968[35:0]         ), //i
    .dout    (fixTo_1007_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1008 (
    .din     (_zz_1969[35:0]         ), //i
    .dout    (fixTo_1008_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1009 (
    .din     (_zz_1970[35:0]         ), //i
    .dout    (fixTo_1009_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1010 (
    .din     (_zz_1971[35:0]         ), //i
    .dout    (fixTo_1010_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1011 (
    .din     (_zz_1972[35:0]         ), //i
    .dout    (fixTo_1011_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1012 (
    .din     (_zz_1973[35:0]         ), //i
    .dout    (fixTo_1012_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1013 (
    .din     (_zz_1974[35:0]         ), //i
    .dout    (fixTo_1013_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1014 (
    .din     (_zz_1975[35:0]         ), //i
    .dout    (fixTo_1014_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1015 (
    .din     (_zz_1976[35:0]         ), //i
    .dout    (fixTo_1015_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1016 (
    .din     (_zz_1977[35:0]         ), //i
    .dout    (fixTo_1016_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1017 (
    .din     (_zz_1978[35:0]         ), //i
    .dout    (fixTo_1017_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1018 (
    .din     (_zz_1979[35:0]         ), //i
    .dout    (fixTo_1018_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1019 (
    .din     (_zz_1980[35:0]         ), //i
    .dout    (fixTo_1019_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1020 (
    .din     (_zz_1981[35:0]         ), //i
    .dout    (fixTo_1020_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1021 (
    .din     (_zz_1982[35:0]         ), //i
    .dout    (fixTo_1021_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1022 (
    .din     (_zz_1983[35:0]         ), //i
    .dout    (fixTo_1022_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1023 (
    .din     (_zz_1984[35:0]         ), //i
    .dout    (fixTo_1023_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1024 (
    .din     (_zz_1985[35:0]         ), //i
    .dout    (fixTo_1024_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1025 (
    .din     (_zz_1986[35:0]         ), //i
    .dout    (fixTo_1025_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1026 (
    .din     (_zz_1987[35:0]         ), //i
    .dout    (fixTo_1026_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1027 (
    .din     (_zz_1988[35:0]         ), //i
    .dout    (fixTo_1027_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1028 (
    .din     (_zz_1989[35:0]         ), //i
    .dout    (fixTo_1028_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1029 (
    .din     (_zz_1990[35:0]         ), //i
    .dout    (fixTo_1029_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1030 (
    .din     (_zz_1991[35:0]         ), //i
    .dout    (fixTo_1030_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1031 (
    .din     (_zz_1992[35:0]         ), //i
    .dout    (fixTo_1031_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1032 (
    .din     (_zz_1993[35:0]         ), //i
    .dout    (fixTo_1032_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1033 (
    .din     (_zz_1994[35:0]         ), //i
    .dout    (fixTo_1033_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1034 (
    .din     (_zz_1995[35:0]         ), //i
    .dout    (fixTo_1034_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1035 (
    .din     (_zz_1996[35:0]         ), //i
    .dout    (fixTo_1035_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1036 (
    .din     (_zz_1997[35:0]         ), //i
    .dout    (fixTo_1036_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1037 (
    .din     (_zz_1998[35:0]         ), //i
    .dout    (fixTo_1037_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1038 (
    .din     (_zz_1999[35:0]         ), //i
    .dout    (fixTo_1038_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1039 (
    .din     (_zz_2000[35:0]         ), //i
    .dout    (fixTo_1039_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1040 (
    .din     (_zz_2001[35:0]         ), //i
    .dout    (fixTo_1040_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1041 (
    .din     (_zz_2002[35:0]         ), //i
    .dout    (fixTo_1041_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1042 (
    .din     (_zz_2003[35:0]         ), //i
    .dout    (fixTo_1042_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1043 (
    .din     (_zz_2004[35:0]         ), //i
    .dout    (fixTo_1043_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1044 (
    .din     (_zz_2005[35:0]         ), //i
    .dout    (fixTo_1044_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1045 (
    .din     (_zz_2006[35:0]         ), //i
    .dout    (fixTo_1045_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1046 (
    .din     (_zz_2007[35:0]         ), //i
    .dout    (fixTo_1046_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1047 (
    .din     (_zz_2008[35:0]         ), //i
    .dout    (fixTo_1047_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1048 (
    .din     (_zz_2009[35:0]         ), //i
    .dout    (fixTo_1048_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1049 (
    .din     (_zz_2010[35:0]         ), //i
    .dout    (fixTo_1049_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1050 (
    .din     (_zz_2011[35:0]         ), //i
    .dout    (fixTo_1050_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1051 (
    .din     (_zz_2012[35:0]         ), //i
    .dout    (fixTo_1051_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1052 (
    .din     (_zz_2013[35:0]         ), //i
    .dout    (fixTo_1052_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1053 (
    .din     (_zz_2014[35:0]         ), //i
    .dout    (fixTo_1053_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1054 (
    .din     (_zz_2015[35:0]         ), //i
    .dout    (fixTo_1054_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1055 (
    .din     (_zz_2016[35:0]         ), //i
    .dout    (fixTo_1055_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1056 (
    .din     (_zz_2017[35:0]         ), //i
    .dout    (fixTo_1056_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1057 (
    .din     (_zz_2018[35:0]         ), //i
    .dout    (fixTo_1057_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1058 (
    .din     (_zz_2019[35:0]         ), //i
    .dout    (fixTo_1058_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1059 (
    .din     (_zz_2020[35:0]         ), //i
    .dout    (fixTo_1059_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1060 (
    .din     (_zz_2021[35:0]         ), //i
    .dout    (fixTo_1060_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1061 (
    .din     (_zz_2022[35:0]         ), //i
    .dout    (fixTo_1061_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1062 (
    .din     (_zz_2023[35:0]         ), //i
    .dout    (fixTo_1062_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1063 (
    .din     (_zz_2024[35:0]         ), //i
    .dout    (fixTo_1063_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1064 (
    .din     (_zz_2025[35:0]         ), //i
    .dout    (fixTo_1064_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1065 (
    .din     (_zz_2026[35:0]         ), //i
    .dout    (fixTo_1065_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1066 (
    .din     (_zz_2027[35:0]         ), //i
    .dout    (fixTo_1066_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1067 (
    .din     (_zz_2028[35:0]         ), //i
    .dout    (fixTo_1067_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1068 (
    .din     (_zz_2029[35:0]         ), //i
    .dout    (fixTo_1068_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1069 (
    .din     (_zz_2030[35:0]         ), //i
    .dout    (fixTo_1069_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1070 (
    .din     (_zz_2031[35:0]         ), //i
    .dout    (fixTo_1070_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1071 (
    .din     (_zz_2032[35:0]         ), //i
    .dout    (fixTo_1071_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1072 (
    .din     (_zz_2033[35:0]         ), //i
    .dout    (fixTo_1072_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1073 (
    .din     (_zz_2034[35:0]         ), //i
    .dout    (fixTo_1073_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1074 (
    .din     (_zz_2035[35:0]         ), //i
    .dout    (fixTo_1074_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1075 (
    .din     (_zz_2036[35:0]         ), //i
    .dout    (fixTo_1075_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1076 (
    .din     (_zz_2037[35:0]         ), //i
    .dout    (fixTo_1076_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1077 (
    .din     (_zz_2038[35:0]         ), //i
    .dout    (fixTo_1077_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1078 (
    .din     (_zz_2039[35:0]         ), //i
    .dout    (fixTo_1078_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1079 (
    .din     (_zz_2040[35:0]         ), //i
    .dout    (fixTo_1079_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1080 (
    .din     (_zz_2041[35:0]         ), //i
    .dout    (fixTo_1080_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1081 (
    .din     (_zz_2042[35:0]         ), //i
    .dout    (fixTo_1081_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1082 (
    .din     (_zz_2043[35:0]         ), //i
    .dout    (fixTo_1082_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1083 (
    .din     (_zz_2044[35:0]         ), //i
    .dout    (fixTo_1083_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1084 (
    .din     (_zz_2045[35:0]         ), //i
    .dout    (fixTo_1084_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1085 (
    .din     (_zz_2046[35:0]         ), //i
    .dout    (fixTo_1085_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1086 (
    .din     (_zz_2047[35:0]         ), //i
    .dout    (fixTo_1086_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1087 (
    .din     (_zz_2048[35:0]         ), //i
    .dout    (fixTo_1087_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1088 (
    .din     (_zz_2049[35:0]         ), //i
    .dout    (fixTo_1088_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1089 (
    .din     (_zz_2050[35:0]         ), //i
    .dout    (fixTo_1089_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1090 (
    .din     (_zz_2051[35:0]         ), //i
    .dout    (fixTo_1090_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1091 (
    .din     (_zz_2052[35:0]         ), //i
    .dout    (fixTo_1091_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1092 (
    .din     (_zz_2053[35:0]         ), //i
    .dout    (fixTo_1092_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1093 (
    .din     (_zz_2054[35:0]         ), //i
    .dout    (fixTo_1093_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1094 (
    .din     (_zz_2055[35:0]         ), //i
    .dout    (fixTo_1094_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1095 (
    .din     (_zz_2056[35:0]         ), //i
    .dout    (fixTo_1095_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1096 (
    .din     (_zz_2057[35:0]         ), //i
    .dout    (fixTo_1096_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1097 (
    .din     (_zz_2058[35:0]         ), //i
    .dout    (fixTo_1097_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1098 (
    .din     (_zz_2059[35:0]         ), //i
    .dout    (fixTo_1098_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1099 (
    .din     (_zz_2060[35:0]         ), //i
    .dout    (fixTo_1099_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1100 (
    .din     (_zz_2061[35:0]         ), //i
    .dout    (fixTo_1100_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1101 (
    .din     (_zz_2062[35:0]         ), //i
    .dout    (fixTo_1101_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1102 (
    .din     (_zz_2063[35:0]         ), //i
    .dout    (fixTo_1102_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1103 (
    .din     (_zz_2064[35:0]         ), //i
    .dout    (fixTo_1103_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1104 (
    .din     (_zz_2065[35:0]         ), //i
    .dout    (fixTo_1104_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1105 (
    .din     (_zz_2066[35:0]         ), //i
    .dout    (fixTo_1105_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1106 (
    .din     (_zz_2067[35:0]         ), //i
    .dout    (fixTo_1106_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1107 (
    .din     (_zz_2068[35:0]         ), //i
    .dout    (fixTo_1107_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1108 (
    .din     (_zz_2069[35:0]         ), //i
    .dout    (fixTo_1108_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1109 (
    .din     (_zz_2070[35:0]         ), //i
    .dout    (fixTo_1109_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1110 (
    .din     (_zz_2071[35:0]         ), //i
    .dout    (fixTo_1110_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1111 (
    .din     (_zz_2072[35:0]         ), //i
    .dout    (fixTo_1111_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1112 (
    .din     (_zz_2073[35:0]         ), //i
    .dout    (fixTo_1112_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1113 (
    .din     (_zz_2074[35:0]         ), //i
    .dout    (fixTo_1113_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1114 (
    .din     (_zz_2075[35:0]         ), //i
    .dout    (fixTo_1114_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1115 (
    .din     (_zz_2076[35:0]         ), //i
    .dout    (fixTo_1115_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1116 (
    .din     (_zz_2077[35:0]         ), //i
    .dout    (fixTo_1116_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1117 (
    .din     (_zz_2078[35:0]         ), //i
    .dout    (fixTo_1117_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1118 (
    .din     (_zz_2079[35:0]         ), //i
    .dout    (fixTo_1118_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1119 (
    .din     (_zz_2080[35:0]         ), //i
    .dout    (fixTo_1119_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1120 (
    .din     (_zz_2081[35:0]         ), //i
    .dout    (fixTo_1120_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1121 (
    .din     (_zz_2082[35:0]         ), //i
    .dout    (fixTo_1121_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1122 (
    .din     (_zz_2083[35:0]         ), //i
    .dout    (fixTo_1122_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1123 (
    .din     (_zz_2084[35:0]         ), //i
    .dout    (fixTo_1123_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1124 (
    .din     (_zz_2085[35:0]         ), //i
    .dout    (fixTo_1124_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1125 (
    .din     (_zz_2086[35:0]         ), //i
    .dout    (fixTo_1125_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1126 (
    .din     (_zz_2087[35:0]         ), //i
    .dout    (fixTo_1126_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1127 (
    .din     (_zz_2088[35:0]         ), //i
    .dout    (fixTo_1127_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1128 (
    .din     (_zz_2089[35:0]         ), //i
    .dout    (fixTo_1128_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1129 (
    .din     (_zz_2090[35:0]         ), //i
    .dout    (fixTo_1129_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1130 (
    .din     (_zz_2091[35:0]         ), //i
    .dout    (fixTo_1130_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1131 (
    .din     (_zz_2092[35:0]         ), //i
    .dout    (fixTo_1131_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1132 (
    .din     (_zz_2093[35:0]         ), //i
    .dout    (fixTo_1132_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1133 (
    .din     (_zz_2094[35:0]         ), //i
    .dout    (fixTo_1133_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1134 (
    .din     (_zz_2095[35:0]         ), //i
    .dout    (fixTo_1134_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1135 (
    .din     (_zz_2096[35:0]         ), //i
    .dout    (fixTo_1135_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1136 (
    .din     (_zz_2097[35:0]         ), //i
    .dout    (fixTo_1136_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1137 (
    .din     (_zz_2098[35:0]         ), //i
    .dout    (fixTo_1137_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1138 (
    .din     (_zz_2099[35:0]         ), //i
    .dout    (fixTo_1138_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1139 (
    .din     (_zz_2100[35:0]         ), //i
    .dout    (fixTo_1139_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1140 (
    .din     (_zz_2101[35:0]         ), //i
    .dout    (fixTo_1140_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1141 (
    .din     (_zz_2102[35:0]         ), //i
    .dout    (fixTo_1141_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1142 (
    .din     (_zz_2103[35:0]         ), //i
    .dout    (fixTo_1142_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1143 (
    .din     (_zz_2104[35:0]         ), //i
    .dout    (fixTo_1143_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1144 (
    .din     (_zz_2105[35:0]         ), //i
    .dout    (fixTo_1144_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1145 (
    .din     (_zz_2106[35:0]         ), //i
    .dout    (fixTo_1145_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1146 (
    .din     (_zz_2107[35:0]         ), //i
    .dout    (fixTo_1146_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1147 (
    .din     (_zz_2108[35:0]         ), //i
    .dout    (fixTo_1147_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1148 (
    .din     (_zz_2109[35:0]         ), //i
    .dout    (fixTo_1148_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1149 (
    .din     (_zz_2110[35:0]         ), //i
    .dout    (fixTo_1149_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1150 (
    .din     (_zz_2111[35:0]         ), //i
    .dout    (fixTo_1150_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1151 (
    .din     (_zz_2112[35:0]         ), //i
    .dout    (fixTo_1151_dout[17:0]  )  //o
  );
  assign twiddle_factor_table_0_real = 18'h00200;
  assign twiddle_factor_table_0_imag = 18'h0;
  assign twiddle_factor_table_1_real = 18'h00200;
  assign twiddle_factor_table_1_imag = 18'h0;
  assign twiddle_factor_table_2_real = 18'h0;
  assign twiddle_factor_table_2_imag = 18'h3fe00;
  assign twiddle_factor_table_3_real = 18'h00200;
  assign twiddle_factor_table_3_imag = 18'h0;
  assign twiddle_factor_table_4_real = 18'h0016a;
  assign twiddle_factor_table_4_imag = 18'h3fe96;
  assign twiddle_factor_table_5_real = 18'h0;
  assign twiddle_factor_table_5_imag = 18'h3fe00;
  assign twiddle_factor_table_6_real = 18'h3fe96;
  assign twiddle_factor_table_6_imag = 18'h3fe96;
  assign twiddle_factor_table_7_real = 18'h00200;
  assign twiddle_factor_table_7_imag = 18'h0;
  assign twiddle_factor_table_8_real = 18'h001d9;
  assign twiddle_factor_table_8_imag = 18'h3ff3d;
  assign twiddle_factor_table_9_real = 18'h0016a;
  assign twiddle_factor_table_9_imag = 18'h3fe96;
  assign twiddle_factor_table_10_real = 18'h000c3;
  assign twiddle_factor_table_10_imag = 18'h3fe27;
  assign twiddle_factor_table_11_real = 18'h0;
  assign twiddle_factor_table_11_imag = 18'h3fe00;
  assign twiddle_factor_table_12_real = 18'h3ff3d;
  assign twiddle_factor_table_12_imag = 18'h3fe27;
  assign twiddle_factor_table_13_real = 18'h3fe96;
  assign twiddle_factor_table_13_imag = 18'h3fe96;
  assign twiddle_factor_table_14_real = 18'h3fe27;
  assign twiddle_factor_table_14_imag = 18'h3ff3d;
  assign twiddle_factor_table_15_real = 18'h00200;
  assign twiddle_factor_table_15_imag = 18'h0;
  assign twiddle_factor_table_16_real = 18'h001f6;
  assign twiddle_factor_table_16_imag = 18'h3ff9d;
  assign twiddle_factor_table_17_real = 18'h001d9;
  assign twiddle_factor_table_17_imag = 18'h3ff3d;
  assign twiddle_factor_table_18_real = 18'h001a9;
  assign twiddle_factor_table_18_imag = 18'h3fee4;
  assign twiddle_factor_table_19_real = 18'h0016a;
  assign twiddle_factor_table_19_imag = 18'h3fe96;
  assign twiddle_factor_table_20_real = 18'h0011c;
  assign twiddle_factor_table_20_imag = 18'h3fe57;
  assign twiddle_factor_table_21_real = 18'h000c3;
  assign twiddle_factor_table_21_imag = 18'h3fe27;
  assign twiddle_factor_table_22_real = 18'h00063;
  assign twiddle_factor_table_22_imag = 18'h3fe0a;
  assign twiddle_factor_table_23_real = 18'h0;
  assign twiddle_factor_table_23_imag = 18'h3fe00;
  assign twiddle_factor_table_24_real = 18'h3ff9d;
  assign twiddle_factor_table_24_imag = 18'h3fe0a;
  assign twiddle_factor_table_25_real = 18'h3ff3d;
  assign twiddle_factor_table_25_imag = 18'h3fe27;
  assign twiddle_factor_table_26_real = 18'h3fee4;
  assign twiddle_factor_table_26_imag = 18'h3fe57;
  assign twiddle_factor_table_27_real = 18'h3fe96;
  assign twiddle_factor_table_27_imag = 18'h3fe96;
  assign twiddle_factor_table_28_real = 18'h3fe57;
  assign twiddle_factor_table_28_imag = 18'h3fee4;
  assign twiddle_factor_table_29_real = 18'h3fe27;
  assign twiddle_factor_table_29_imag = 18'h3ff3d;
  assign twiddle_factor_table_30_real = 18'h3fe0a;
  assign twiddle_factor_table_30_imag = 18'h3ff9d;
  assign twiddle_factor_table_31_real = 18'h00200;
  assign twiddle_factor_table_31_imag = 18'h0;
  assign twiddle_factor_table_32_real = 18'h001fd;
  assign twiddle_factor_table_32_imag = 18'h3ffce;
  assign twiddle_factor_table_33_real = 18'h001f6;
  assign twiddle_factor_table_33_imag = 18'h3ff9d;
  assign twiddle_factor_table_34_real = 18'h001e9;
  assign twiddle_factor_table_34_imag = 18'h3ff6c;
  assign twiddle_factor_table_35_real = 18'h001d9;
  assign twiddle_factor_table_35_imag = 18'h3ff3d;
  assign twiddle_factor_table_36_real = 18'h001c3;
  assign twiddle_factor_table_36_imag = 18'h3ff0f;
  assign twiddle_factor_table_37_real = 18'h001a9;
  assign twiddle_factor_table_37_imag = 18'h3fee4;
  assign twiddle_factor_table_38_real = 18'h0018b;
  assign twiddle_factor_table_38_imag = 18'h3febc;
  assign twiddle_factor_table_39_real = 18'h0016a;
  assign twiddle_factor_table_39_imag = 18'h3fe96;
  assign twiddle_factor_table_40_real = 18'h00144;
  assign twiddle_factor_table_40_imag = 18'h3fe75;
  assign twiddle_factor_table_41_real = 18'h0011c;
  assign twiddle_factor_table_41_imag = 18'h3fe57;
  assign twiddle_factor_table_42_real = 18'h000f1;
  assign twiddle_factor_table_42_imag = 18'h3fe3d;
  assign twiddle_factor_table_43_real = 18'h000c3;
  assign twiddle_factor_table_43_imag = 18'h3fe27;
  assign twiddle_factor_table_44_real = 18'h00094;
  assign twiddle_factor_table_44_imag = 18'h3fe17;
  assign twiddle_factor_table_45_real = 18'h00063;
  assign twiddle_factor_table_45_imag = 18'h3fe0a;
  assign twiddle_factor_table_46_real = 18'h00032;
  assign twiddle_factor_table_46_imag = 18'h3fe03;
  assign twiddle_factor_table_47_real = 18'h0;
  assign twiddle_factor_table_47_imag = 18'h3fe00;
  assign twiddle_factor_table_48_real = 18'h3ffce;
  assign twiddle_factor_table_48_imag = 18'h3fe03;
  assign twiddle_factor_table_49_real = 18'h3ff9d;
  assign twiddle_factor_table_49_imag = 18'h3fe0a;
  assign twiddle_factor_table_50_real = 18'h3ff6c;
  assign twiddle_factor_table_50_imag = 18'h3fe17;
  assign twiddle_factor_table_51_real = 18'h3ff3d;
  assign twiddle_factor_table_51_imag = 18'h3fe27;
  assign twiddle_factor_table_52_real = 18'h3ff0f;
  assign twiddle_factor_table_52_imag = 18'h3fe3d;
  assign twiddle_factor_table_53_real = 18'h3fee4;
  assign twiddle_factor_table_53_imag = 18'h3fe57;
  assign twiddle_factor_table_54_real = 18'h3febc;
  assign twiddle_factor_table_54_imag = 18'h3fe75;
  assign twiddle_factor_table_55_real = 18'h3fe96;
  assign twiddle_factor_table_55_imag = 18'h3fe96;
  assign twiddle_factor_table_56_real = 18'h3fe75;
  assign twiddle_factor_table_56_imag = 18'h3febc;
  assign twiddle_factor_table_57_real = 18'h3fe57;
  assign twiddle_factor_table_57_imag = 18'h3fee4;
  assign twiddle_factor_table_58_real = 18'h3fe3d;
  assign twiddle_factor_table_58_imag = 18'h3ff0f;
  assign twiddle_factor_table_59_real = 18'h3fe27;
  assign twiddle_factor_table_59_imag = 18'h3ff3d;
  assign twiddle_factor_table_60_real = 18'h3fe17;
  assign twiddle_factor_table_60_imag = 18'h3ff6c;
  assign twiddle_factor_table_61_real = 18'h3fe0a;
  assign twiddle_factor_table_61_imag = 18'h3ff9d;
  assign twiddle_factor_table_62_real = 18'h3fe03;
  assign twiddle_factor_table_62_imag = 18'h3ffce;
  assign data_reorder_0_real = data_in_0_real;
  assign data_reorder_0_imag = data_in_0_imag;
  assign data_reorder_32_real = data_in_1_real;
  assign data_reorder_32_imag = data_in_1_imag;
  assign data_reorder_16_real = data_in_2_real;
  assign data_reorder_16_imag = data_in_2_imag;
  assign data_reorder_48_real = data_in_3_real;
  assign data_reorder_48_imag = data_in_3_imag;
  assign data_reorder_8_real = data_in_4_real;
  assign data_reorder_8_imag = data_in_4_imag;
  assign data_reorder_40_real = data_in_5_real;
  assign data_reorder_40_imag = data_in_5_imag;
  assign data_reorder_24_real = data_in_6_real;
  assign data_reorder_24_imag = data_in_6_imag;
  assign data_reorder_56_real = data_in_7_real;
  assign data_reorder_56_imag = data_in_7_imag;
  assign data_reorder_4_real = data_in_8_real;
  assign data_reorder_4_imag = data_in_8_imag;
  assign data_reorder_36_real = data_in_9_real;
  assign data_reorder_36_imag = data_in_9_imag;
  assign data_reorder_20_real = data_in_10_real;
  assign data_reorder_20_imag = data_in_10_imag;
  assign data_reorder_52_real = data_in_11_real;
  assign data_reorder_52_imag = data_in_11_imag;
  assign data_reorder_12_real = data_in_12_real;
  assign data_reorder_12_imag = data_in_12_imag;
  assign data_reorder_44_real = data_in_13_real;
  assign data_reorder_44_imag = data_in_13_imag;
  assign data_reorder_28_real = data_in_14_real;
  assign data_reorder_28_imag = data_in_14_imag;
  assign data_reorder_60_real = data_in_15_real;
  assign data_reorder_60_imag = data_in_15_imag;
  assign data_reorder_2_real = data_in_16_real;
  assign data_reorder_2_imag = data_in_16_imag;
  assign data_reorder_34_real = data_in_17_real;
  assign data_reorder_34_imag = data_in_17_imag;
  assign data_reorder_18_real = data_in_18_real;
  assign data_reorder_18_imag = data_in_18_imag;
  assign data_reorder_50_real = data_in_19_real;
  assign data_reorder_50_imag = data_in_19_imag;
  assign data_reorder_10_real = data_in_20_real;
  assign data_reorder_10_imag = data_in_20_imag;
  assign data_reorder_42_real = data_in_21_real;
  assign data_reorder_42_imag = data_in_21_imag;
  assign data_reorder_26_real = data_in_22_real;
  assign data_reorder_26_imag = data_in_22_imag;
  assign data_reorder_58_real = data_in_23_real;
  assign data_reorder_58_imag = data_in_23_imag;
  assign data_reorder_6_real = data_in_24_real;
  assign data_reorder_6_imag = data_in_24_imag;
  assign data_reorder_38_real = data_in_25_real;
  assign data_reorder_38_imag = data_in_25_imag;
  assign data_reorder_22_real = data_in_26_real;
  assign data_reorder_22_imag = data_in_26_imag;
  assign data_reorder_54_real = data_in_27_real;
  assign data_reorder_54_imag = data_in_27_imag;
  assign data_reorder_14_real = data_in_28_real;
  assign data_reorder_14_imag = data_in_28_imag;
  assign data_reorder_46_real = data_in_29_real;
  assign data_reorder_46_imag = data_in_29_imag;
  assign data_reorder_30_real = data_in_30_real;
  assign data_reorder_30_imag = data_in_30_imag;
  assign data_reorder_62_real = data_in_31_real;
  assign data_reorder_62_imag = data_in_31_imag;
  assign data_reorder_1_real = data_in_32_real;
  assign data_reorder_1_imag = data_in_32_imag;
  assign data_reorder_33_real = data_in_33_real;
  assign data_reorder_33_imag = data_in_33_imag;
  assign data_reorder_17_real = data_in_34_real;
  assign data_reorder_17_imag = data_in_34_imag;
  assign data_reorder_49_real = data_in_35_real;
  assign data_reorder_49_imag = data_in_35_imag;
  assign data_reorder_9_real = data_in_36_real;
  assign data_reorder_9_imag = data_in_36_imag;
  assign data_reorder_41_real = data_in_37_real;
  assign data_reorder_41_imag = data_in_37_imag;
  assign data_reorder_25_real = data_in_38_real;
  assign data_reorder_25_imag = data_in_38_imag;
  assign data_reorder_57_real = data_in_39_real;
  assign data_reorder_57_imag = data_in_39_imag;
  assign data_reorder_5_real = data_in_40_real;
  assign data_reorder_5_imag = data_in_40_imag;
  assign data_reorder_37_real = data_in_41_real;
  assign data_reorder_37_imag = data_in_41_imag;
  assign data_reorder_21_real = data_in_42_real;
  assign data_reorder_21_imag = data_in_42_imag;
  assign data_reorder_53_real = data_in_43_real;
  assign data_reorder_53_imag = data_in_43_imag;
  assign data_reorder_13_real = data_in_44_real;
  assign data_reorder_13_imag = data_in_44_imag;
  assign data_reorder_45_real = data_in_45_real;
  assign data_reorder_45_imag = data_in_45_imag;
  assign data_reorder_29_real = data_in_46_real;
  assign data_reorder_29_imag = data_in_46_imag;
  assign data_reorder_61_real = data_in_47_real;
  assign data_reorder_61_imag = data_in_47_imag;
  assign data_reorder_3_real = data_in_48_real;
  assign data_reorder_3_imag = data_in_48_imag;
  assign data_reorder_35_real = data_in_49_real;
  assign data_reorder_35_imag = data_in_49_imag;
  assign data_reorder_19_real = data_in_50_real;
  assign data_reorder_19_imag = data_in_50_imag;
  assign data_reorder_51_real = data_in_51_real;
  assign data_reorder_51_imag = data_in_51_imag;
  assign data_reorder_11_real = data_in_52_real;
  assign data_reorder_11_imag = data_in_52_imag;
  assign data_reorder_43_real = data_in_53_real;
  assign data_reorder_43_imag = data_in_53_imag;
  assign data_reorder_27_real = data_in_54_real;
  assign data_reorder_27_imag = data_in_54_imag;
  assign data_reorder_59_real = data_in_55_real;
  assign data_reorder_59_imag = data_in_55_imag;
  assign data_reorder_7_real = data_in_56_real;
  assign data_reorder_7_imag = data_in_56_imag;
  assign data_reorder_39_real = data_in_57_real;
  assign data_reorder_39_imag = data_in_57_imag;
  assign data_reorder_23_real = data_in_58_real;
  assign data_reorder_23_imag = data_in_58_imag;
  assign data_reorder_55_real = data_in_59_real;
  assign data_reorder_55_imag = data_in_59_imag;
  assign data_reorder_15_real = data_in_60_real;
  assign data_reorder_15_imag = data_in_60_imag;
  assign data_reorder_47_real = data_in_61_real;
  assign data_reorder_47_imag = data_in_61_imag;
  assign data_reorder_31_real = data_in_62_real;
  assign data_reorder_31_imag = data_in_62_imag;
  assign data_reorder_63_real = data_in_63_real;
  assign data_reorder_63_imag = data_in_63_imag;
  assign _zz_3 = ($signed(_zz_2113) * $signed(data_mid_0_1_real));
  assign _zz_961 = _zz_2114;
  assign _zz_1 = _zz_2117[35 : 0];
  assign _zz_962 = _zz_2118;
  assign _zz_2 = _zz_2121[35 : 0];
  assign _zz_4 = 1'b1;
  assign _zz_963 = _zz_2122;
  assign _zz_964 = _zz_2130;
  assign _zz_5 = 1'b1;
  assign _zz_965 = _zz_2138;
  assign _zz_966 = _zz_2146;
  assign _zz_8 = ($signed(_zz_2154) * $signed(data_mid_0_3_real));
  assign _zz_967 = _zz_2155;
  assign _zz_6 = _zz_2158[35 : 0];
  assign _zz_968 = _zz_2159;
  assign _zz_7 = _zz_2162[35 : 0];
  assign _zz_9 = 1'b1;
  assign _zz_969 = _zz_2163;
  assign _zz_970 = _zz_2171;
  assign _zz_10 = 1'b1;
  assign _zz_971 = _zz_2179;
  assign _zz_972 = _zz_2187;
  assign _zz_13 = ($signed(_zz_2195) * $signed(data_mid_0_5_real));
  assign _zz_973 = _zz_2196;
  assign _zz_11 = _zz_2199[35 : 0];
  assign _zz_974 = _zz_2200;
  assign _zz_12 = _zz_2203[35 : 0];
  assign _zz_14 = 1'b1;
  assign _zz_975 = _zz_2204;
  assign _zz_976 = _zz_2212;
  assign _zz_15 = 1'b1;
  assign _zz_977 = _zz_2220;
  assign _zz_978 = _zz_2228;
  assign _zz_18 = ($signed(_zz_2236) * $signed(data_mid_0_7_real));
  assign _zz_979 = _zz_2237;
  assign _zz_16 = _zz_2240[35 : 0];
  assign _zz_980 = _zz_2241;
  assign _zz_17 = _zz_2244[35 : 0];
  assign _zz_19 = 1'b1;
  assign _zz_981 = _zz_2245;
  assign _zz_982 = _zz_2253;
  assign _zz_20 = 1'b1;
  assign _zz_983 = _zz_2261;
  assign _zz_984 = _zz_2269;
  assign _zz_23 = ($signed(_zz_2277) * $signed(data_mid_0_9_real));
  assign _zz_985 = _zz_2278;
  assign _zz_21 = _zz_2281[35 : 0];
  assign _zz_986 = _zz_2282;
  assign _zz_22 = _zz_2285[35 : 0];
  assign _zz_24 = 1'b1;
  assign _zz_987 = _zz_2286;
  assign _zz_988 = _zz_2294;
  assign _zz_25 = 1'b1;
  assign _zz_989 = _zz_2302;
  assign _zz_990 = _zz_2310;
  assign _zz_28 = ($signed(_zz_2318) * $signed(data_mid_0_11_real));
  assign _zz_991 = _zz_2319;
  assign _zz_26 = _zz_2322[35 : 0];
  assign _zz_992 = _zz_2323;
  assign _zz_27 = _zz_2326[35 : 0];
  assign _zz_29 = 1'b1;
  assign _zz_993 = _zz_2327;
  assign _zz_994 = _zz_2335;
  assign _zz_30 = 1'b1;
  assign _zz_995 = _zz_2343;
  assign _zz_996 = _zz_2351;
  assign _zz_33 = ($signed(_zz_2359) * $signed(data_mid_0_13_real));
  assign _zz_997 = _zz_2360;
  assign _zz_31 = _zz_2363[35 : 0];
  assign _zz_998 = _zz_2364;
  assign _zz_32 = _zz_2367[35 : 0];
  assign _zz_34 = 1'b1;
  assign _zz_999 = _zz_2368;
  assign _zz_1000 = _zz_2376;
  assign _zz_35 = 1'b1;
  assign _zz_1001 = _zz_2384;
  assign _zz_1002 = _zz_2392;
  assign _zz_38 = ($signed(_zz_2400) * $signed(data_mid_0_15_real));
  assign _zz_1003 = _zz_2401;
  assign _zz_36 = _zz_2404[35 : 0];
  assign _zz_1004 = _zz_2405;
  assign _zz_37 = _zz_2408[35 : 0];
  assign _zz_39 = 1'b1;
  assign _zz_1005 = _zz_2409;
  assign _zz_1006 = _zz_2417;
  assign _zz_40 = 1'b1;
  assign _zz_1007 = _zz_2425;
  assign _zz_1008 = _zz_2433;
  assign _zz_43 = ($signed(_zz_2441) * $signed(data_mid_0_17_real));
  assign _zz_1009 = _zz_2442;
  assign _zz_41 = _zz_2445[35 : 0];
  assign _zz_1010 = _zz_2446;
  assign _zz_42 = _zz_2449[35 : 0];
  assign _zz_44 = 1'b1;
  assign _zz_1011 = _zz_2450;
  assign _zz_1012 = _zz_2458;
  assign _zz_45 = 1'b1;
  assign _zz_1013 = _zz_2466;
  assign _zz_1014 = _zz_2474;
  assign _zz_48 = ($signed(_zz_2482) * $signed(data_mid_0_19_real));
  assign _zz_1015 = _zz_2483;
  assign _zz_46 = _zz_2486[35 : 0];
  assign _zz_1016 = _zz_2487;
  assign _zz_47 = _zz_2490[35 : 0];
  assign _zz_49 = 1'b1;
  assign _zz_1017 = _zz_2491;
  assign _zz_1018 = _zz_2499;
  assign _zz_50 = 1'b1;
  assign _zz_1019 = _zz_2507;
  assign _zz_1020 = _zz_2515;
  assign _zz_53 = ($signed(_zz_2523) * $signed(data_mid_0_21_real));
  assign _zz_1021 = _zz_2524;
  assign _zz_51 = _zz_2527[35 : 0];
  assign _zz_1022 = _zz_2528;
  assign _zz_52 = _zz_2531[35 : 0];
  assign _zz_54 = 1'b1;
  assign _zz_1023 = _zz_2532;
  assign _zz_1024 = _zz_2540;
  assign _zz_55 = 1'b1;
  assign _zz_1025 = _zz_2548;
  assign _zz_1026 = _zz_2556;
  assign _zz_58 = ($signed(_zz_2564) * $signed(data_mid_0_23_real));
  assign _zz_1027 = _zz_2565;
  assign _zz_56 = _zz_2568[35 : 0];
  assign _zz_1028 = _zz_2569;
  assign _zz_57 = _zz_2572[35 : 0];
  assign _zz_59 = 1'b1;
  assign _zz_1029 = _zz_2573;
  assign _zz_1030 = _zz_2581;
  assign _zz_60 = 1'b1;
  assign _zz_1031 = _zz_2589;
  assign _zz_1032 = _zz_2597;
  assign _zz_63 = ($signed(_zz_2605) * $signed(data_mid_0_25_real));
  assign _zz_1033 = _zz_2606;
  assign _zz_61 = _zz_2609[35 : 0];
  assign _zz_1034 = _zz_2610;
  assign _zz_62 = _zz_2613[35 : 0];
  assign _zz_64 = 1'b1;
  assign _zz_1035 = _zz_2614;
  assign _zz_1036 = _zz_2622;
  assign _zz_65 = 1'b1;
  assign _zz_1037 = _zz_2630;
  assign _zz_1038 = _zz_2638;
  assign _zz_68 = ($signed(_zz_2646) * $signed(data_mid_0_27_real));
  assign _zz_1039 = _zz_2647;
  assign _zz_66 = _zz_2650[35 : 0];
  assign _zz_1040 = _zz_2651;
  assign _zz_67 = _zz_2654[35 : 0];
  assign _zz_69 = 1'b1;
  assign _zz_1041 = _zz_2655;
  assign _zz_1042 = _zz_2663;
  assign _zz_70 = 1'b1;
  assign _zz_1043 = _zz_2671;
  assign _zz_1044 = _zz_2679;
  assign _zz_73 = ($signed(_zz_2687) * $signed(data_mid_0_29_real));
  assign _zz_1045 = _zz_2688;
  assign _zz_71 = _zz_2691[35 : 0];
  assign _zz_1046 = _zz_2692;
  assign _zz_72 = _zz_2695[35 : 0];
  assign _zz_74 = 1'b1;
  assign _zz_1047 = _zz_2696;
  assign _zz_1048 = _zz_2704;
  assign _zz_75 = 1'b1;
  assign _zz_1049 = _zz_2712;
  assign _zz_1050 = _zz_2720;
  assign _zz_78 = ($signed(_zz_2728) * $signed(data_mid_0_31_real));
  assign _zz_1051 = _zz_2729;
  assign _zz_76 = _zz_2732[35 : 0];
  assign _zz_1052 = _zz_2733;
  assign _zz_77 = _zz_2736[35 : 0];
  assign _zz_79 = 1'b1;
  assign _zz_1053 = _zz_2737;
  assign _zz_1054 = _zz_2745;
  assign _zz_80 = 1'b1;
  assign _zz_1055 = _zz_2753;
  assign _zz_1056 = _zz_2761;
  assign _zz_83 = ($signed(_zz_2769) * $signed(data_mid_0_33_real));
  assign _zz_1057 = _zz_2770;
  assign _zz_81 = _zz_2773[35 : 0];
  assign _zz_1058 = _zz_2774;
  assign _zz_82 = _zz_2777[35 : 0];
  assign _zz_84 = 1'b1;
  assign _zz_1059 = _zz_2778;
  assign _zz_1060 = _zz_2786;
  assign _zz_85 = 1'b1;
  assign _zz_1061 = _zz_2794;
  assign _zz_1062 = _zz_2802;
  assign _zz_88 = ($signed(_zz_2810) * $signed(data_mid_0_35_real));
  assign _zz_1063 = _zz_2811;
  assign _zz_86 = _zz_2814[35 : 0];
  assign _zz_1064 = _zz_2815;
  assign _zz_87 = _zz_2818[35 : 0];
  assign _zz_89 = 1'b1;
  assign _zz_1065 = _zz_2819;
  assign _zz_1066 = _zz_2827;
  assign _zz_90 = 1'b1;
  assign _zz_1067 = _zz_2835;
  assign _zz_1068 = _zz_2843;
  assign _zz_93 = ($signed(_zz_2851) * $signed(data_mid_0_37_real));
  assign _zz_1069 = _zz_2852;
  assign _zz_91 = _zz_2855[35 : 0];
  assign _zz_1070 = _zz_2856;
  assign _zz_92 = _zz_2859[35 : 0];
  assign _zz_94 = 1'b1;
  assign _zz_1071 = _zz_2860;
  assign _zz_1072 = _zz_2868;
  assign _zz_95 = 1'b1;
  assign _zz_1073 = _zz_2876;
  assign _zz_1074 = _zz_2884;
  assign _zz_98 = ($signed(_zz_2892) * $signed(data_mid_0_39_real));
  assign _zz_1075 = _zz_2893;
  assign _zz_96 = _zz_2896[35 : 0];
  assign _zz_1076 = _zz_2897;
  assign _zz_97 = _zz_2900[35 : 0];
  assign _zz_99 = 1'b1;
  assign _zz_1077 = _zz_2901;
  assign _zz_1078 = _zz_2909;
  assign _zz_100 = 1'b1;
  assign _zz_1079 = _zz_2917;
  assign _zz_1080 = _zz_2925;
  assign _zz_103 = ($signed(_zz_2933) * $signed(data_mid_0_41_real));
  assign _zz_1081 = _zz_2934;
  assign _zz_101 = _zz_2937[35 : 0];
  assign _zz_1082 = _zz_2938;
  assign _zz_102 = _zz_2941[35 : 0];
  assign _zz_104 = 1'b1;
  assign _zz_1083 = _zz_2942;
  assign _zz_1084 = _zz_2950;
  assign _zz_105 = 1'b1;
  assign _zz_1085 = _zz_2958;
  assign _zz_1086 = _zz_2966;
  assign _zz_108 = ($signed(_zz_2974) * $signed(data_mid_0_43_real));
  assign _zz_1087 = _zz_2975;
  assign _zz_106 = _zz_2978[35 : 0];
  assign _zz_1088 = _zz_2979;
  assign _zz_107 = _zz_2982[35 : 0];
  assign _zz_109 = 1'b1;
  assign _zz_1089 = _zz_2983;
  assign _zz_1090 = _zz_2991;
  assign _zz_110 = 1'b1;
  assign _zz_1091 = _zz_2999;
  assign _zz_1092 = _zz_3007;
  assign _zz_113 = ($signed(_zz_3015) * $signed(data_mid_0_45_real));
  assign _zz_1093 = _zz_3016;
  assign _zz_111 = _zz_3019[35 : 0];
  assign _zz_1094 = _zz_3020;
  assign _zz_112 = _zz_3023[35 : 0];
  assign _zz_114 = 1'b1;
  assign _zz_1095 = _zz_3024;
  assign _zz_1096 = _zz_3032;
  assign _zz_115 = 1'b1;
  assign _zz_1097 = _zz_3040;
  assign _zz_1098 = _zz_3048;
  assign _zz_118 = ($signed(_zz_3056) * $signed(data_mid_0_47_real));
  assign _zz_1099 = _zz_3057;
  assign _zz_116 = _zz_3060[35 : 0];
  assign _zz_1100 = _zz_3061;
  assign _zz_117 = _zz_3064[35 : 0];
  assign _zz_119 = 1'b1;
  assign _zz_1101 = _zz_3065;
  assign _zz_1102 = _zz_3073;
  assign _zz_120 = 1'b1;
  assign _zz_1103 = _zz_3081;
  assign _zz_1104 = _zz_3089;
  assign _zz_123 = ($signed(_zz_3097) * $signed(data_mid_0_49_real));
  assign _zz_1105 = _zz_3098;
  assign _zz_121 = _zz_3101[35 : 0];
  assign _zz_1106 = _zz_3102;
  assign _zz_122 = _zz_3105[35 : 0];
  assign _zz_124 = 1'b1;
  assign _zz_1107 = _zz_3106;
  assign _zz_1108 = _zz_3114;
  assign _zz_125 = 1'b1;
  assign _zz_1109 = _zz_3122;
  assign _zz_1110 = _zz_3130;
  assign _zz_128 = ($signed(_zz_3138) * $signed(data_mid_0_51_real));
  assign _zz_1111 = _zz_3139;
  assign _zz_126 = _zz_3142[35 : 0];
  assign _zz_1112 = _zz_3143;
  assign _zz_127 = _zz_3146[35 : 0];
  assign _zz_129 = 1'b1;
  assign _zz_1113 = _zz_3147;
  assign _zz_1114 = _zz_3155;
  assign _zz_130 = 1'b1;
  assign _zz_1115 = _zz_3163;
  assign _zz_1116 = _zz_3171;
  assign _zz_133 = ($signed(_zz_3179) * $signed(data_mid_0_53_real));
  assign _zz_1117 = _zz_3180;
  assign _zz_131 = _zz_3183[35 : 0];
  assign _zz_1118 = _zz_3184;
  assign _zz_132 = _zz_3187[35 : 0];
  assign _zz_134 = 1'b1;
  assign _zz_1119 = _zz_3188;
  assign _zz_1120 = _zz_3196;
  assign _zz_135 = 1'b1;
  assign _zz_1121 = _zz_3204;
  assign _zz_1122 = _zz_3212;
  assign _zz_138 = ($signed(_zz_3220) * $signed(data_mid_0_55_real));
  assign _zz_1123 = _zz_3221;
  assign _zz_136 = _zz_3224[35 : 0];
  assign _zz_1124 = _zz_3225;
  assign _zz_137 = _zz_3228[35 : 0];
  assign _zz_139 = 1'b1;
  assign _zz_1125 = _zz_3229;
  assign _zz_1126 = _zz_3237;
  assign _zz_140 = 1'b1;
  assign _zz_1127 = _zz_3245;
  assign _zz_1128 = _zz_3253;
  assign _zz_143 = ($signed(_zz_3261) * $signed(data_mid_0_57_real));
  assign _zz_1129 = _zz_3262;
  assign _zz_141 = _zz_3265[35 : 0];
  assign _zz_1130 = _zz_3266;
  assign _zz_142 = _zz_3269[35 : 0];
  assign _zz_144 = 1'b1;
  assign _zz_1131 = _zz_3270;
  assign _zz_1132 = _zz_3278;
  assign _zz_145 = 1'b1;
  assign _zz_1133 = _zz_3286;
  assign _zz_1134 = _zz_3294;
  assign _zz_148 = ($signed(_zz_3302) * $signed(data_mid_0_59_real));
  assign _zz_1135 = _zz_3303;
  assign _zz_146 = _zz_3306[35 : 0];
  assign _zz_1136 = _zz_3307;
  assign _zz_147 = _zz_3310[35 : 0];
  assign _zz_149 = 1'b1;
  assign _zz_1137 = _zz_3311;
  assign _zz_1138 = _zz_3319;
  assign _zz_150 = 1'b1;
  assign _zz_1139 = _zz_3327;
  assign _zz_1140 = _zz_3335;
  assign _zz_153 = ($signed(_zz_3343) * $signed(data_mid_0_61_real));
  assign _zz_1141 = _zz_3344;
  assign _zz_151 = _zz_3347[35 : 0];
  assign _zz_1142 = _zz_3348;
  assign _zz_152 = _zz_3351[35 : 0];
  assign _zz_154 = 1'b1;
  assign _zz_1143 = _zz_3352;
  assign _zz_1144 = _zz_3360;
  assign _zz_155 = 1'b1;
  assign _zz_1145 = _zz_3368;
  assign _zz_1146 = _zz_3376;
  assign _zz_158 = ($signed(_zz_3384) * $signed(data_mid_0_63_real));
  assign _zz_1147 = _zz_3385;
  assign _zz_156 = _zz_3388[35 : 0];
  assign _zz_1148 = _zz_3389;
  assign _zz_157 = _zz_3392[35 : 0];
  assign _zz_159 = 1'b1;
  assign _zz_1149 = _zz_3393;
  assign _zz_1150 = _zz_3401;
  assign _zz_160 = 1'b1;
  assign _zz_1151 = _zz_3409;
  assign _zz_1152 = _zz_3417;
  assign _zz_163 = ($signed(_zz_3425) * $signed(data_mid_1_2_real));
  assign _zz_1153 = _zz_3426;
  assign _zz_161 = _zz_3429[35 : 0];
  assign _zz_1154 = _zz_3430;
  assign _zz_162 = _zz_3433[35 : 0];
  assign _zz_164 = 1'b1;
  assign _zz_1155 = _zz_3434;
  assign _zz_1156 = _zz_3442;
  assign _zz_165 = 1'b1;
  assign _zz_1157 = _zz_3450;
  assign _zz_1158 = _zz_3458;
  assign _zz_168 = ($signed(_zz_3466) * $signed(data_mid_1_3_real));
  assign _zz_1159 = _zz_3467;
  assign _zz_166 = _zz_3470[35 : 0];
  assign _zz_1160 = _zz_3471;
  assign _zz_167 = _zz_3474[35 : 0];
  assign _zz_169 = 1'b1;
  assign _zz_1161 = _zz_3475;
  assign _zz_1162 = _zz_3483;
  assign _zz_170 = 1'b1;
  assign _zz_1163 = _zz_3491;
  assign _zz_1164 = _zz_3499;
  assign _zz_173 = ($signed(_zz_3507) * $signed(data_mid_1_6_real));
  assign _zz_1165 = _zz_3508;
  assign _zz_171 = _zz_3511[35 : 0];
  assign _zz_1166 = _zz_3512;
  assign _zz_172 = _zz_3515[35 : 0];
  assign _zz_174 = 1'b1;
  assign _zz_1167 = _zz_3516;
  assign _zz_1168 = _zz_3524;
  assign _zz_175 = 1'b1;
  assign _zz_1169 = _zz_3532;
  assign _zz_1170 = _zz_3540;
  assign _zz_178 = ($signed(_zz_3548) * $signed(data_mid_1_7_real));
  assign _zz_1171 = _zz_3549;
  assign _zz_176 = _zz_3552[35 : 0];
  assign _zz_1172 = _zz_3553;
  assign _zz_177 = _zz_3556[35 : 0];
  assign _zz_179 = 1'b1;
  assign _zz_1173 = _zz_3557;
  assign _zz_1174 = _zz_3565;
  assign _zz_180 = 1'b1;
  assign _zz_1175 = _zz_3573;
  assign _zz_1176 = _zz_3581;
  assign _zz_183 = ($signed(_zz_3589) * $signed(data_mid_1_10_real));
  assign _zz_1177 = _zz_3590;
  assign _zz_181 = _zz_3593[35 : 0];
  assign _zz_1178 = _zz_3594;
  assign _zz_182 = _zz_3597[35 : 0];
  assign _zz_184 = 1'b1;
  assign _zz_1179 = _zz_3598;
  assign _zz_1180 = _zz_3606;
  assign _zz_185 = 1'b1;
  assign _zz_1181 = _zz_3614;
  assign _zz_1182 = _zz_3622;
  assign _zz_188 = ($signed(_zz_3630) * $signed(data_mid_1_11_real));
  assign _zz_1183 = _zz_3631;
  assign _zz_186 = _zz_3634[35 : 0];
  assign _zz_1184 = _zz_3635;
  assign _zz_187 = _zz_3638[35 : 0];
  assign _zz_189 = 1'b1;
  assign _zz_1185 = _zz_3639;
  assign _zz_1186 = _zz_3647;
  assign _zz_190 = 1'b1;
  assign _zz_1187 = _zz_3655;
  assign _zz_1188 = _zz_3663;
  assign _zz_193 = ($signed(_zz_3671) * $signed(data_mid_1_14_real));
  assign _zz_1189 = _zz_3672;
  assign _zz_191 = _zz_3675[35 : 0];
  assign _zz_1190 = _zz_3676;
  assign _zz_192 = _zz_3679[35 : 0];
  assign _zz_194 = 1'b1;
  assign _zz_1191 = _zz_3680;
  assign _zz_1192 = _zz_3688;
  assign _zz_195 = 1'b1;
  assign _zz_1193 = _zz_3696;
  assign _zz_1194 = _zz_3704;
  assign _zz_198 = ($signed(_zz_3712) * $signed(data_mid_1_15_real));
  assign _zz_1195 = _zz_3713;
  assign _zz_196 = _zz_3716[35 : 0];
  assign _zz_1196 = _zz_3717;
  assign _zz_197 = _zz_3720[35 : 0];
  assign _zz_199 = 1'b1;
  assign _zz_1197 = _zz_3721;
  assign _zz_1198 = _zz_3729;
  assign _zz_200 = 1'b1;
  assign _zz_1199 = _zz_3737;
  assign _zz_1200 = _zz_3745;
  assign _zz_203 = ($signed(_zz_3753) * $signed(data_mid_1_18_real));
  assign _zz_1201 = _zz_3754;
  assign _zz_201 = _zz_3757[35 : 0];
  assign _zz_1202 = _zz_3758;
  assign _zz_202 = _zz_3761[35 : 0];
  assign _zz_204 = 1'b1;
  assign _zz_1203 = _zz_3762;
  assign _zz_1204 = _zz_3770;
  assign _zz_205 = 1'b1;
  assign _zz_1205 = _zz_3778;
  assign _zz_1206 = _zz_3786;
  assign _zz_208 = ($signed(_zz_3794) * $signed(data_mid_1_19_real));
  assign _zz_1207 = _zz_3795;
  assign _zz_206 = _zz_3798[35 : 0];
  assign _zz_1208 = _zz_3799;
  assign _zz_207 = _zz_3802[35 : 0];
  assign _zz_209 = 1'b1;
  assign _zz_1209 = _zz_3803;
  assign _zz_1210 = _zz_3811;
  assign _zz_210 = 1'b1;
  assign _zz_1211 = _zz_3819;
  assign _zz_1212 = _zz_3827;
  assign _zz_213 = ($signed(_zz_3835) * $signed(data_mid_1_22_real));
  assign _zz_1213 = _zz_3836;
  assign _zz_211 = _zz_3839[35 : 0];
  assign _zz_1214 = _zz_3840;
  assign _zz_212 = _zz_3843[35 : 0];
  assign _zz_214 = 1'b1;
  assign _zz_1215 = _zz_3844;
  assign _zz_1216 = _zz_3852;
  assign _zz_215 = 1'b1;
  assign _zz_1217 = _zz_3860;
  assign _zz_1218 = _zz_3868;
  assign _zz_218 = ($signed(_zz_3876) * $signed(data_mid_1_23_real));
  assign _zz_1219 = _zz_3877;
  assign _zz_216 = _zz_3880[35 : 0];
  assign _zz_1220 = _zz_3881;
  assign _zz_217 = _zz_3884[35 : 0];
  assign _zz_219 = 1'b1;
  assign _zz_1221 = _zz_3885;
  assign _zz_1222 = _zz_3893;
  assign _zz_220 = 1'b1;
  assign _zz_1223 = _zz_3901;
  assign _zz_1224 = _zz_3909;
  assign _zz_223 = ($signed(_zz_3917) * $signed(data_mid_1_26_real));
  assign _zz_1225 = _zz_3918;
  assign _zz_221 = _zz_3921[35 : 0];
  assign _zz_1226 = _zz_3922;
  assign _zz_222 = _zz_3925[35 : 0];
  assign _zz_224 = 1'b1;
  assign _zz_1227 = _zz_3926;
  assign _zz_1228 = _zz_3934;
  assign _zz_225 = 1'b1;
  assign _zz_1229 = _zz_3942;
  assign _zz_1230 = _zz_3950;
  assign _zz_228 = ($signed(_zz_3958) * $signed(data_mid_1_27_real));
  assign _zz_1231 = _zz_3959;
  assign _zz_226 = _zz_3962[35 : 0];
  assign _zz_1232 = _zz_3963;
  assign _zz_227 = _zz_3966[35 : 0];
  assign _zz_229 = 1'b1;
  assign _zz_1233 = _zz_3967;
  assign _zz_1234 = _zz_3975;
  assign _zz_230 = 1'b1;
  assign _zz_1235 = _zz_3983;
  assign _zz_1236 = _zz_3991;
  assign _zz_233 = ($signed(_zz_3999) * $signed(data_mid_1_30_real));
  assign _zz_1237 = _zz_4000;
  assign _zz_231 = _zz_4003[35 : 0];
  assign _zz_1238 = _zz_4004;
  assign _zz_232 = _zz_4007[35 : 0];
  assign _zz_234 = 1'b1;
  assign _zz_1239 = _zz_4008;
  assign _zz_1240 = _zz_4016;
  assign _zz_235 = 1'b1;
  assign _zz_1241 = _zz_4024;
  assign _zz_1242 = _zz_4032;
  assign _zz_238 = ($signed(_zz_4040) * $signed(data_mid_1_31_real));
  assign _zz_1243 = _zz_4041;
  assign _zz_236 = _zz_4044[35 : 0];
  assign _zz_1244 = _zz_4045;
  assign _zz_237 = _zz_4048[35 : 0];
  assign _zz_239 = 1'b1;
  assign _zz_1245 = _zz_4049;
  assign _zz_1246 = _zz_4057;
  assign _zz_240 = 1'b1;
  assign _zz_1247 = _zz_4065;
  assign _zz_1248 = _zz_4073;
  assign _zz_243 = ($signed(_zz_4081) * $signed(data_mid_1_34_real));
  assign _zz_1249 = _zz_4082;
  assign _zz_241 = _zz_4085[35 : 0];
  assign _zz_1250 = _zz_4086;
  assign _zz_242 = _zz_4089[35 : 0];
  assign _zz_244 = 1'b1;
  assign _zz_1251 = _zz_4090;
  assign _zz_1252 = _zz_4098;
  assign _zz_245 = 1'b1;
  assign _zz_1253 = _zz_4106;
  assign _zz_1254 = _zz_4114;
  assign _zz_248 = ($signed(_zz_4122) * $signed(data_mid_1_35_real));
  assign _zz_1255 = _zz_4123;
  assign _zz_246 = _zz_4126[35 : 0];
  assign _zz_1256 = _zz_4127;
  assign _zz_247 = _zz_4130[35 : 0];
  assign _zz_249 = 1'b1;
  assign _zz_1257 = _zz_4131;
  assign _zz_1258 = _zz_4139;
  assign _zz_250 = 1'b1;
  assign _zz_1259 = _zz_4147;
  assign _zz_1260 = _zz_4155;
  assign _zz_253 = ($signed(_zz_4163) * $signed(data_mid_1_38_real));
  assign _zz_1261 = _zz_4164;
  assign _zz_251 = _zz_4167[35 : 0];
  assign _zz_1262 = _zz_4168;
  assign _zz_252 = _zz_4171[35 : 0];
  assign _zz_254 = 1'b1;
  assign _zz_1263 = _zz_4172;
  assign _zz_1264 = _zz_4180;
  assign _zz_255 = 1'b1;
  assign _zz_1265 = _zz_4188;
  assign _zz_1266 = _zz_4196;
  assign _zz_258 = ($signed(_zz_4204) * $signed(data_mid_1_39_real));
  assign _zz_1267 = _zz_4205;
  assign _zz_256 = _zz_4208[35 : 0];
  assign _zz_1268 = _zz_4209;
  assign _zz_257 = _zz_4212[35 : 0];
  assign _zz_259 = 1'b1;
  assign _zz_1269 = _zz_4213;
  assign _zz_1270 = _zz_4221;
  assign _zz_260 = 1'b1;
  assign _zz_1271 = _zz_4229;
  assign _zz_1272 = _zz_4237;
  assign _zz_263 = ($signed(_zz_4245) * $signed(data_mid_1_42_real));
  assign _zz_1273 = _zz_4246;
  assign _zz_261 = _zz_4249[35 : 0];
  assign _zz_1274 = _zz_4250;
  assign _zz_262 = _zz_4253[35 : 0];
  assign _zz_264 = 1'b1;
  assign _zz_1275 = _zz_4254;
  assign _zz_1276 = _zz_4262;
  assign _zz_265 = 1'b1;
  assign _zz_1277 = _zz_4270;
  assign _zz_1278 = _zz_4278;
  assign _zz_268 = ($signed(_zz_4286) * $signed(data_mid_1_43_real));
  assign _zz_1279 = _zz_4287;
  assign _zz_266 = _zz_4290[35 : 0];
  assign _zz_1280 = _zz_4291;
  assign _zz_267 = _zz_4294[35 : 0];
  assign _zz_269 = 1'b1;
  assign _zz_1281 = _zz_4295;
  assign _zz_1282 = _zz_4303;
  assign _zz_270 = 1'b1;
  assign _zz_1283 = _zz_4311;
  assign _zz_1284 = _zz_4319;
  assign _zz_273 = ($signed(_zz_4327) * $signed(data_mid_1_46_real));
  assign _zz_1285 = _zz_4328;
  assign _zz_271 = _zz_4331[35 : 0];
  assign _zz_1286 = _zz_4332;
  assign _zz_272 = _zz_4335[35 : 0];
  assign _zz_274 = 1'b1;
  assign _zz_1287 = _zz_4336;
  assign _zz_1288 = _zz_4344;
  assign _zz_275 = 1'b1;
  assign _zz_1289 = _zz_4352;
  assign _zz_1290 = _zz_4360;
  assign _zz_278 = ($signed(_zz_4368) * $signed(data_mid_1_47_real));
  assign _zz_1291 = _zz_4369;
  assign _zz_276 = _zz_4372[35 : 0];
  assign _zz_1292 = _zz_4373;
  assign _zz_277 = _zz_4376[35 : 0];
  assign _zz_279 = 1'b1;
  assign _zz_1293 = _zz_4377;
  assign _zz_1294 = _zz_4385;
  assign _zz_280 = 1'b1;
  assign _zz_1295 = _zz_4393;
  assign _zz_1296 = _zz_4401;
  assign _zz_283 = ($signed(_zz_4409) * $signed(data_mid_1_50_real));
  assign _zz_1297 = _zz_4410;
  assign _zz_281 = _zz_4413[35 : 0];
  assign _zz_1298 = _zz_4414;
  assign _zz_282 = _zz_4417[35 : 0];
  assign _zz_284 = 1'b1;
  assign _zz_1299 = _zz_4418;
  assign _zz_1300 = _zz_4426;
  assign _zz_285 = 1'b1;
  assign _zz_1301 = _zz_4434;
  assign _zz_1302 = _zz_4442;
  assign _zz_288 = ($signed(_zz_4450) * $signed(data_mid_1_51_real));
  assign _zz_1303 = _zz_4451;
  assign _zz_286 = _zz_4454[35 : 0];
  assign _zz_1304 = _zz_4455;
  assign _zz_287 = _zz_4458[35 : 0];
  assign _zz_289 = 1'b1;
  assign _zz_1305 = _zz_4459;
  assign _zz_1306 = _zz_4467;
  assign _zz_290 = 1'b1;
  assign _zz_1307 = _zz_4475;
  assign _zz_1308 = _zz_4483;
  assign _zz_293 = ($signed(_zz_4491) * $signed(data_mid_1_54_real));
  assign _zz_1309 = _zz_4492;
  assign _zz_291 = _zz_4495[35 : 0];
  assign _zz_1310 = _zz_4496;
  assign _zz_292 = _zz_4499[35 : 0];
  assign _zz_294 = 1'b1;
  assign _zz_1311 = _zz_4500;
  assign _zz_1312 = _zz_4508;
  assign _zz_295 = 1'b1;
  assign _zz_1313 = _zz_4516;
  assign _zz_1314 = _zz_4524;
  assign _zz_298 = ($signed(_zz_4532) * $signed(data_mid_1_55_real));
  assign _zz_1315 = _zz_4533;
  assign _zz_296 = _zz_4536[35 : 0];
  assign _zz_1316 = _zz_4537;
  assign _zz_297 = _zz_4540[35 : 0];
  assign _zz_299 = 1'b1;
  assign _zz_1317 = _zz_4541;
  assign _zz_1318 = _zz_4549;
  assign _zz_300 = 1'b1;
  assign _zz_1319 = _zz_4557;
  assign _zz_1320 = _zz_4565;
  assign _zz_303 = ($signed(_zz_4573) * $signed(data_mid_1_58_real));
  assign _zz_1321 = _zz_4574;
  assign _zz_301 = _zz_4577[35 : 0];
  assign _zz_1322 = _zz_4578;
  assign _zz_302 = _zz_4581[35 : 0];
  assign _zz_304 = 1'b1;
  assign _zz_1323 = _zz_4582;
  assign _zz_1324 = _zz_4590;
  assign _zz_305 = 1'b1;
  assign _zz_1325 = _zz_4598;
  assign _zz_1326 = _zz_4606;
  assign _zz_308 = ($signed(_zz_4614) * $signed(data_mid_1_59_real));
  assign _zz_1327 = _zz_4615;
  assign _zz_306 = _zz_4618[35 : 0];
  assign _zz_1328 = _zz_4619;
  assign _zz_307 = _zz_4622[35 : 0];
  assign _zz_309 = 1'b1;
  assign _zz_1329 = _zz_4623;
  assign _zz_1330 = _zz_4631;
  assign _zz_310 = 1'b1;
  assign _zz_1331 = _zz_4639;
  assign _zz_1332 = _zz_4647;
  assign _zz_313 = ($signed(_zz_4655) * $signed(data_mid_1_62_real));
  assign _zz_1333 = _zz_4656;
  assign _zz_311 = _zz_4659[35 : 0];
  assign _zz_1334 = _zz_4660;
  assign _zz_312 = _zz_4663[35 : 0];
  assign _zz_314 = 1'b1;
  assign _zz_1335 = _zz_4664;
  assign _zz_1336 = _zz_4672;
  assign _zz_315 = 1'b1;
  assign _zz_1337 = _zz_4680;
  assign _zz_1338 = _zz_4688;
  assign _zz_318 = ($signed(_zz_4696) * $signed(data_mid_1_63_real));
  assign _zz_1339 = _zz_4697;
  assign _zz_316 = _zz_4700[35 : 0];
  assign _zz_1340 = _zz_4701;
  assign _zz_317 = _zz_4704[35 : 0];
  assign _zz_319 = 1'b1;
  assign _zz_1341 = _zz_4705;
  assign _zz_1342 = _zz_4713;
  assign _zz_320 = 1'b1;
  assign _zz_1343 = _zz_4721;
  assign _zz_1344 = _zz_4729;
  assign _zz_323 = ($signed(_zz_4737) * $signed(data_mid_2_4_real));
  assign _zz_1345 = _zz_4738;
  assign _zz_321 = _zz_4741[35 : 0];
  assign _zz_1346 = _zz_4742;
  assign _zz_322 = _zz_4745[35 : 0];
  assign _zz_324 = 1'b1;
  assign _zz_1347 = _zz_4746;
  assign _zz_1348 = _zz_4754;
  assign _zz_325 = 1'b1;
  assign _zz_1349 = _zz_4762;
  assign _zz_1350 = _zz_4770;
  assign _zz_328 = ($signed(_zz_4778) * $signed(data_mid_2_5_real));
  assign _zz_1351 = _zz_4779;
  assign _zz_326 = _zz_4782[35 : 0];
  assign _zz_1352 = _zz_4783;
  assign _zz_327 = _zz_4786[35 : 0];
  assign _zz_329 = 1'b1;
  assign _zz_1353 = _zz_4787;
  assign _zz_1354 = _zz_4795;
  assign _zz_330 = 1'b1;
  assign _zz_1355 = _zz_4803;
  assign _zz_1356 = _zz_4811;
  assign _zz_333 = ($signed(_zz_4819) * $signed(data_mid_2_6_real));
  assign _zz_1357 = _zz_4820;
  assign _zz_331 = _zz_4823[35 : 0];
  assign _zz_1358 = _zz_4824;
  assign _zz_332 = _zz_4827[35 : 0];
  assign _zz_334 = 1'b1;
  assign _zz_1359 = _zz_4828;
  assign _zz_1360 = _zz_4836;
  assign _zz_335 = 1'b1;
  assign _zz_1361 = _zz_4844;
  assign _zz_1362 = _zz_4852;
  assign _zz_338 = ($signed(_zz_4860) * $signed(data_mid_2_7_real));
  assign _zz_1363 = _zz_4861;
  assign _zz_336 = _zz_4864[35 : 0];
  assign _zz_1364 = _zz_4865;
  assign _zz_337 = _zz_4868[35 : 0];
  assign _zz_339 = 1'b1;
  assign _zz_1365 = _zz_4869;
  assign _zz_1366 = _zz_4877;
  assign _zz_340 = 1'b1;
  assign _zz_1367 = _zz_4885;
  assign _zz_1368 = _zz_4893;
  assign _zz_343 = ($signed(_zz_4901) * $signed(data_mid_2_12_real));
  assign _zz_1369 = _zz_4902;
  assign _zz_341 = _zz_4905[35 : 0];
  assign _zz_1370 = _zz_4906;
  assign _zz_342 = _zz_4909[35 : 0];
  assign _zz_344 = 1'b1;
  assign _zz_1371 = _zz_4910;
  assign _zz_1372 = _zz_4918;
  assign _zz_345 = 1'b1;
  assign _zz_1373 = _zz_4926;
  assign _zz_1374 = _zz_4934;
  assign _zz_348 = ($signed(_zz_4942) * $signed(data_mid_2_13_real));
  assign _zz_1375 = _zz_4943;
  assign _zz_346 = _zz_4946[35 : 0];
  assign _zz_1376 = _zz_4947;
  assign _zz_347 = _zz_4950[35 : 0];
  assign _zz_349 = 1'b1;
  assign _zz_1377 = _zz_4951;
  assign _zz_1378 = _zz_4959;
  assign _zz_350 = 1'b1;
  assign _zz_1379 = _zz_4967;
  assign _zz_1380 = _zz_4975;
  assign _zz_353 = ($signed(_zz_4983) * $signed(data_mid_2_14_real));
  assign _zz_1381 = _zz_4984;
  assign _zz_351 = _zz_4987[35 : 0];
  assign _zz_1382 = _zz_4988;
  assign _zz_352 = _zz_4991[35 : 0];
  assign _zz_354 = 1'b1;
  assign _zz_1383 = _zz_4992;
  assign _zz_1384 = _zz_5000;
  assign _zz_355 = 1'b1;
  assign _zz_1385 = _zz_5008;
  assign _zz_1386 = _zz_5016;
  assign _zz_358 = ($signed(_zz_5024) * $signed(data_mid_2_15_real));
  assign _zz_1387 = _zz_5025;
  assign _zz_356 = _zz_5028[35 : 0];
  assign _zz_1388 = _zz_5029;
  assign _zz_357 = _zz_5032[35 : 0];
  assign _zz_359 = 1'b1;
  assign _zz_1389 = _zz_5033;
  assign _zz_1390 = _zz_5041;
  assign _zz_360 = 1'b1;
  assign _zz_1391 = _zz_5049;
  assign _zz_1392 = _zz_5057;
  assign _zz_363 = ($signed(_zz_5065) * $signed(data_mid_2_20_real));
  assign _zz_1393 = _zz_5066;
  assign _zz_361 = _zz_5069[35 : 0];
  assign _zz_1394 = _zz_5070;
  assign _zz_362 = _zz_5073[35 : 0];
  assign _zz_364 = 1'b1;
  assign _zz_1395 = _zz_5074;
  assign _zz_1396 = _zz_5082;
  assign _zz_365 = 1'b1;
  assign _zz_1397 = _zz_5090;
  assign _zz_1398 = _zz_5098;
  assign _zz_368 = ($signed(_zz_5106) * $signed(data_mid_2_21_real));
  assign _zz_1399 = _zz_5107;
  assign _zz_366 = _zz_5110[35 : 0];
  assign _zz_1400 = _zz_5111;
  assign _zz_367 = _zz_5114[35 : 0];
  assign _zz_369 = 1'b1;
  assign _zz_1401 = _zz_5115;
  assign _zz_1402 = _zz_5123;
  assign _zz_370 = 1'b1;
  assign _zz_1403 = _zz_5131;
  assign _zz_1404 = _zz_5139;
  assign _zz_373 = ($signed(_zz_5147) * $signed(data_mid_2_22_real));
  assign _zz_1405 = _zz_5148;
  assign _zz_371 = _zz_5151[35 : 0];
  assign _zz_1406 = _zz_5152;
  assign _zz_372 = _zz_5155[35 : 0];
  assign _zz_374 = 1'b1;
  assign _zz_1407 = _zz_5156;
  assign _zz_1408 = _zz_5164;
  assign _zz_375 = 1'b1;
  assign _zz_1409 = _zz_5172;
  assign _zz_1410 = _zz_5180;
  assign _zz_378 = ($signed(_zz_5188) * $signed(data_mid_2_23_real));
  assign _zz_1411 = _zz_5189;
  assign _zz_376 = _zz_5192[35 : 0];
  assign _zz_1412 = _zz_5193;
  assign _zz_377 = _zz_5196[35 : 0];
  assign _zz_379 = 1'b1;
  assign _zz_1413 = _zz_5197;
  assign _zz_1414 = _zz_5205;
  assign _zz_380 = 1'b1;
  assign _zz_1415 = _zz_5213;
  assign _zz_1416 = _zz_5221;
  assign _zz_383 = ($signed(_zz_5229) * $signed(data_mid_2_28_real));
  assign _zz_1417 = _zz_5230;
  assign _zz_381 = _zz_5233[35 : 0];
  assign _zz_1418 = _zz_5234;
  assign _zz_382 = _zz_5237[35 : 0];
  assign _zz_384 = 1'b1;
  assign _zz_1419 = _zz_5238;
  assign _zz_1420 = _zz_5246;
  assign _zz_385 = 1'b1;
  assign _zz_1421 = _zz_5254;
  assign _zz_1422 = _zz_5262;
  assign _zz_388 = ($signed(_zz_5270) * $signed(data_mid_2_29_real));
  assign _zz_1423 = _zz_5271;
  assign _zz_386 = _zz_5274[35 : 0];
  assign _zz_1424 = _zz_5275;
  assign _zz_387 = _zz_5278[35 : 0];
  assign _zz_389 = 1'b1;
  assign _zz_1425 = _zz_5279;
  assign _zz_1426 = _zz_5287;
  assign _zz_390 = 1'b1;
  assign _zz_1427 = _zz_5295;
  assign _zz_1428 = _zz_5303;
  assign _zz_393 = ($signed(_zz_5311) * $signed(data_mid_2_30_real));
  assign _zz_1429 = _zz_5312;
  assign _zz_391 = _zz_5315[35 : 0];
  assign _zz_1430 = _zz_5316;
  assign _zz_392 = _zz_5319[35 : 0];
  assign _zz_394 = 1'b1;
  assign _zz_1431 = _zz_5320;
  assign _zz_1432 = _zz_5328;
  assign _zz_395 = 1'b1;
  assign _zz_1433 = _zz_5336;
  assign _zz_1434 = _zz_5344;
  assign _zz_398 = ($signed(_zz_5352) * $signed(data_mid_2_31_real));
  assign _zz_1435 = _zz_5353;
  assign _zz_396 = _zz_5356[35 : 0];
  assign _zz_1436 = _zz_5357;
  assign _zz_397 = _zz_5360[35 : 0];
  assign _zz_399 = 1'b1;
  assign _zz_1437 = _zz_5361;
  assign _zz_1438 = _zz_5369;
  assign _zz_400 = 1'b1;
  assign _zz_1439 = _zz_5377;
  assign _zz_1440 = _zz_5385;
  assign _zz_403 = ($signed(_zz_5393) * $signed(data_mid_2_36_real));
  assign _zz_1441 = _zz_5394;
  assign _zz_401 = _zz_5397[35 : 0];
  assign _zz_1442 = _zz_5398;
  assign _zz_402 = _zz_5401[35 : 0];
  assign _zz_404 = 1'b1;
  assign _zz_1443 = _zz_5402;
  assign _zz_1444 = _zz_5410;
  assign _zz_405 = 1'b1;
  assign _zz_1445 = _zz_5418;
  assign _zz_1446 = _zz_5426;
  assign _zz_408 = ($signed(_zz_5434) * $signed(data_mid_2_37_real));
  assign _zz_1447 = _zz_5435;
  assign _zz_406 = _zz_5438[35 : 0];
  assign _zz_1448 = _zz_5439;
  assign _zz_407 = _zz_5442[35 : 0];
  assign _zz_409 = 1'b1;
  assign _zz_1449 = _zz_5443;
  assign _zz_1450 = _zz_5451;
  assign _zz_410 = 1'b1;
  assign _zz_1451 = _zz_5459;
  assign _zz_1452 = _zz_5467;
  assign _zz_413 = ($signed(_zz_5475) * $signed(data_mid_2_38_real));
  assign _zz_1453 = _zz_5476;
  assign _zz_411 = _zz_5479[35 : 0];
  assign _zz_1454 = _zz_5480;
  assign _zz_412 = _zz_5483[35 : 0];
  assign _zz_414 = 1'b1;
  assign _zz_1455 = _zz_5484;
  assign _zz_1456 = _zz_5492;
  assign _zz_415 = 1'b1;
  assign _zz_1457 = _zz_5500;
  assign _zz_1458 = _zz_5508;
  assign _zz_418 = ($signed(_zz_5516) * $signed(data_mid_2_39_real));
  assign _zz_1459 = _zz_5517;
  assign _zz_416 = _zz_5520[35 : 0];
  assign _zz_1460 = _zz_5521;
  assign _zz_417 = _zz_5524[35 : 0];
  assign _zz_419 = 1'b1;
  assign _zz_1461 = _zz_5525;
  assign _zz_1462 = _zz_5533;
  assign _zz_420 = 1'b1;
  assign _zz_1463 = _zz_5541;
  assign _zz_1464 = _zz_5549;
  assign _zz_423 = ($signed(_zz_5557) * $signed(data_mid_2_44_real));
  assign _zz_1465 = _zz_5558;
  assign _zz_421 = _zz_5561[35 : 0];
  assign _zz_1466 = _zz_5562;
  assign _zz_422 = _zz_5565[35 : 0];
  assign _zz_424 = 1'b1;
  assign _zz_1467 = _zz_5566;
  assign _zz_1468 = _zz_5574;
  assign _zz_425 = 1'b1;
  assign _zz_1469 = _zz_5582;
  assign _zz_1470 = _zz_5590;
  assign _zz_428 = ($signed(_zz_5598) * $signed(data_mid_2_45_real));
  assign _zz_1471 = _zz_5599;
  assign _zz_426 = _zz_5602[35 : 0];
  assign _zz_1472 = _zz_5603;
  assign _zz_427 = _zz_5606[35 : 0];
  assign _zz_429 = 1'b1;
  assign _zz_1473 = _zz_5607;
  assign _zz_1474 = _zz_5615;
  assign _zz_430 = 1'b1;
  assign _zz_1475 = _zz_5623;
  assign _zz_1476 = _zz_5631;
  assign _zz_433 = ($signed(_zz_5639) * $signed(data_mid_2_46_real));
  assign _zz_1477 = _zz_5640;
  assign _zz_431 = _zz_5643[35 : 0];
  assign _zz_1478 = _zz_5644;
  assign _zz_432 = _zz_5647[35 : 0];
  assign _zz_434 = 1'b1;
  assign _zz_1479 = _zz_5648;
  assign _zz_1480 = _zz_5656;
  assign _zz_435 = 1'b1;
  assign _zz_1481 = _zz_5664;
  assign _zz_1482 = _zz_5672;
  assign _zz_438 = ($signed(_zz_5680) * $signed(data_mid_2_47_real));
  assign _zz_1483 = _zz_5681;
  assign _zz_436 = _zz_5684[35 : 0];
  assign _zz_1484 = _zz_5685;
  assign _zz_437 = _zz_5688[35 : 0];
  assign _zz_439 = 1'b1;
  assign _zz_1485 = _zz_5689;
  assign _zz_1486 = _zz_5697;
  assign _zz_440 = 1'b1;
  assign _zz_1487 = _zz_5705;
  assign _zz_1488 = _zz_5713;
  assign _zz_443 = ($signed(_zz_5721) * $signed(data_mid_2_52_real));
  assign _zz_1489 = _zz_5722;
  assign _zz_441 = _zz_5725[35 : 0];
  assign _zz_1490 = _zz_5726;
  assign _zz_442 = _zz_5729[35 : 0];
  assign _zz_444 = 1'b1;
  assign _zz_1491 = _zz_5730;
  assign _zz_1492 = _zz_5738;
  assign _zz_445 = 1'b1;
  assign _zz_1493 = _zz_5746;
  assign _zz_1494 = _zz_5754;
  assign _zz_448 = ($signed(_zz_5762) * $signed(data_mid_2_53_real));
  assign _zz_1495 = _zz_5763;
  assign _zz_446 = _zz_5766[35 : 0];
  assign _zz_1496 = _zz_5767;
  assign _zz_447 = _zz_5770[35 : 0];
  assign _zz_449 = 1'b1;
  assign _zz_1497 = _zz_5771;
  assign _zz_1498 = _zz_5779;
  assign _zz_450 = 1'b1;
  assign _zz_1499 = _zz_5787;
  assign _zz_1500 = _zz_5795;
  assign _zz_453 = ($signed(_zz_5803) * $signed(data_mid_2_54_real));
  assign _zz_1501 = _zz_5804;
  assign _zz_451 = _zz_5807[35 : 0];
  assign _zz_1502 = _zz_5808;
  assign _zz_452 = _zz_5811[35 : 0];
  assign _zz_454 = 1'b1;
  assign _zz_1503 = _zz_5812;
  assign _zz_1504 = _zz_5820;
  assign _zz_455 = 1'b1;
  assign _zz_1505 = _zz_5828;
  assign _zz_1506 = _zz_5836;
  assign _zz_458 = ($signed(_zz_5844) * $signed(data_mid_2_55_real));
  assign _zz_1507 = _zz_5845;
  assign _zz_456 = _zz_5848[35 : 0];
  assign _zz_1508 = _zz_5849;
  assign _zz_457 = _zz_5852[35 : 0];
  assign _zz_459 = 1'b1;
  assign _zz_1509 = _zz_5853;
  assign _zz_1510 = _zz_5861;
  assign _zz_460 = 1'b1;
  assign _zz_1511 = _zz_5869;
  assign _zz_1512 = _zz_5877;
  assign _zz_463 = ($signed(_zz_5885) * $signed(data_mid_2_60_real));
  assign _zz_1513 = _zz_5886;
  assign _zz_461 = _zz_5889[35 : 0];
  assign _zz_1514 = _zz_5890;
  assign _zz_462 = _zz_5893[35 : 0];
  assign _zz_464 = 1'b1;
  assign _zz_1515 = _zz_5894;
  assign _zz_1516 = _zz_5902;
  assign _zz_465 = 1'b1;
  assign _zz_1517 = _zz_5910;
  assign _zz_1518 = _zz_5918;
  assign _zz_468 = ($signed(_zz_5926) * $signed(data_mid_2_61_real));
  assign _zz_1519 = _zz_5927;
  assign _zz_466 = _zz_5930[35 : 0];
  assign _zz_1520 = _zz_5931;
  assign _zz_467 = _zz_5934[35 : 0];
  assign _zz_469 = 1'b1;
  assign _zz_1521 = _zz_5935;
  assign _zz_1522 = _zz_5943;
  assign _zz_470 = 1'b1;
  assign _zz_1523 = _zz_5951;
  assign _zz_1524 = _zz_5959;
  assign _zz_473 = ($signed(_zz_5967) * $signed(data_mid_2_62_real));
  assign _zz_1525 = _zz_5968;
  assign _zz_471 = _zz_5971[35 : 0];
  assign _zz_1526 = _zz_5972;
  assign _zz_472 = _zz_5975[35 : 0];
  assign _zz_474 = 1'b1;
  assign _zz_1527 = _zz_5976;
  assign _zz_1528 = _zz_5984;
  assign _zz_475 = 1'b1;
  assign _zz_1529 = _zz_5992;
  assign _zz_1530 = _zz_6000;
  assign _zz_478 = ($signed(_zz_6008) * $signed(data_mid_2_63_real));
  assign _zz_1531 = _zz_6009;
  assign _zz_476 = _zz_6012[35 : 0];
  assign _zz_1532 = _zz_6013;
  assign _zz_477 = _zz_6016[35 : 0];
  assign _zz_479 = 1'b1;
  assign _zz_1533 = _zz_6017;
  assign _zz_1534 = _zz_6025;
  assign _zz_480 = 1'b1;
  assign _zz_1535 = _zz_6033;
  assign _zz_1536 = _zz_6041;
  assign _zz_483 = ($signed(_zz_6049) * $signed(data_mid_3_8_real));
  assign _zz_1537 = _zz_6050;
  assign _zz_481 = _zz_6053[35 : 0];
  assign _zz_1538 = _zz_6054;
  assign _zz_482 = _zz_6057[35 : 0];
  assign _zz_484 = 1'b1;
  assign _zz_1539 = _zz_6058;
  assign _zz_1540 = _zz_6066;
  assign _zz_485 = 1'b1;
  assign _zz_1541 = _zz_6074;
  assign _zz_1542 = _zz_6082;
  assign _zz_488 = ($signed(_zz_6090) * $signed(data_mid_3_9_real));
  assign _zz_1543 = _zz_6091;
  assign _zz_486 = _zz_6094[35 : 0];
  assign _zz_1544 = _zz_6095;
  assign _zz_487 = _zz_6098[35 : 0];
  assign _zz_489 = 1'b1;
  assign _zz_1545 = _zz_6099;
  assign _zz_1546 = _zz_6107;
  assign _zz_490 = 1'b1;
  assign _zz_1547 = _zz_6115;
  assign _zz_1548 = _zz_6123;
  assign _zz_493 = ($signed(_zz_6131) * $signed(data_mid_3_10_real));
  assign _zz_1549 = _zz_6132;
  assign _zz_491 = _zz_6135[35 : 0];
  assign _zz_1550 = _zz_6136;
  assign _zz_492 = _zz_6139[35 : 0];
  assign _zz_494 = 1'b1;
  assign _zz_1551 = _zz_6140;
  assign _zz_1552 = _zz_6148;
  assign _zz_495 = 1'b1;
  assign _zz_1553 = _zz_6156;
  assign _zz_1554 = _zz_6164;
  assign _zz_498 = ($signed(_zz_6172) * $signed(data_mid_3_11_real));
  assign _zz_1555 = _zz_6173;
  assign _zz_496 = _zz_6176[35 : 0];
  assign _zz_1556 = _zz_6177;
  assign _zz_497 = _zz_6180[35 : 0];
  assign _zz_499 = 1'b1;
  assign _zz_1557 = _zz_6181;
  assign _zz_1558 = _zz_6189;
  assign _zz_500 = 1'b1;
  assign _zz_1559 = _zz_6197;
  assign _zz_1560 = _zz_6205;
  assign _zz_503 = ($signed(_zz_6213) * $signed(data_mid_3_12_real));
  assign _zz_1561 = _zz_6214;
  assign _zz_501 = _zz_6217[35 : 0];
  assign _zz_1562 = _zz_6218;
  assign _zz_502 = _zz_6221[35 : 0];
  assign _zz_504 = 1'b1;
  assign _zz_1563 = _zz_6222;
  assign _zz_1564 = _zz_6230;
  assign _zz_505 = 1'b1;
  assign _zz_1565 = _zz_6238;
  assign _zz_1566 = _zz_6246;
  assign _zz_508 = ($signed(_zz_6254) * $signed(data_mid_3_13_real));
  assign _zz_1567 = _zz_6255;
  assign _zz_506 = _zz_6258[35 : 0];
  assign _zz_1568 = _zz_6259;
  assign _zz_507 = _zz_6262[35 : 0];
  assign _zz_509 = 1'b1;
  assign _zz_1569 = _zz_6263;
  assign _zz_1570 = _zz_6271;
  assign _zz_510 = 1'b1;
  assign _zz_1571 = _zz_6279;
  assign _zz_1572 = _zz_6287;
  assign _zz_513 = ($signed(_zz_6295) * $signed(data_mid_3_14_real));
  assign _zz_1573 = _zz_6296;
  assign _zz_511 = _zz_6299[35 : 0];
  assign _zz_1574 = _zz_6300;
  assign _zz_512 = _zz_6303[35 : 0];
  assign _zz_514 = 1'b1;
  assign _zz_1575 = _zz_6304;
  assign _zz_1576 = _zz_6312;
  assign _zz_515 = 1'b1;
  assign _zz_1577 = _zz_6320;
  assign _zz_1578 = _zz_6328;
  assign _zz_518 = ($signed(_zz_6336) * $signed(data_mid_3_15_real));
  assign _zz_1579 = _zz_6337;
  assign _zz_516 = _zz_6340[35 : 0];
  assign _zz_1580 = _zz_6341;
  assign _zz_517 = _zz_6344[35 : 0];
  assign _zz_519 = 1'b1;
  assign _zz_1581 = _zz_6345;
  assign _zz_1582 = _zz_6353;
  assign _zz_520 = 1'b1;
  assign _zz_1583 = _zz_6361;
  assign _zz_1584 = _zz_6369;
  assign _zz_523 = ($signed(_zz_6377) * $signed(data_mid_3_24_real));
  assign _zz_1585 = _zz_6378;
  assign _zz_521 = _zz_6381[35 : 0];
  assign _zz_1586 = _zz_6382;
  assign _zz_522 = _zz_6385[35 : 0];
  assign _zz_524 = 1'b1;
  assign _zz_1587 = _zz_6386;
  assign _zz_1588 = _zz_6394;
  assign _zz_525 = 1'b1;
  assign _zz_1589 = _zz_6402;
  assign _zz_1590 = _zz_6410;
  assign _zz_528 = ($signed(_zz_6418) * $signed(data_mid_3_25_real));
  assign _zz_1591 = _zz_6419;
  assign _zz_526 = _zz_6422[35 : 0];
  assign _zz_1592 = _zz_6423;
  assign _zz_527 = _zz_6426[35 : 0];
  assign _zz_529 = 1'b1;
  assign _zz_1593 = _zz_6427;
  assign _zz_1594 = _zz_6435;
  assign _zz_530 = 1'b1;
  assign _zz_1595 = _zz_6443;
  assign _zz_1596 = _zz_6451;
  assign _zz_533 = ($signed(_zz_6459) * $signed(data_mid_3_26_real));
  assign _zz_1597 = _zz_6460;
  assign _zz_531 = _zz_6463[35 : 0];
  assign _zz_1598 = _zz_6464;
  assign _zz_532 = _zz_6467[35 : 0];
  assign _zz_534 = 1'b1;
  assign _zz_1599 = _zz_6468;
  assign _zz_1600 = _zz_6476;
  assign _zz_535 = 1'b1;
  assign _zz_1601 = _zz_6484;
  assign _zz_1602 = _zz_6492;
  assign _zz_538 = ($signed(_zz_6500) * $signed(data_mid_3_27_real));
  assign _zz_1603 = _zz_6501;
  assign _zz_536 = _zz_6504[35 : 0];
  assign _zz_1604 = _zz_6505;
  assign _zz_537 = _zz_6508[35 : 0];
  assign _zz_539 = 1'b1;
  assign _zz_1605 = _zz_6509;
  assign _zz_1606 = _zz_6517;
  assign _zz_540 = 1'b1;
  assign _zz_1607 = _zz_6525;
  assign _zz_1608 = _zz_6533;
  assign _zz_543 = ($signed(_zz_6541) * $signed(data_mid_3_28_real));
  assign _zz_1609 = _zz_6542;
  assign _zz_541 = _zz_6545[35 : 0];
  assign _zz_1610 = _zz_6546;
  assign _zz_542 = _zz_6549[35 : 0];
  assign _zz_544 = 1'b1;
  assign _zz_1611 = _zz_6550;
  assign _zz_1612 = _zz_6558;
  assign _zz_545 = 1'b1;
  assign _zz_1613 = _zz_6566;
  assign _zz_1614 = _zz_6574;
  assign _zz_548 = ($signed(_zz_6582) * $signed(data_mid_3_29_real));
  assign _zz_1615 = _zz_6583;
  assign _zz_546 = _zz_6586[35 : 0];
  assign _zz_1616 = _zz_6587;
  assign _zz_547 = _zz_6590[35 : 0];
  assign _zz_549 = 1'b1;
  assign _zz_1617 = _zz_6591;
  assign _zz_1618 = _zz_6599;
  assign _zz_550 = 1'b1;
  assign _zz_1619 = _zz_6607;
  assign _zz_1620 = _zz_6615;
  assign _zz_553 = ($signed(_zz_6623) * $signed(data_mid_3_30_real));
  assign _zz_1621 = _zz_6624;
  assign _zz_551 = _zz_6627[35 : 0];
  assign _zz_1622 = _zz_6628;
  assign _zz_552 = _zz_6631[35 : 0];
  assign _zz_554 = 1'b1;
  assign _zz_1623 = _zz_6632;
  assign _zz_1624 = _zz_6640;
  assign _zz_555 = 1'b1;
  assign _zz_1625 = _zz_6648;
  assign _zz_1626 = _zz_6656;
  assign _zz_558 = ($signed(_zz_6664) * $signed(data_mid_3_31_real));
  assign _zz_1627 = _zz_6665;
  assign _zz_556 = _zz_6668[35 : 0];
  assign _zz_1628 = _zz_6669;
  assign _zz_557 = _zz_6672[35 : 0];
  assign _zz_559 = 1'b1;
  assign _zz_1629 = _zz_6673;
  assign _zz_1630 = _zz_6681;
  assign _zz_560 = 1'b1;
  assign _zz_1631 = _zz_6689;
  assign _zz_1632 = _zz_6697;
  assign _zz_563 = ($signed(_zz_6705) * $signed(data_mid_3_40_real));
  assign _zz_1633 = _zz_6706;
  assign _zz_561 = _zz_6709[35 : 0];
  assign _zz_1634 = _zz_6710;
  assign _zz_562 = _zz_6713[35 : 0];
  assign _zz_564 = 1'b1;
  assign _zz_1635 = _zz_6714;
  assign _zz_1636 = _zz_6722;
  assign _zz_565 = 1'b1;
  assign _zz_1637 = _zz_6730;
  assign _zz_1638 = _zz_6738;
  assign _zz_568 = ($signed(_zz_6746) * $signed(data_mid_3_41_real));
  assign _zz_1639 = _zz_6747;
  assign _zz_566 = _zz_6750[35 : 0];
  assign _zz_1640 = _zz_6751;
  assign _zz_567 = _zz_6754[35 : 0];
  assign _zz_569 = 1'b1;
  assign _zz_1641 = _zz_6755;
  assign _zz_1642 = _zz_6763;
  assign _zz_570 = 1'b1;
  assign _zz_1643 = _zz_6771;
  assign _zz_1644 = _zz_6779;
  assign _zz_573 = ($signed(_zz_6787) * $signed(data_mid_3_42_real));
  assign _zz_1645 = _zz_6788;
  assign _zz_571 = _zz_6791[35 : 0];
  assign _zz_1646 = _zz_6792;
  assign _zz_572 = _zz_6795[35 : 0];
  assign _zz_574 = 1'b1;
  assign _zz_1647 = _zz_6796;
  assign _zz_1648 = _zz_6804;
  assign _zz_575 = 1'b1;
  assign _zz_1649 = _zz_6812;
  assign _zz_1650 = _zz_6820;
  assign _zz_578 = ($signed(_zz_6828) * $signed(data_mid_3_43_real));
  assign _zz_1651 = _zz_6829;
  assign _zz_576 = _zz_6832[35 : 0];
  assign _zz_1652 = _zz_6833;
  assign _zz_577 = _zz_6836[35 : 0];
  assign _zz_579 = 1'b1;
  assign _zz_1653 = _zz_6837;
  assign _zz_1654 = _zz_6845;
  assign _zz_580 = 1'b1;
  assign _zz_1655 = _zz_6853;
  assign _zz_1656 = _zz_6861;
  assign _zz_583 = ($signed(_zz_6869) * $signed(data_mid_3_44_real));
  assign _zz_1657 = _zz_6870;
  assign _zz_581 = _zz_6873[35 : 0];
  assign _zz_1658 = _zz_6874;
  assign _zz_582 = _zz_6877[35 : 0];
  assign _zz_584 = 1'b1;
  assign _zz_1659 = _zz_6878;
  assign _zz_1660 = _zz_6886;
  assign _zz_585 = 1'b1;
  assign _zz_1661 = _zz_6894;
  assign _zz_1662 = _zz_6902;
  assign _zz_588 = ($signed(_zz_6910) * $signed(data_mid_3_45_real));
  assign _zz_1663 = _zz_6911;
  assign _zz_586 = _zz_6914[35 : 0];
  assign _zz_1664 = _zz_6915;
  assign _zz_587 = _zz_6918[35 : 0];
  assign _zz_589 = 1'b1;
  assign _zz_1665 = _zz_6919;
  assign _zz_1666 = _zz_6927;
  assign _zz_590 = 1'b1;
  assign _zz_1667 = _zz_6935;
  assign _zz_1668 = _zz_6943;
  assign _zz_593 = ($signed(_zz_6951) * $signed(data_mid_3_46_real));
  assign _zz_1669 = _zz_6952;
  assign _zz_591 = _zz_6955[35 : 0];
  assign _zz_1670 = _zz_6956;
  assign _zz_592 = _zz_6959[35 : 0];
  assign _zz_594 = 1'b1;
  assign _zz_1671 = _zz_6960;
  assign _zz_1672 = _zz_6968;
  assign _zz_595 = 1'b1;
  assign _zz_1673 = _zz_6976;
  assign _zz_1674 = _zz_6984;
  assign _zz_598 = ($signed(_zz_6992) * $signed(data_mid_3_47_real));
  assign _zz_1675 = _zz_6993;
  assign _zz_596 = _zz_6996[35 : 0];
  assign _zz_1676 = _zz_6997;
  assign _zz_597 = _zz_7000[35 : 0];
  assign _zz_599 = 1'b1;
  assign _zz_1677 = _zz_7001;
  assign _zz_1678 = _zz_7009;
  assign _zz_600 = 1'b1;
  assign _zz_1679 = _zz_7017;
  assign _zz_1680 = _zz_7025;
  assign _zz_603 = ($signed(_zz_7033) * $signed(data_mid_3_56_real));
  assign _zz_1681 = _zz_7034;
  assign _zz_601 = _zz_7037[35 : 0];
  assign _zz_1682 = _zz_7038;
  assign _zz_602 = _zz_7041[35 : 0];
  assign _zz_604 = 1'b1;
  assign _zz_1683 = _zz_7042;
  assign _zz_1684 = _zz_7050;
  assign _zz_605 = 1'b1;
  assign _zz_1685 = _zz_7058;
  assign _zz_1686 = _zz_7066;
  assign _zz_608 = ($signed(_zz_7074) * $signed(data_mid_3_57_real));
  assign _zz_1687 = _zz_7075;
  assign _zz_606 = _zz_7078[35 : 0];
  assign _zz_1688 = _zz_7079;
  assign _zz_607 = _zz_7082[35 : 0];
  assign _zz_609 = 1'b1;
  assign _zz_1689 = _zz_7083;
  assign _zz_1690 = _zz_7091;
  assign _zz_610 = 1'b1;
  assign _zz_1691 = _zz_7099;
  assign _zz_1692 = _zz_7107;
  assign _zz_613 = ($signed(_zz_7115) * $signed(data_mid_3_58_real));
  assign _zz_1693 = _zz_7116;
  assign _zz_611 = _zz_7119[35 : 0];
  assign _zz_1694 = _zz_7120;
  assign _zz_612 = _zz_7123[35 : 0];
  assign _zz_614 = 1'b1;
  assign _zz_1695 = _zz_7124;
  assign _zz_1696 = _zz_7132;
  assign _zz_615 = 1'b1;
  assign _zz_1697 = _zz_7140;
  assign _zz_1698 = _zz_7148;
  assign _zz_618 = ($signed(_zz_7156) * $signed(data_mid_3_59_real));
  assign _zz_1699 = _zz_7157;
  assign _zz_616 = _zz_7160[35 : 0];
  assign _zz_1700 = _zz_7161;
  assign _zz_617 = _zz_7164[35 : 0];
  assign _zz_619 = 1'b1;
  assign _zz_1701 = _zz_7165;
  assign _zz_1702 = _zz_7173;
  assign _zz_620 = 1'b1;
  assign _zz_1703 = _zz_7181;
  assign _zz_1704 = _zz_7189;
  assign _zz_623 = ($signed(_zz_7197) * $signed(data_mid_3_60_real));
  assign _zz_1705 = _zz_7198;
  assign _zz_621 = _zz_7201[35 : 0];
  assign _zz_1706 = _zz_7202;
  assign _zz_622 = _zz_7205[35 : 0];
  assign _zz_624 = 1'b1;
  assign _zz_1707 = _zz_7206;
  assign _zz_1708 = _zz_7214;
  assign _zz_625 = 1'b1;
  assign _zz_1709 = _zz_7222;
  assign _zz_1710 = _zz_7230;
  assign _zz_628 = ($signed(_zz_7238) * $signed(data_mid_3_61_real));
  assign _zz_1711 = _zz_7239;
  assign _zz_626 = _zz_7242[35 : 0];
  assign _zz_1712 = _zz_7243;
  assign _zz_627 = _zz_7246[35 : 0];
  assign _zz_629 = 1'b1;
  assign _zz_1713 = _zz_7247;
  assign _zz_1714 = _zz_7255;
  assign _zz_630 = 1'b1;
  assign _zz_1715 = _zz_7263;
  assign _zz_1716 = _zz_7271;
  assign _zz_633 = ($signed(_zz_7279) * $signed(data_mid_3_62_real));
  assign _zz_1717 = _zz_7280;
  assign _zz_631 = _zz_7283[35 : 0];
  assign _zz_1718 = _zz_7284;
  assign _zz_632 = _zz_7287[35 : 0];
  assign _zz_634 = 1'b1;
  assign _zz_1719 = _zz_7288;
  assign _zz_1720 = _zz_7296;
  assign _zz_635 = 1'b1;
  assign _zz_1721 = _zz_7304;
  assign _zz_1722 = _zz_7312;
  assign _zz_638 = ($signed(_zz_7320) * $signed(data_mid_3_63_real));
  assign _zz_1723 = _zz_7321;
  assign _zz_636 = _zz_7324[35 : 0];
  assign _zz_1724 = _zz_7325;
  assign _zz_637 = _zz_7328[35 : 0];
  assign _zz_639 = 1'b1;
  assign _zz_1725 = _zz_7329;
  assign _zz_1726 = _zz_7337;
  assign _zz_640 = 1'b1;
  assign _zz_1727 = _zz_7345;
  assign _zz_1728 = _zz_7353;
  assign _zz_643 = ($signed(_zz_7361) * $signed(data_mid_4_16_real));
  assign _zz_1729 = _zz_7362;
  assign _zz_641 = _zz_7365[35 : 0];
  assign _zz_1730 = _zz_7366;
  assign _zz_642 = _zz_7369[35 : 0];
  assign _zz_644 = 1'b1;
  assign _zz_1731 = _zz_7370;
  assign _zz_1732 = _zz_7378;
  assign _zz_645 = 1'b1;
  assign _zz_1733 = _zz_7386;
  assign _zz_1734 = _zz_7394;
  assign _zz_648 = ($signed(_zz_7402) * $signed(data_mid_4_17_real));
  assign _zz_1735 = _zz_7403;
  assign _zz_646 = _zz_7406[35 : 0];
  assign _zz_1736 = _zz_7407;
  assign _zz_647 = _zz_7410[35 : 0];
  assign _zz_649 = 1'b1;
  assign _zz_1737 = _zz_7411;
  assign _zz_1738 = _zz_7419;
  assign _zz_650 = 1'b1;
  assign _zz_1739 = _zz_7427;
  assign _zz_1740 = _zz_7435;
  assign _zz_653 = ($signed(_zz_7443) * $signed(data_mid_4_18_real));
  assign _zz_1741 = _zz_7444;
  assign _zz_651 = _zz_7447[35 : 0];
  assign _zz_1742 = _zz_7448;
  assign _zz_652 = _zz_7451[35 : 0];
  assign _zz_654 = 1'b1;
  assign _zz_1743 = _zz_7452;
  assign _zz_1744 = _zz_7460;
  assign _zz_655 = 1'b1;
  assign _zz_1745 = _zz_7468;
  assign _zz_1746 = _zz_7476;
  assign _zz_658 = ($signed(_zz_7484) * $signed(data_mid_4_19_real));
  assign _zz_1747 = _zz_7485;
  assign _zz_656 = _zz_7488[35 : 0];
  assign _zz_1748 = _zz_7489;
  assign _zz_657 = _zz_7492[35 : 0];
  assign _zz_659 = 1'b1;
  assign _zz_1749 = _zz_7493;
  assign _zz_1750 = _zz_7501;
  assign _zz_660 = 1'b1;
  assign _zz_1751 = _zz_7509;
  assign _zz_1752 = _zz_7517;
  assign _zz_663 = ($signed(_zz_7525) * $signed(data_mid_4_20_real));
  assign _zz_1753 = _zz_7526;
  assign _zz_661 = _zz_7529[35 : 0];
  assign _zz_1754 = _zz_7530;
  assign _zz_662 = _zz_7533[35 : 0];
  assign _zz_664 = 1'b1;
  assign _zz_1755 = _zz_7534;
  assign _zz_1756 = _zz_7542;
  assign _zz_665 = 1'b1;
  assign _zz_1757 = _zz_7550;
  assign _zz_1758 = _zz_7558;
  assign _zz_668 = ($signed(_zz_7566) * $signed(data_mid_4_21_real));
  assign _zz_1759 = _zz_7567;
  assign _zz_666 = _zz_7570[35 : 0];
  assign _zz_1760 = _zz_7571;
  assign _zz_667 = _zz_7574[35 : 0];
  assign _zz_669 = 1'b1;
  assign _zz_1761 = _zz_7575;
  assign _zz_1762 = _zz_7583;
  assign _zz_670 = 1'b1;
  assign _zz_1763 = _zz_7591;
  assign _zz_1764 = _zz_7599;
  assign _zz_673 = ($signed(_zz_7607) * $signed(data_mid_4_22_real));
  assign _zz_1765 = _zz_7608;
  assign _zz_671 = _zz_7611[35 : 0];
  assign _zz_1766 = _zz_7612;
  assign _zz_672 = _zz_7615[35 : 0];
  assign _zz_674 = 1'b1;
  assign _zz_1767 = _zz_7616;
  assign _zz_1768 = _zz_7624;
  assign _zz_675 = 1'b1;
  assign _zz_1769 = _zz_7632;
  assign _zz_1770 = _zz_7640;
  assign _zz_678 = ($signed(_zz_7648) * $signed(data_mid_4_23_real));
  assign _zz_1771 = _zz_7649;
  assign _zz_676 = _zz_7652[35 : 0];
  assign _zz_1772 = _zz_7653;
  assign _zz_677 = _zz_7656[35 : 0];
  assign _zz_679 = 1'b1;
  assign _zz_1773 = _zz_7657;
  assign _zz_1774 = _zz_7665;
  assign _zz_680 = 1'b1;
  assign _zz_1775 = _zz_7673;
  assign _zz_1776 = _zz_7681;
  assign _zz_683 = ($signed(_zz_7689) * $signed(data_mid_4_24_real));
  assign _zz_1777 = _zz_7690;
  assign _zz_681 = _zz_7693[35 : 0];
  assign _zz_1778 = _zz_7694;
  assign _zz_682 = _zz_7697[35 : 0];
  assign _zz_684 = 1'b1;
  assign _zz_1779 = _zz_7698;
  assign _zz_1780 = _zz_7706;
  assign _zz_685 = 1'b1;
  assign _zz_1781 = _zz_7714;
  assign _zz_1782 = _zz_7722;
  assign _zz_688 = ($signed(_zz_7730) * $signed(data_mid_4_25_real));
  assign _zz_1783 = _zz_7731;
  assign _zz_686 = _zz_7734[35 : 0];
  assign _zz_1784 = _zz_7735;
  assign _zz_687 = _zz_7738[35 : 0];
  assign _zz_689 = 1'b1;
  assign _zz_1785 = _zz_7739;
  assign _zz_1786 = _zz_7747;
  assign _zz_690 = 1'b1;
  assign _zz_1787 = _zz_7755;
  assign _zz_1788 = _zz_7763;
  assign _zz_693 = ($signed(_zz_7771) * $signed(data_mid_4_26_real));
  assign _zz_1789 = _zz_7772;
  assign _zz_691 = _zz_7775[35 : 0];
  assign _zz_1790 = _zz_7776;
  assign _zz_692 = _zz_7779[35 : 0];
  assign _zz_694 = 1'b1;
  assign _zz_1791 = _zz_7780;
  assign _zz_1792 = _zz_7788;
  assign _zz_695 = 1'b1;
  assign _zz_1793 = _zz_7796;
  assign _zz_1794 = _zz_7804;
  assign _zz_698 = ($signed(_zz_7812) * $signed(data_mid_4_27_real));
  assign _zz_1795 = _zz_7813;
  assign _zz_696 = _zz_7816[35 : 0];
  assign _zz_1796 = _zz_7817;
  assign _zz_697 = _zz_7820[35 : 0];
  assign _zz_699 = 1'b1;
  assign _zz_1797 = _zz_7821;
  assign _zz_1798 = _zz_7829;
  assign _zz_700 = 1'b1;
  assign _zz_1799 = _zz_7837;
  assign _zz_1800 = _zz_7845;
  assign _zz_703 = ($signed(_zz_7853) * $signed(data_mid_4_28_real));
  assign _zz_1801 = _zz_7854;
  assign _zz_701 = _zz_7857[35 : 0];
  assign _zz_1802 = _zz_7858;
  assign _zz_702 = _zz_7861[35 : 0];
  assign _zz_704 = 1'b1;
  assign _zz_1803 = _zz_7862;
  assign _zz_1804 = _zz_7870;
  assign _zz_705 = 1'b1;
  assign _zz_1805 = _zz_7878;
  assign _zz_1806 = _zz_7886;
  assign _zz_708 = ($signed(_zz_7894) * $signed(data_mid_4_29_real));
  assign _zz_1807 = _zz_7895;
  assign _zz_706 = _zz_7898[35 : 0];
  assign _zz_1808 = _zz_7899;
  assign _zz_707 = _zz_7902[35 : 0];
  assign _zz_709 = 1'b1;
  assign _zz_1809 = _zz_7903;
  assign _zz_1810 = _zz_7911;
  assign _zz_710 = 1'b1;
  assign _zz_1811 = _zz_7919;
  assign _zz_1812 = _zz_7927;
  assign _zz_713 = ($signed(_zz_7935) * $signed(data_mid_4_30_real));
  assign _zz_1813 = _zz_7936;
  assign _zz_711 = _zz_7939[35 : 0];
  assign _zz_1814 = _zz_7940;
  assign _zz_712 = _zz_7943[35 : 0];
  assign _zz_714 = 1'b1;
  assign _zz_1815 = _zz_7944;
  assign _zz_1816 = _zz_7952;
  assign _zz_715 = 1'b1;
  assign _zz_1817 = _zz_7960;
  assign _zz_1818 = _zz_7968;
  assign _zz_718 = ($signed(_zz_7976) * $signed(data_mid_4_31_real));
  assign _zz_1819 = _zz_7977;
  assign _zz_716 = _zz_7980[35 : 0];
  assign _zz_1820 = _zz_7981;
  assign _zz_717 = _zz_7984[35 : 0];
  assign _zz_719 = 1'b1;
  assign _zz_1821 = _zz_7985;
  assign _zz_1822 = _zz_7993;
  assign _zz_720 = 1'b1;
  assign _zz_1823 = _zz_8001;
  assign _zz_1824 = _zz_8009;
  assign _zz_723 = ($signed(_zz_8017) * $signed(data_mid_4_48_real));
  assign _zz_1825 = _zz_8018;
  assign _zz_721 = _zz_8021[35 : 0];
  assign _zz_1826 = _zz_8022;
  assign _zz_722 = _zz_8025[35 : 0];
  assign _zz_724 = 1'b1;
  assign _zz_1827 = _zz_8026;
  assign _zz_1828 = _zz_8034;
  assign _zz_725 = 1'b1;
  assign _zz_1829 = _zz_8042;
  assign _zz_1830 = _zz_8050;
  assign _zz_728 = ($signed(_zz_8058) * $signed(data_mid_4_49_real));
  assign _zz_1831 = _zz_8059;
  assign _zz_726 = _zz_8062[35 : 0];
  assign _zz_1832 = _zz_8063;
  assign _zz_727 = _zz_8066[35 : 0];
  assign _zz_729 = 1'b1;
  assign _zz_1833 = _zz_8067;
  assign _zz_1834 = _zz_8075;
  assign _zz_730 = 1'b1;
  assign _zz_1835 = _zz_8083;
  assign _zz_1836 = _zz_8091;
  assign _zz_733 = ($signed(_zz_8099) * $signed(data_mid_4_50_real));
  assign _zz_1837 = _zz_8100;
  assign _zz_731 = _zz_8103[35 : 0];
  assign _zz_1838 = _zz_8104;
  assign _zz_732 = _zz_8107[35 : 0];
  assign _zz_734 = 1'b1;
  assign _zz_1839 = _zz_8108;
  assign _zz_1840 = _zz_8116;
  assign _zz_735 = 1'b1;
  assign _zz_1841 = _zz_8124;
  assign _zz_1842 = _zz_8132;
  assign _zz_738 = ($signed(_zz_8140) * $signed(data_mid_4_51_real));
  assign _zz_1843 = _zz_8141;
  assign _zz_736 = _zz_8144[35 : 0];
  assign _zz_1844 = _zz_8145;
  assign _zz_737 = _zz_8148[35 : 0];
  assign _zz_739 = 1'b1;
  assign _zz_1845 = _zz_8149;
  assign _zz_1846 = _zz_8157;
  assign _zz_740 = 1'b1;
  assign _zz_1847 = _zz_8165;
  assign _zz_1848 = _zz_8173;
  assign _zz_743 = ($signed(_zz_8181) * $signed(data_mid_4_52_real));
  assign _zz_1849 = _zz_8182;
  assign _zz_741 = _zz_8185[35 : 0];
  assign _zz_1850 = _zz_8186;
  assign _zz_742 = _zz_8189[35 : 0];
  assign _zz_744 = 1'b1;
  assign _zz_1851 = _zz_8190;
  assign _zz_1852 = _zz_8198;
  assign _zz_745 = 1'b1;
  assign _zz_1853 = _zz_8206;
  assign _zz_1854 = _zz_8214;
  assign _zz_748 = ($signed(_zz_8222) * $signed(data_mid_4_53_real));
  assign _zz_1855 = _zz_8223;
  assign _zz_746 = _zz_8226[35 : 0];
  assign _zz_1856 = _zz_8227;
  assign _zz_747 = _zz_8230[35 : 0];
  assign _zz_749 = 1'b1;
  assign _zz_1857 = _zz_8231;
  assign _zz_1858 = _zz_8239;
  assign _zz_750 = 1'b1;
  assign _zz_1859 = _zz_8247;
  assign _zz_1860 = _zz_8255;
  assign _zz_753 = ($signed(_zz_8263) * $signed(data_mid_4_54_real));
  assign _zz_1861 = _zz_8264;
  assign _zz_751 = _zz_8267[35 : 0];
  assign _zz_1862 = _zz_8268;
  assign _zz_752 = _zz_8271[35 : 0];
  assign _zz_754 = 1'b1;
  assign _zz_1863 = _zz_8272;
  assign _zz_1864 = _zz_8280;
  assign _zz_755 = 1'b1;
  assign _zz_1865 = _zz_8288;
  assign _zz_1866 = _zz_8296;
  assign _zz_758 = ($signed(_zz_8304) * $signed(data_mid_4_55_real));
  assign _zz_1867 = _zz_8305;
  assign _zz_756 = _zz_8308[35 : 0];
  assign _zz_1868 = _zz_8309;
  assign _zz_757 = _zz_8312[35 : 0];
  assign _zz_759 = 1'b1;
  assign _zz_1869 = _zz_8313;
  assign _zz_1870 = _zz_8321;
  assign _zz_760 = 1'b1;
  assign _zz_1871 = _zz_8329;
  assign _zz_1872 = _zz_8337;
  assign _zz_763 = ($signed(_zz_8345) * $signed(data_mid_4_56_real));
  assign _zz_1873 = _zz_8346;
  assign _zz_761 = _zz_8349[35 : 0];
  assign _zz_1874 = _zz_8350;
  assign _zz_762 = _zz_8353[35 : 0];
  assign _zz_764 = 1'b1;
  assign _zz_1875 = _zz_8354;
  assign _zz_1876 = _zz_8362;
  assign _zz_765 = 1'b1;
  assign _zz_1877 = _zz_8370;
  assign _zz_1878 = _zz_8378;
  assign _zz_768 = ($signed(_zz_8386) * $signed(data_mid_4_57_real));
  assign _zz_1879 = _zz_8387;
  assign _zz_766 = _zz_8390[35 : 0];
  assign _zz_1880 = _zz_8391;
  assign _zz_767 = _zz_8394[35 : 0];
  assign _zz_769 = 1'b1;
  assign _zz_1881 = _zz_8395;
  assign _zz_1882 = _zz_8403;
  assign _zz_770 = 1'b1;
  assign _zz_1883 = _zz_8411;
  assign _zz_1884 = _zz_8419;
  assign _zz_773 = ($signed(_zz_8427) * $signed(data_mid_4_58_real));
  assign _zz_1885 = _zz_8428;
  assign _zz_771 = _zz_8431[35 : 0];
  assign _zz_1886 = _zz_8432;
  assign _zz_772 = _zz_8435[35 : 0];
  assign _zz_774 = 1'b1;
  assign _zz_1887 = _zz_8436;
  assign _zz_1888 = _zz_8444;
  assign _zz_775 = 1'b1;
  assign _zz_1889 = _zz_8452;
  assign _zz_1890 = _zz_8460;
  assign _zz_778 = ($signed(_zz_8468) * $signed(data_mid_4_59_real));
  assign _zz_1891 = _zz_8469;
  assign _zz_776 = _zz_8472[35 : 0];
  assign _zz_1892 = _zz_8473;
  assign _zz_777 = _zz_8476[35 : 0];
  assign _zz_779 = 1'b1;
  assign _zz_1893 = _zz_8477;
  assign _zz_1894 = _zz_8485;
  assign _zz_780 = 1'b1;
  assign _zz_1895 = _zz_8493;
  assign _zz_1896 = _zz_8501;
  assign _zz_783 = ($signed(_zz_8509) * $signed(data_mid_4_60_real));
  assign _zz_1897 = _zz_8510;
  assign _zz_781 = _zz_8513[35 : 0];
  assign _zz_1898 = _zz_8514;
  assign _zz_782 = _zz_8517[35 : 0];
  assign _zz_784 = 1'b1;
  assign _zz_1899 = _zz_8518;
  assign _zz_1900 = _zz_8526;
  assign _zz_785 = 1'b1;
  assign _zz_1901 = _zz_8534;
  assign _zz_1902 = _zz_8542;
  assign _zz_788 = ($signed(_zz_8550) * $signed(data_mid_4_61_real));
  assign _zz_1903 = _zz_8551;
  assign _zz_786 = _zz_8554[35 : 0];
  assign _zz_1904 = _zz_8555;
  assign _zz_787 = _zz_8558[35 : 0];
  assign _zz_789 = 1'b1;
  assign _zz_1905 = _zz_8559;
  assign _zz_1906 = _zz_8567;
  assign _zz_790 = 1'b1;
  assign _zz_1907 = _zz_8575;
  assign _zz_1908 = _zz_8583;
  assign _zz_793 = ($signed(_zz_8591) * $signed(data_mid_4_62_real));
  assign _zz_1909 = _zz_8592;
  assign _zz_791 = _zz_8595[35 : 0];
  assign _zz_1910 = _zz_8596;
  assign _zz_792 = _zz_8599[35 : 0];
  assign _zz_794 = 1'b1;
  assign _zz_1911 = _zz_8600;
  assign _zz_1912 = _zz_8608;
  assign _zz_795 = 1'b1;
  assign _zz_1913 = _zz_8616;
  assign _zz_1914 = _zz_8624;
  assign _zz_798 = ($signed(_zz_8632) * $signed(data_mid_4_63_real));
  assign _zz_1915 = _zz_8633;
  assign _zz_796 = _zz_8636[35 : 0];
  assign _zz_1916 = _zz_8637;
  assign _zz_797 = _zz_8640[35 : 0];
  assign _zz_799 = 1'b1;
  assign _zz_1917 = _zz_8641;
  assign _zz_1918 = _zz_8649;
  assign _zz_800 = 1'b1;
  assign _zz_1919 = _zz_8657;
  assign _zz_1920 = _zz_8665;
  assign _zz_803 = ($signed(_zz_8673) * $signed(data_mid_5_32_real));
  assign _zz_1921 = _zz_8674;
  assign _zz_801 = _zz_8677[35 : 0];
  assign _zz_1922 = _zz_8678;
  assign _zz_802 = _zz_8681[35 : 0];
  assign _zz_804 = 1'b1;
  assign _zz_1923 = _zz_8682;
  assign _zz_1924 = _zz_8690;
  assign _zz_805 = 1'b1;
  assign _zz_1925 = _zz_8698;
  assign _zz_1926 = _zz_8706;
  assign _zz_808 = ($signed(_zz_8714) * $signed(data_mid_5_33_real));
  assign _zz_1927 = _zz_8715;
  assign _zz_806 = _zz_8718[35 : 0];
  assign _zz_1928 = _zz_8719;
  assign _zz_807 = _zz_8722[35 : 0];
  assign _zz_809 = 1'b1;
  assign _zz_1929 = _zz_8723;
  assign _zz_1930 = _zz_8731;
  assign _zz_810 = 1'b1;
  assign _zz_1931 = _zz_8739;
  assign _zz_1932 = _zz_8747;
  assign _zz_813 = ($signed(_zz_8755) * $signed(data_mid_5_34_real));
  assign _zz_1933 = _zz_8756;
  assign _zz_811 = _zz_8759[35 : 0];
  assign _zz_1934 = _zz_8760;
  assign _zz_812 = _zz_8763[35 : 0];
  assign _zz_814 = 1'b1;
  assign _zz_1935 = _zz_8764;
  assign _zz_1936 = _zz_8772;
  assign _zz_815 = 1'b1;
  assign _zz_1937 = _zz_8780;
  assign _zz_1938 = _zz_8788;
  assign _zz_818 = ($signed(_zz_8796) * $signed(data_mid_5_35_real));
  assign _zz_1939 = _zz_8797;
  assign _zz_816 = _zz_8800[35 : 0];
  assign _zz_1940 = _zz_8801;
  assign _zz_817 = _zz_8804[35 : 0];
  assign _zz_819 = 1'b1;
  assign _zz_1941 = _zz_8805;
  assign _zz_1942 = _zz_8813;
  assign _zz_820 = 1'b1;
  assign _zz_1943 = _zz_8821;
  assign _zz_1944 = _zz_8829;
  assign _zz_823 = ($signed(_zz_8837) * $signed(data_mid_5_36_real));
  assign _zz_1945 = _zz_8838;
  assign _zz_821 = _zz_8841[35 : 0];
  assign _zz_1946 = _zz_8842;
  assign _zz_822 = _zz_8845[35 : 0];
  assign _zz_824 = 1'b1;
  assign _zz_1947 = _zz_8846;
  assign _zz_1948 = _zz_8854;
  assign _zz_825 = 1'b1;
  assign _zz_1949 = _zz_8862;
  assign _zz_1950 = _zz_8870;
  assign _zz_828 = ($signed(_zz_8878) * $signed(data_mid_5_37_real));
  assign _zz_1951 = _zz_8879;
  assign _zz_826 = _zz_8882[35 : 0];
  assign _zz_1952 = _zz_8883;
  assign _zz_827 = _zz_8886[35 : 0];
  assign _zz_829 = 1'b1;
  assign _zz_1953 = _zz_8887;
  assign _zz_1954 = _zz_8895;
  assign _zz_830 = 1'b1;
  assign _zz_1955 = _zz_8903;
  assign _zz_1956 = _zz_8911;
  assign _zz_833 = ($signed(_zz_8919) * $signed(data_mid_5_38_real));
  assign _zz_1957 = _zz_8920;
  assign _zz_831 = _zz_8923[35 : 0];
  assign _zz_1958 = _zz_8924;
  assign _zz_832 = _zz_8927[35 : 0];
  assign _zz_834 = 1'b1;
  assign _zz_1959 = _zz_8928;
  assign _zz_1960 = _zz_8936;
  assign _zz_835 = 1'b1;
  assign _zz_1961 = _zz_8944;
  assign _zz_1962 = _zz_8952;
  assign _zz_838 = ($signed(_zz_8960) * $signed(data_mid_5_39_real));
  assign _zz_1963 = _zz_8961;
  assign _zz_836 = _zz_8964[35 : 0];
  assign _zz_1964 = _zz_8965;
  assign _zz_837 = _zz_8968[35 : 0];
  assign _zz_839 = 1'b1;
  assign _zz_1965 = _zz_8969;
  assign _zz_1966 = _zz_8977;
  assign _zz_840 = 1'b1;
  assign _zz_1967 = _zz_8985;
  assign _zz_1968 = _zz_8993;
  assign _zz_843 = ($signed(_zz_9001) * $signed(data_mid_5_40_real));
  assign _zz_1969 = _zz_9002;
  assign _zz_841 = _zz_9005[35 : 0];
  assign _zz_1970 = _zz_9006;
  assign _zz_842 = _zz_9009[35 : 0];
  assign _zz_844 = 1'b1;
  assign _zz_1971 = _zz_9010;
  assign _zz_1972 = _zz_9018;
  assign _zz_845 = 1'b1;
  assign _zz_1973 = _zz_9026;
  assign _zz_1974 = _zz_9034;
  assign _zz_848 = ($signed(_zz_9042) * $signed(data_mid_5_41_real));
  assign _zz_1975 = _zz_9043;
  assign _zz_846 = _zz_9046[35 : 0];
  assign _zz_1976 = _zz_9047;
  assign _zz_847 = _zz_9050[35 : 0];
  assign _zz_849 = 1'b1;
  assign _zz_1977 = _zz_9051;
  assign _zz_1978 = _zz_9059;
  assign _zz_850 = 1'b1;
  assign _zz_1979 = _zz_9067;
  assign _zz_1980 = _zz_9075;
  assign _zz_853 = ($signed(_zz_9083) * $signed(data_mid_5_42_real));
  assign _zz_1981 = _zz_9084;
  assign _zz_851 = _zz_9087[35 : 0];
  assign _zz_1982 = _zz_9088;
  assign _zz_852 = _zz_9091[35 : 0];
  assign _zz_854 = 1'b1;
  assign _zz_1983 = _zz_9092;
  assign _zz_1984 = _zz_9100;
  assign _zz_855 = 1'b1;
  assign _zz_1985 = _zz_9108;
  assign _zz_1986 = _zz_9116;
  assign _zz_858 = ($signed(_zz_9124) * $signed(data_mid_5_43_real));
  assign _zz_1987 = _zz_9125;
  assign _zz_856 = _zz_9128[35 : 0];
  assign _zz_1988 = _zz_9129;
  assign _zz_857 = _zz_9132[35 : 0];
  assign _zz_859 = 1'b1;
  assign _zz_1989 = _zz_9133;
  assign _zz_1990 = _zz_9141;
  assign _zz_860 = 1'b1;
  assign _zz_1991 = _zz_9149;
  assign _zz_1992 = _zz_9157;
  assign _zz_863 = ($signed(_zz_9165) * $signed(data_mid_5_44_real));
  assign _zz_1993 = _zz_9166;
  assign _zz_861 = _zz_9169[35 : 0];
  assign _zz_1994 = _zz_9170;
  assign _zz_862 = _zz_9173[35 : 0];
  assign _zz_864 = 1'b1;
  assign _zz_1995 = _zz_9174;
  assign _zz_1996 = _zz_9182;
  assign _zz_865 = 1'b1;
  assign _zz_1997 = _zz_9190;
  assign _zz_1998 = _zz_9198;
  assign _zz_868 = ($signed(_zz_9206) * $signed(data_mid_5_45_real));
  assign _zz_1999 = _zz_9207;
  assign _zz_866 = _zz_9210[35 : 0];
  assign _zz_2000 = _zz_9211;
  assign _zz_867 = _zz_9214[35 : 0];
  assign _zz_869 = 1'b1;
  assign _zz_2001 = _zz_9215;
  assign _zz_2002 = _zz_9223;
  assign _zz_870 = 1'b1;
  assign _zz_2003 = _zz_9231;
  assign _zz_2004 = _zz_9239;
  assign _zz_873 = ($signed(_zz_9247) * $signed(data_mid_5_46_real));
  assign _zz_2005 = _zz_9248;
  assign _zz_871 = _zz_9251[35 : 0];
  assign _zz_2006 = _zz_9252;
  assign _zz_872 = _zz_9255[35 : 0];
  assign _zz_874 = 1'b1;
  assign _zz_2007 = _zz_9256;
  assign _zz_2008 = _zz_9264;
  assign _zz_875 = 1'b1;
  assign _zz_2009 = _zz_9272;
  assign _zz_2010 = _zz_9280;
  assign _zz_878 = ($signed(_zz_9288) * $signed(data_mid_5_47_real));
  assign _zz_2011 = _zz_9289;
  assign _zz_876 = _zz_9292[35 : 0];
  assign _zz_2012 = _zz_9293;
  assign _zz_877 = _zz_9296[35 : 0];
  assign _zz_879 = 1'b1;
  assign _zz_2013 = _zz_9297;
  assign _zz_2014 = _zz_9305;
  assign _zz_880 = 1'b1;
  assign _zz_2015 = _zz_9313;
  assign _zz_2016 = _zz_9321;
  assign _zz_883 = ($signed(_zz_9329) * $signed(data_mid_5_48_real));
  assign _zz_2017 = _zz_9330;
  assign _zz_881 = _zz_9333[35 : 0];
  assign _zz_2018 = _zz_9334;
  assign _zz_882 = _zz_9337[35 : 0];
  assign _zz_884 = 1'b1;
  assign _zz_2019 = _zz_9338;
  assign _zz_2020 = _zz_9346;
  assign _zz_885 = 1'b1;
  assign _zz_2021 = _zz_9354;
  assign _zz_2022 = _zz_9362;
  assign _zz_888 = ($signed(_zz_9370) * $signed(data_mid_5_49_real));
  assign _zz_2023 = _zz_9371;
  assign _zz_886 = _zz_9374[35 : 0];
  assign _zz_2024 = _zz_9375;
  assign _zz_887 = _zz_9378[35 : 0];
  assign _zz_889 = 1'b1;
  assign _zz_2025 = _zz_9379;
  assign _zz_2026 = _zz_9387;
  assign _zz_890 = 1'b1;
  assign _zz_2027 = _zz_9395;
  assign _zz_2028 = _zz_9403;
  assign _zz_893 = ($signed(_zz_9411) * $signed(data_mid_5_50_real));
  assign _zz_2029 = _zz_9412;
  assign _zz_891 = _zz_9415[35 : 0];
  assign _zz_2030 = _zz_9416;
  assign _zz_892 = _zz_9419[35 : 0];
  assign _zz_894 = 1'b1;
  assign _zz_2031 = _zz_9420;
  assign _zz_2032 = _zz_9428;
  assign _zz_895 = 1'b1;
  assign _zz_2033 = _zz_9436;
  assign _zz_2034 = _zz_9444;
  assign _zz_898 = ($signed(_zz_9452) * $signed(data_mid_5_51_real));
  assign _zz_2035 = _zz_9453;
  assign _zz_896 = _zz_9456[35 : 0];
  assign _zz_2036 = _zz_9457;
  assign _zz_897 = _zz_9460[35 : 0];
  assign _zz_899 = 1'b1;
  assign _zz_2037 = _zz_9461;
  assign _zz_2038 = _zz_9469;
  assign _zz_900 = 1'b1;
  assign _zz_2039 = _zz_9477;
  assign _zz_2040 = _zz_9485;
  assign _zz_903 = ($signed(_zz_9493) * $signed(data_mid_5_52_real));
  assign _zz_2041 = _zz_9494;
  assign _zz_901 = _zz_9497[35 : 0];
  assign _zz_2042 = _zz_9498;
  assign _zz_902 = _zz_9501[35 : 0];
  assign _zz_904 = 1'b1;
  assign _zz_2043 = _zz_9502;
  assign _zz_2044 = _zz_9510;
  assign _zz_905 = 1'b1;
  assign _zz_2045 = _zz_9518;
  assign _zz_2046 = _zz_9526;
  assign _zz_908 = ($signed(_zz_9534) * $signed(data_mid_5_53_real));
  assign _zz_2047 = _zz_9535;
  assign _zz_906 = _zz_9538[35 : 0];
  assign _zz_2048 = _zz_9539;
  assign _zz_907 = _zz_9542[35 : 0];
  assign _zz_909 = 1'b1;
  assign _zz_2049 = _zz_9543;
  assign _zz_2050 = _zz_9551;
  assign _zz_910 = 1'b1;
  assign _zz_2051 = _zz_9559;
  assign _zz_2052 = _zz_9567;
  assign _zz_913 = ($signed(_zz_9575) * $signed(data_mid_5_54_real));
  assign _zz_2053 = _zz_9576;
  assign _zz_911 = _zz_9579[35 : 0];
  assign _zz_2054 = _zz_9580;
  assign _zz_912 = _zz_9583[35 : 0];
  assign _zz_914 = 1'b1;
  assign _zz_2055 = _zz_9584;
  assign _zz_2056 = _zz_9592;
  assign _zz_915 = 1'b1;
  assign _zz_2057 = _zz_9600;
  assign _zz_2058 = _zz_9608;
  assign _zz_918 = ($signed(_zz_9616) * $signed(data_mid_5_55_real));
  assign _zz_2059 = _zz_9617;
  assign _zz_916 = _zz_9620[35 : 0];
  assign _zz_2060 = _zz_9621;
  assign _zz_917 = _zz_9624[35 : 0];
  assign _zz_919 = 1'b1;
  assign _zz_2061 = _zz_9625;
  assign _zz_2062 = _zz_9633;
  assign _zz_920 = 1'b1;
  assign _zz_2063 = _zz_9641;
  assign _zz_2064 = _zz_9649;
  assign _zz_923 = ($signed(_zz_9657) * $signed(data_mid_5_56_real));
  assign _zz_2065 = _zz_9658;
  assign _zz_921 = _zz_9661[35 : 0];
  assign _zz_2066 = _zz_9662;
  assign _zz_922 = _zz_9665[35 : 0];
  assign _zz_924 = 1'b1;
  assign _zz_2067 = _zz_9666;
  assign _zz_2068 = _zz_9674;
  assign _zz_925 = 1'b1;
  assign _zz_2069 = _zz_9682;
  assign _zz_2070 = _zz_9690;
  assign _zz_928 = ($signed(_zz_9698) * $signed(data_mid_5_57_real));
  assign _zz_2071 = _zz_9699;
  assign _zz_926 = _zz_9702[35 : 0];
  assign _zz_2072 = _zz_9703;
  assign _zz_927 = _zz_9706[35 : 0];
  assign _zz_929 = 1'b1;
  assign _zz_2073 = _zz_9707;
  assign _zz_2074 = _zz_9715;
  assign _zz_930 = 1'b1;
  assign _zz_2075 = _zz_9723;
  assign _zz_2076 = _zz_9731;
  assign _zz_933 = ($signed(_zz_9739) * $signed(data_mid_5_58_real));
  assign _zz_2077 = _zz_9740;
  assign _zz_931 = _zz_9743[35 : 0];
  assign _zz_2078 = _zz_9744;
  assign _zz_932 = _zz_9747[35 : 0];
  assign _zz_934 = 1'b1;
  assign _zz_2079 = _zz_9748;
  assign _zz_2080 = _zz_9756;
  assign _zz_935 = 1'b1;
  assign _zz_2081 = _zz_9764;
  assign _zz_2082 = _zz_9772;
  assign _zz_938 = ($signed(_zz_9780) * $signed(data_mid_5_59_real));
  assign _zz_2083 = _zz_9781;
  assign _zz_936 = _zz_9784[35 : 0];
  assign _zz_2084 = _zz_9785;
  assign _zz_937 = _zz_9788[35 : 0];
  assign _zz_939 = 1'b1;
  assign _zz_2085 = _zz_9789;
  assign _zz_2086 = _zz_9797;
  assign _zz_940 = 1'b1;
  assign _zz_2087 = _zz_9805;
  assign _zz_2088 = _zz_9813;
  assign _zz_943 = ($signed(_zz_9821) * $signed(data_mid_5_60_real));
  assign _zz_2089 = _zz_9822;
  assign _zz_941 = _zz_9825[35 : 0];
  assign _zz_2090 = _zz_9826;
  assign _zz_942 = _zz_9829[35 : 0];
  assign _zz_944 = 1'b1;
  assign _zz_2091 = _zz_9830;
  assign _zz_2092 = _zz_9838;
  assign _zz_945 = 1'b1;
  assign _zz_2093 = _zz_9846;
  assign _zz_2094 = _zz_9854;
  assign _zz_948 = ($signed(_zz_9862) * $signed(data_mid_5_61_real));
  assign _zz_2095 = _zz_9863;
  assign _zz_946 = _zz_9866[35 : 0];
  assign _zz_2096 = _zz_9867;
  assign _zz_947 = _zz_9870[35 : 0];
  assign _zz_949 = 1'b1;
  assign _zz_2097 = _zz_9871;
  assign _zz_2098 = _zz_9879;
  assign _zz_950 = 1'b1;
  assign _zz_2099 = _zz_9887;
  assign _zz_2100 = _zz_9895;
  assign _zz_953 = ($signed(_zz_9903) * $signed(data_mid_5_62_real));
  assign _zz_2101 = _zz_9904;
  assign _zz_951 = _zz_9907[35 : 0];
  assign _zz_2102 = _zz_9908;
  assign _zz_952 = _zz_9911[35 : 0];
  assign _zz_954 = 1'b1;
  assign _zz_2103 = _zz_9912;
  assign _zz_2104 = _zz_9920;
  assign _zz_955 = 1'b1;
  assign _zz_2105 = _zz_9928;
  assign _zz_2106 = _zz_9936;
  assign _zz_958 = ($signed(_zz_9944) * $signed(data_mid_5_63_real));
  assign _zz_2107 = _zz_9945;
  assign _zz_956 = _zz_9948[35 : 0];
  assign _zz_2108 = _zz_9949;
  assign _zz_957 = _zz_9952[35 : 0];
  assign _zz_959 = 1'b1;
  assign _zz_2109 = _zz_9953;
  assign _zz_2110 = _zz_9961;
  assign _zz_960 = 1'b1;
  assign _zz_2111 = _zz_9969;
  assign _zz_2112 = _zz_9977;
  assign fft_col_out_valid = io_data_in_valid_delay_8;
  assign fft_col_out_payload_0_real = data_mid_6_0_real;
  assign fft_col_out_payload_0_imag = data_mid_6_0_imag;
  assign fft_col_out_payload_1_real = data_mid_6_1_real;
  assign fft_col_out_payload_1_imag = data_mid_6_1_imag;
  assign fft_col_out_payload_2_real = data_mid_6_2_real;
  assign fft_col_out_payload_2_imag = data_mid_6_2_imag;
  assign fft_col_out_payload_3_real = data_mid_6_3_real;
  assign fft_col_out_payload_3_imag = data_mid_6_3_imag;
  assign fft_col_out_payload_4_real = data_mid_6_4_real;
  assign fft_col_out_payload_4_imag = data_mid_6_4_imag;
  assign fft_col_out_payload_5_real = data_mid_6_5_real;
  assign fft_col_out_payload_5_imag = data_mid_6_5_imag;
  assign fft_col_out_payload_6_real = data_mid_6_6_real;
  assign fft_col_out_payload_6_imag = data_mid_6_6_imag;
  assign fft_col_out_payload_7_real = data_mid_6_7_real;
  assign fft_col_out_payload_7_imag = data_mid_6_7_imag;
  assign fft_col_out_payload_8_real = data_mid_6_8_real;
  assign fft_col_out_payload_8_imag = data_mid_6_8_imag;
  assign fft_col_out_payload_9_real = data_mid_6_9_real;
  assign fft_col_out_payload_9_imag = data_mid_6_9_imag;
  assign fft_col_out_payload_10_real = data_mid_6_10_real;
  assign fft_col_out_payload_10_imag = data_mid_6_10_imag;
  assign fft_col_out_payload_11_real = data_mid_6_11_real;
  assign fft_col_out_payload_11_imag = data_mid_6_11_imag;
  assign fft_col_out_payload_12_real = data_mid_6_12_real;
  assign fft_col_out_payload_12_imag = data_mid_6_12_imag;
  assign fft_col_out_payload_13_real = data_mid_6_13_real;
  assign fft_col_out_payload_13_imag = data_mid_6_13_imag;
  assign fft_col_out_payload_14_real = data_mid_6_14_real;
  assign fft_col_out_payload_14_imag = data_mid_6_14_imag;
  assign fft_col_out_payload_15_real = data_mid_6_15_real;
  assign fft_col_out_payload_15_imag = data_mid_6_15_imag;
  assign fft_col_out_payload_16_real = data_mid_6_16_real;
  assign fft_col_out_payload_16_imag = data_mid_6_16_imag;
  assign fft_col_out_payload_17_real = data_mid_6_17_real;
  assign fft_col_out_payload_17_imag = data_mid_6_17_imag;
  assign fft_col_out_payload_18_real = data_mid_6_18_real;
  assign fft_col_out_payload_18_imag = data_mid_6_18_imag;
  assign fft_col_out_payload_19_real = data_mid_6_19_real;
  assign fft_col_out_payload_19_imag = data_mid_6_19_imag;
  assign fft_col_out_payload_20_real = data_mid_6_20_real;
  assign fft_col_out_payload_20_imag = data_mid_6_20_imag;
  assign fft_col_out_payload_21_real = data_mid_6_21_real;
  assign fft_col_out_payload_21_imag = data_mid_6_21_imag;
  assign fft_col_out_payload_22_real = data_mid_6_22_real;
  assign fft_col_out_payload_22_imag = data_mid_6_22_imag;
  assign fft_col_out_payload_23_real = data_mid_6_23_real;
  assign fft_col_out_payload_23_imag = data_mid_6_23_imag;
  assign fft_col_out_payload_24_real = data_mid_6_24_real;
  assign fft_col_out_payload_24_imag = data_mid_6_24_imag;
  assign fft_col_out_payload_25_real = data_mid_6_25_real;
  assign fft_col_out_payload_25_imag = data_mid_6_25_imag;
  assign fft_col_out_payload_26_real = data_mid_6_26_real;
  assign fft_col_out_payload_26_imag = data_mid_6_26_imag;
  assign fft_col_out_payload_27_real = data_mid_6_27_real;
  assign fft_col_out_payload_27_imag = data_mid_6_27_imag;
  assign fft_col_out_payload_28_real = data_mid_6_28_real;
  assign fft_col_out_payload_28_imag = data_mid_6_28_imag;
  assign fft_col_out_payload_29_real = data_mid_6_29_real;
  assign fft_col_out_payload_29_imag = data_mid_6_29_imag;
  assign fft_col_out_payload_30_real = data_mid_6_30_real;
  assign fft_col_out_payload_30_imag = data_mid_6_30_imag;
  assign fft_col_out_payload_31_real = data_mid_6_31_real;
  assign fft_col_out_payload_31_imag = data_mid_6_31_imag;
  assign fft_col_out_payload_32_real = data_mid_6_32_real;
  assign fft_col_out_payload_32_imag = data_mid_6_32_imag;
  assign fft_col_out_payload_33_real = data_mid_6_33_real;
  assign fft_col_out_payload_33_imag = data_mid_6_33_imag;
  assign fft_col_out_payload_34_real = data_mid_6_34_real;
  assign fft_col_out_payload_34_imag = data_mid_6_34_imag;
  assign fft_col_out_payload_35_real = data_mid_6_35_real;
  assign fft_col_out_payload_35_imag = data_mid_6_35_imag;
  assign fft_col_out_payload_36_real = data_mid_6_36_real;
  assign fft_col_out_payload_36_imag = data_mid_6_36_imag;
  assign fft_col_out_payload_37_real = data_mid_6_37_real;
  assign fft_col_out_payload_37_imag = data_mid_6_37_imag;
  assign fft_col_out_payload_38_real = data_mid_6_38_real;
  assign fft_col_out_payload_38_imag = data_mid_6_38_imag;
  assign fft_col_out_payload_39_real = data_mid_6_39_real;
  assign fft_col_out_payload_39_imag = data_mid_6_39_imag;
  assign fft_col_out_payload_40_real = data_mid_6_40_real;
  assign fft_col_out_payload_40_imag = data_mid_6_40_imag;
  assign fft_col_out_payload_41_real = data_mid_6_41_real;
  assign fft_col_out_payload_41_imag = data_mid_6_41_imag;
  assign fft_col_out_payload_42_real = data_mid_6_42_real;
  assign fft_col_out_payload_42_imag = data_mid_6_42_imag;
  assign fft_col_out_payload_43_real = data_mid_6_43_real;
  assign fft_col_out_payload_43_imag = data_mid_6_43_imag;
  assign fft_col_out_payload_44_real = data_mid_6_44_real;
  assign fft_col_out_payload_44_imag = data_mid_6_44_imag;
  assign fft_col_out_payload_45_real = data_mid_6_45_real;
  assign fft_col_out_payload_45_imag = data_mid_6_45_imag;
  assign fft_col_out_payload_46_real = data_mid_6_46_real;
  assign fft_col_out_payload_46_imag = data_mid_6_46_imag;
  assign fft_col_out_payload_47_real = data_mid_6_47_real;
  assign fft_col_out_payload_47_imag = data_mid_6_47_imag;
  assign fft_col_out_payload_48_real = data_mid_6_48_real;
  assign fft_col_out_payload_48_imag = data_mid_6_48_imag;
  assign fft_col_out_payload_49_real = data_mid_6_49_real;
  assign fft_col_out_payload_49_imag = data_mid_6_49_imag;
  assign fft_col_out_payload_50_real = data_mid_6_50_real;
  assign fft_col_out_payload_50_imag = data_mid_6_50_imag;
  assign fft_col_out_payload_51_real = data_mid_6_51_real;
  assign fft_col_out_payload_51_imag = data_mid_6_51_imag;
  assign fft_col_out_payload_52_real = data_mid_6_52_real;
  assign fft_col_out_payload_52_imag = data_mid_6_52_imag;
  assign fft_col_out_payload_53_real = data_mid_6_53_real;
  assign fft_col_out_payload_53_imag = data_mid_6_53_imag;
  assign fft_col_out_payload_54_real = data_mid_6_54_real;
  assign fft_col_out_payload_54_imag = data_mid_6_54_imag;
  assign fft_col_out_payload_55_real = data_mid_6_55_real;
  assign fft_col_out_payload_55_imag = data_mid_6_55_imag;
  assign fft_col_out_payload_56_real = data_mid_6_56_real;
  assign fft_col_out_payload_56_imag = data_mid_6_56_imag;
  assign fft_col_out_payload_57_real = data_mid_6_57_real;
  assign fft_col_out_payload_57_imag = data_mid_6_57_imag;
  assign fft_col_out_payload_58_real = data_mid_6_58_real;
  assign fft_col_out_payload_58_imag = data_mid_6_58_imag;
  assign fft_col_out_payload_59_real = data_mid_6_59_real;
  assign fft_col_out_payload_59_imag = data_mid_6_59_imag;
  assign fft_col_out_payload_60_real = data_mid_6_60_real;
  assign fft_col_out_payload_60_imag = data_mid_6_60_imag;
  assign fft_col_out_payload_61_real = data_mid_6_61_real;
  assign fft_col_out_payload_61_imag = data_mid_6_61_imag;
  assign fft_col_out_payload_62_real = data_mid_6_62_real;
  assign fft_col_out_payload_62_imag = data_mid_6_62_imag;
  assign fft_col_out_payload_63_real = data_mid_6_63_real;
  assign fft_col_out_payload_63_imag = data_mid_6_63_imag;
  always @ (posedge clk) begin
    if(io_data_in_valid)begin
      data_in_0_real <= io_data_in_payload_0_real;
      data_in_0_imag <= io_data_in_payload_0_imag;
      data_in_1_real <= io_data_in_payload_1_real;
      data_in_1_imag <= io_data_in_payload_1_imag;
      data_in_2_real <= io_data_in_payload_2_real;
      data_in_2_imag <= io_data_in_payload_2_imag;
      data_in_3_real <= io_data_in_payload_3_real;
      data_in_3_imag <= io_data_in_payload_3_imag;
      data_in_4_real <= io_data_in_payload_4_real;
      data_in_4_imag <= io_data_in_payload_4_imag;
      data_in_5_real <= io_data_in_payload_5_real;
      data_in_5_imag <= io_data_in_payload_5_imag;
      data_in_6_real <= io_data_in_payload_6_real;
      data_in_6_imag <= io_data_in_payload_6_imag;
      data_in_7_real <= io_data_in_payload_7_real;
      data_in_7_imag <= io_data_in_payload_7_imag;
      data_in_8_real <= io_data_in_payload_8_real;
      data_in_8_imag <= io_data_in_payload_8_imag;
      data_in_9_real <= io_data_in_payload_9_real;
      data_in_9_imag <= io_data_in_payload_9_imag;
      data_in_10_real <= io_data_in_payload_10_real;
      data_in_10_imag <= io_data_in_payload_10_imag;
      data_in_11_real <= io_data_in_payload_11_real;
      data_in_11_imag <= io_data_in_payload_11_imag;
      data_in_12_real <= io_data_in_payload_12_real;
      data_in_12_imag <= io_data_in_payload_12_imag;
      data_in_13_real <= io_data_in_payload_13_real;
      data_in_13_imag <= io_data_in_payload_13_imag;
      data_in_14_real <= io_data_in_payload_14_real;
      data_in_14_imag <= io_data_in_payload_14_imag;
      data_in_15_real <= io_data_in_payload_15_real;
      data_in_15_imag <= io_data_in_payload_15_imag;
      data_in_16_real <= io_data_in_payload_16_real;
      data_in_16_imag <= io_data_in_payload_16_imag;
      data_in_17_real <= io_data_in_payload_17_real;
      data_in_17_imag <= io_data_in_payload_17_imag;
      data_in_18_real <= io_data_in_payload_18_real;
      data_in_18_imag <= io_data_in_payload_18_imag;
      data_in_19_real <= io_data_in_payload_19_real;
      data_in_19_imag <= io_data_in_payload_19_imag;
      data_in_20_real <= io_data_in_payload_20_real;
      data_in_20_imag <= io_data_in_payload_20_imag;
      data_in_21_real <= io_data_in_payload_21_real;
      data_in_21_imag <= io_data_in_payload_21_imag;
      data_in_22_real <= io_data_in_payload_22_real;
      data_in_22_imag <= io_data_in_payload_22_imag;
      data_in_23_real <= io_data_in_payload_23_real;
      data_in_23_imag <= io_data_in_payload_23_imag;
      data_in_24_real <= io_data_in_payload_24_real;
      data_in_24_imag <= io_data_in_payload_24_imag;
      data_in_25_real <= io_data_in_payload_25_real;
      data_in_25_imag <= io_data_in_payload_25_imag;
      data_in_26_real <= io_data_in_payload_26_real;
      data_in_26_imag <= io_data_in_payload_26_imag;
      data_in_27_real <= io_data_in_payload_27_real;
      data_in_27_imag <= io_data_in_payload_27_imag;
      data_in_28_real <= io_data_in_payload_28_real;
      data_in_28_imag <= io_data_in_payload_28_imag;
      data_in_29_real <= io_data_in_payload_29_real;
      data_in_29_imag <= io_data_in_payload_29_imag;
      data_in_30_real <= io_data_in_payload_30_real;
      data_in_30_imag <= io_data_in_payload_30_imag;
      data_in_31_real <= io_data_in_payload_31_real;
      data_in_31_imag <= io_data_in_payload_31_imag;
      data_in_32_real <= io_data_in_payload_32_real;
      data_in_32_imag <= io_data_in_payload_32_imag;
      data_in_33_real <= io_data_in_payload_33_real;
      data_in_33_imag <= io_data_in_payload_33_imag;
      data_in_34_real <= io_data_in_payload_34_real;
      data_in_34_imag <= io_data_in_payload_34_imag;
      data_in_35_real <= io_data_in_payload_35_real;
      data_in_35_imag <= io_data_in_payload_35_imag;
      data_in_36_real <= io_data_in_payload_36_real;
      data_in_36_imag <= io_data_in_payload_36_imag;
      data_in_37_real <= io_data_in_payload_37_real;
      data_in_37_imag <= io_data_in_payload_37_imag;
      data_in_38_real <= io_data_in_payload_38_real;
      data_in_38_imag <= io_data_in_payload_38_imag;
      data_in_39_real <= io_data_in_payload_39_real;
      data_in_39_imag <= io_data_in_payload_39_imag;
      data_in_40_real <= io_data_in_payload_40_real;
      data_in_40_imag <= io_data_in_payload_40_imag;
      data_in_41_real <= io_data_in_payload_41_real;
      data_in_41_imag <= io_data_in_payload_41_imag;
      data_in_42_real <= io_data_in_payload_42_real;
      data_in_42_imag <= io_data_in_payload_42_imag;
      data_in_43_real <= io_data_in_payload_43_real;
      data_in_43_imag <= io_data_in_payload_43_imag;
      data_in_44_real <= io_data_in_payload_44_real;
      data_in_44_imag <= io_data_in_payload_44_imag;
      data_in_45_real <= io_data_in_payload_45_real;
      data_in_45_imag <= io_data_in_payload_45_imag;
      data_in_46_real <= io_data_in_payload_46_real;
      data_in_46_imag <= io_data_in_payload_46_imag;
      data_in_47_real <= io_data_in_payload_47_real;
      data_in_47_imag <= io_data_in_payload_47_imag;
      data_in_48_real <= io_data_in_payload_48_real;
      data_in_48_imag <= io_data_in_payload_48_imag;
      data_in_49_real <= io_data_in_payload_49_real;
      data_in_49_imag <= io_data_in_payload_49_imag;
      data_in_50_real <= io_data_in_payload_50_real;
      data_in_50_imag <= io_data_in_payload_50_imag;
      data_in_51_real <= io_data_in_payload_51_real;
      data_in_51_imag <= io_data_in_payload_51_imag;
      data_in_52_real <= io_data_in_payload_52_real;
      data_in_52_imag <= io_data_in_payload_52_imag;
      data_in_53_real <= io_data_in_payload_53_real;
      data_in_53_imag <= io_data_in_payload_53_imag;
      data_in_54_real <= io_data_in_payload_54_real;
      data_in_54_imag <= io_data_in_payload_54_imag;
      data_in_55_real <= io_data_in_payload_55_real;
      data_in_55_imag <= io_data_in_payload_55_imag;
      data_in_56_real <= io_data_in_payload_56_real;
      data_in_56_imag <= io_data_in_payload_56_imag;
      data_in_57_real <= io_data_in_payload_57_real;
      data_in_57_imag <= io_data_in_payload_57_imag;
      data_in_58_real <= io_data_in_payload_58_real;
      data_in_58_imag <= io_data_in_payload_58_imag;
      data_in_59_real <= io_data_in_payload_59_real;
      data_in_59_imag <= io_data_in_payload_59_imag;
      data_in_60_real <= io_data_in_payload_60_real;
      data_in_60_imag <= io_data_in_payload_60_imag;
      data_in_61_real <= io_data_in_payload_61_real;
      data_in_61_imag <= io_data_in_payload_61_imag;
      data_in_62_real <= io_data_in_payload_62_real;
      data_in_62_imag <= io_data_in_payload_62_imag;
      data_in_63_real <= io_data_in_payload_63_real;
      data_in_63_imag <= io_data_in_payload_63_imag;
    end
    data_mid_0_0_real <= data_reorder_0_real;
    data_mid_0_0_imag <= data_reorder_0_imag;
    data_mid_0_1_real <= data_reorder_1_real;
    data_mid_0_1_imag <= data_reorder_1_imag;
    data_mid_0_2_real <= data_reorder_2_real;
    data_mid_0_2_imag <= data_reorder_2_imag;
    data_mid_0_3_real <= data_reorder_3_real;
    data_mid_0_3_imag <= data_reorder_3_imag;
    data_mid_0_4_real <= data_reorder_4_real;
    data_mid_0_4_imag <= data_reorder_4_imag;
    data_mid_0_5_real <= data_reorder_5_real;
    data_mid_0_5_imag <= data_reorder_5_imag;
    data_mid_0_6_real <= data_reorder_6_real;
    data_mid_0_6_imag <= data_reorder_6_imag;
    data_mid_0_7_real <= data_reorder_7_real;
    data_mid_0_7_imag <= data_reorder_7_imag;
    data_mid_0_8_real <= data_reorder_8_real;
    data_mid_0_8_imag <= data_reorder_8_imag;
    data_mid_0_9_real <= data_reorder_9_real;
    data_mid_0_9_imag <= data_reorder_9_imag;
    data_mid_0_10_real <= data_reorder_10_real;
    data_mid_0_10_imag <= data_reorder_10_imag;
    data_mid_0_11_real <= data_reorder_11_real;
    data_mid_0_11_imag <= data_reorder_11_imag;
    data_mid_0_12_real <= data_reorder_12_real;
    data_mid_0_12_imag <= data_reorder_12_imag;
    data_mid_0_13_real <= data_reorder_13_real;
    data_mid_0_13_imag <= data_reorder_13_imag;
    data_mid_0_14_real <= data_reorder_14_real;
    data_mid_0_14_imag <= data_reorder_14_imag;
    data_mid_0_15_real <= data_reorder_15_real;
    data_mid_0_15_imag <= data_reorder_15_imag;
    data_mid_0_16_real <= data_reorder_16_real;
    data_mid_0_16_imag <= data_reorder_16_imag;
    data_mid_0_17_real <= data_reorder_17_real;
    data_mid_0_17_imag <= data_reorder_17_imag;
    data_mid_0_18_real <= data_reorder_18_real;
    data_mid_0_18_imag <= data_reorder_18_imag;
    data_mid_0_19_real <= data_reorder_19_real;
    data_mid_0_19_imag <= data_reorder_19_imag;
    data_mid_0_20_real <= data_reorder_20_real;
    data_mid_0_20_imag <= data_reorder_20_imag;
    data_mid_0_21_real <= data_reorder_21_real;
    data_mid_0_21_imag <= data_reorder_21_imag;
    data_mid_0_22_real <= data_reorder_22_real;
    data_mid_0_22_imag <= data_reorder_22_imag;
    data_mid_0_23_real <= data_reorder_23_real;
    data_mid_0_23_imag <= data_reorder_23_imag;
    data_mid_0_24_real <= data_reorder_24_real;
    data_mid_0_24_imag <= data_reorder_24_imag;
    data_mid_0_25_real <= data_reorder_25_real;
    data_mid_0_25_imag <= data_reorder_25_imag;
    data_mid_0_26_real <= data_reorder_26_real;
    data_mid_0_26_imag <= data_reorder_26_imag;
    data_mid_0_27_real <= data_reorder_27_real;
    data_mid_0_27_imag <= data_reorder_27_imag;
    data_mid_0_28_real <= data_reorder_28_real;
    data_mid_0_28_imag <= data_reorder_28_imag;
    data_mid_0_29_real <= data_reorder_29_real;
    data_mid_0_29_imag <= data_reorder_29_imag;
    data_mid_0_30_real <= data_reorder_30_real;
    data_mid_0_30_imag <= data_reorder_30_imag;
    data_mid_0_31_real <= data_reorder_31_real;
    data_mid_0_31_imag <= data_reorder_31_imag;
    data_mid_0_32_real <= data_reorder_32_real;
    data_mid_0_32_imag <= data_reorder_32_imag;
    data_mid_0_33_real <= data_reorder_33_real;
    data_mid_0_33_imag <= data_reorder_33_imag;
    data_mid_0_34_real <= data_reorder_34_real;
    data_mid_0_34_imag <= data_reorder_34_imag;
    data_mid_0_35_real <= data_reorder_35_real;
    data_mid_0_35_imag <= data_reorder_35_imag;
    data_mid_0_36_real <= data_reorder_36_real;
    data_mid_0_36_imag <= data_reorder_36_imag;
    data_mid_0_37_real <= data_reorder_37_real;
    data_mid_0_37_imag <= data_reorder_37_imag;
    data_mid_0_38_real <= data_reorder_38_real;
    data_mid_0_38_imag <= data_reorder_38_imag;
    data_mid_0_39_real <= data_reorder_39_real;
    data_mid_0_39_imag <= data_reorder_39_imag;
    data_mid_0_40_real <= data_reorder_40_real;
    data_mid_0_40_imag <= data_reorder_40_imag;
    data_mid_0_41_real <= data_reorder_41_real;
    data_mid_0_41_imag <= data_reorder_41_imag;
    data_mid_0_42_real <= data_reorder_42_real;
    data_mid_0_42_imag <= data_reorder_42_imag;
    data_mid_0_43_real <= data_reorder_43_real;
    data_mid_0_43_imag <= data_reorder_43_imag;
    data_mid_0_44_real <= data_reorder_44_real;
    data_mid_0_44_imag <= data_reorder_44_imag;
    data_mid_0_45_real <= data_reorder_45_real;
    data_mid_0_45_imag <= data_reorder_45_imag;
    data_mid_0_46_real <= data_reorder_46_real;
    data_mid_0_46_imag <= data_reorder_46_imag;
    data_mid_0_47_real <= data_reorder_47_real;
    data_mid_0_47_imag <= data_reorder_47_imag;
    data_mid_0_48_real <= data_reorder_48_real;
    data_mid_0_48_imag <= data_reorder_48_imag;
    data_mid_0_49_real <= data_reorder_49_real;
    data_mid_0_49_imag <= data_reorder_49_imag;
    data_mid_0_50_real <= data_reorder_50_real;
    data_mid_0_50_imag <= data_reorder_50_imag;
    data_mid_0_51_real <= data_reorder_51_real;
    data_mid_0_51_imag <= data_reorder_51_imag;
    data_mid_0_52_real <= data_reorder_52_real;
    data_mid_0_52_imag <= data_reorder_52_imag;
    data_mid_0_53_real <= data_reorder_53_real;
    data_mid_0_53_imag <= data_reorder_53_imag;
    data_mid_0_54_real <= data_reorder_54_real;
    data_mid_0_54_imag <= data_reorder_54_imag;
    data_mid_0_55_real <= data_reorder_55_real;
    data_mid_0_55_imag <= data_reorder_55_imag;
    data_mid_0_56_real <= data_reorder_56_real;
    data_mid_0_56_imag <= data_reorder_56_imag;
    data_mid_0_57_real <= data_reorder_57_real;
    data_mid_0_57_imag <= data_reorder_57_imag;
    data_mid_0_58_real <= data_reorder_58_real;
    data_mid_0_58_imag <= data_reorder_58_imag;
    data_mid_0_59_real <= data_reorder_59_real;
    data_mid_0_59_imag <= data_reorder_59_imag;
    data_mid_0_60_real <= data_reorder_60_real;
    data_mid_0_60_imag <= data_reorder_60_imag;
    data_mid_0_61_real <= data_reorder_61_real;
    data_mid_0_61_imag <= data_reorder_61_imag;
    data_mid_0_62_real <= data_reorder_62_real;
    data_mid_0_62_imag <= data_reorder_62_imag;
    data_mid_0_63_real <= data_reorder_63_real;
    data_mid_0_63_imag <= data_reorder_63_imag;
    data_mid_1_1_real <= _zz_2129[17 : 0];
    data_mid_1_1_imag <= _zz_2137[17 : 0];
    data_mid_1_0_real <= _zz_2145[17 : 0];
    data_mid_1_0_imag <= _zz_2153[17 : 0];
    data_mid_1_3_real <= _zz_2170[17 : 0];
    data_mid_1_3_imag <= _zz_2178[17 : 0];
    data_mid_1_2_real <= _zz_2186[17 : 0];
    data_mid_1_2_imag <= _zz_2194[17 : 0];
    data_mid_1_5_real <= _zz_2211[17 : 0];
    data_mid_1_5_imag <= _zz_2219[17 : 0];
    data_mid_1_4_real <= _zz_2227[17 : 0];
    data_mid_1_4_imag <= _zz_2235[17 : 0];
    data_mid_1_7_real <= _zz_2252[17 : 0];
    data_mid_1_7_imag <= _zz_2260[17 : 0];
    data_mid_1_6_real <= _zz_2268[17 : 0];
    data_mid_1_6_imag <= _zz_2276[17 : 0];
    data_mid_1_9_real <= _zz_2293[17 : 0];
    data_mid_1_9_imag <= _zz_2301[17 : 0];
    data_mid_1_8_real <= _zz_2309[17 : 0];
    data_mid_1_8_imag <= _zz_2317[17 : 0];
    data_mid_1_11_real <= _zz_2334[17 : 0];
    data_mid_1_11_imag <= _zz_2342[17 : 0];
    data_mid_1_10_real <= _zz_2350[17 : 0];
    data_mid_1_10_imag <= _zz_2358[17 : 0];
    data_mid_1_13_real <= _zz_2375[17 : 0];
    data_mid_1_13_imag <= _zz_2383[17 : 0];
    data_mid_1_12_real <= _zz_2391[17 : 0];
    data_mid_1_12_imag <= _zz_2399[17 : 0];
    data_mid_1_15_real <= _zz_2416[17 : 0];
    data_mid_1_15_imag <= _zz_2424[17 : 0];
    data_mid_1_14_real <= _zz_2432[17 : 0];
    data_mid_1_14_imag <= _zz_2440[17 : 0];
    data_mid_1_17_real <= _zz_2457[17 : 0];
    data_mid_1_17_imag <= _zz_2465[17 : 0];
    data_mid_1_16_real <= _zz_2473[17 : 0];
    data_mid_1_16_imag <= _zz_2481[17 : 0];
    data_mid_1_19_real <= _zz_2498[17 : 0];
    data_mid_1_19_imag <= _zz_2506[17 : 0];
    data_mid_1_18_real <= _zz_2514[17 : 0];
    data_mid_1_18_imag <= _zz_2522[17 : 0];
    data_mid_1_21_real <= _zz_2539[17 : 0];
    data_mid_1_21_imag <= _zz_2547[17 : 0];
    data_mid_1_20_real <= _zz_2555[17 : 0];
    data_mid_1_20_imag <= _zz_2563[17 : 0];
    data_mid_1_23_real <= _zz_2580[17 : 0];
    data_mid_1_23_imag <= _zz_2588[17 : 0];
    data_mid_1_22_real <= _zz_2596[17 : 0];
    data_mid_1_22_imag <= _zz_2604[17 : 0];
    data_mid_1_25_real <= _zz_2621[17 : 0];
    data_mid_1_25_imag <= _zz_2629[17 : 0];
    data_mid_1_24_real <= _zz_2637[17 : 0];
    data_mid_1_24_imag <= _zz_2645[17 : 0];
    data_mid_1_27_real <= _zz_2662[17 : 0];
    data_mid_1_27_imag <= _zz_2670[17 : 0];
    data_mid_1_26_real <= _zz_2678[17 : 0];
    data_mid_1_26_imag <= _zz_2686[17 : 0];
    data_mid_1_29_real <= _zz_2703[17 : 0];
    data_mid_1_29_imag <= _zz_2711[17 : 0];
    data_mid_1_28_real <= _zz_2719[17 : 0];
    data_mid_1_28_imag <= _zz_2727[17 : 0];
    data_mid_1_31_real <= _zz_2744[17 : 0];
    data_mid_1_31_imag <= _zz_2752[17 : 0];
    data_mid_1_30_real <= _zz_2760[17 : 0];
    data_mid_1_30_imag <= _zz_2768[17 : 0];
    data_mid_1_33_real <= _zz_2785[17 : 0];
    data_mid_1_33_imag <= _zz_2793[17 : 0];
    data_mid_1_32_real <= _zz_2801[17 : 0];
    data_mid_1_32_imag <= _zz_2809[17 : 0];
    data_mid_1_35_real <= _zz_2826[17 : 0];
    data_mid_1_35_imag <= _zz_2834[17 : 0];
    data_mid_1_34_real <= _zz_2842[17 : 0];
    data_mid_1_34_imag <= _zz_2850[17 : 0];
    data_mid_1_37_real <= _zz_2867[17 : 0];
    data_mid_1_37_imag <= _zz_2875[17 : 0];
    data_mid_1_36_real <= _zz_2883[17 : 0];
    data_mid_1_36_imag <= _zz_2891[17 : 0];
    data_mid_1_39_real <= _zz_2908[17 : 0];
    data_mid_1_39_imag <= _zz_2916[17 : 0];
    data_mid_1_38_real <= _zz_2924[17 : 0];
    data_mid_1_38_imag <= _zz_2932[17 : 0];
    data_mid_1_41_real <= _zz_2949[17 : 0];
    data_mid_1_41_imag <= _zz_2957[17 : 0];
    data_mid_1_40_real <= _zz_2965[17 : 0];
    data_mid_1_40_imag <= _zz_2973[17 : 0];
    data_mid_1_43_real <= _zz_2990[17 : 0];
    data_mid_1_43_imag <= _zz_2998[17 : 0];
    data_mid_1_42_real <= _zz_3006[17 : 0];
    data_mid_1_42_imag <= _zz_3014[17 : 0];
    data_mid_1_45_real <= _zz_3031[17 : 0];
    data_mid_1_45_imag <= _zz_3039[17 : 0];
    data_mid_1_44_real <= _zz_3047[17 : 0];
    data_mid_1_44_imag <= _zz_3055[17 : 0];
    data_mid_1_47_real <= _zz_3072[17 : 0];
    data_mid_1_47_imag <= _zz_3080[17 : 0];
    data_mid_1_46_real <= _zz_3088[17 : 0];
    data_mid_1_46_imag <= _zz_3096[17 : 0];
    data_mid_1_49_real <= _zz_3113[17 : 0];
    data_mid_1_49_imag <= _zz_3121[17 : 0];
    data_mid_1_48_real <= _zz_3129[17 : 0];
    data_mid_1_48_imag <= _zz_3137[17 : 0];
    data_mid_1_51_real <= _zz_3154[17 : 0];
    data_mid_1_51_imag <= _zz_3162[17 : 0];
    data_mid_1_50_real <= _zz_3170[17 : 0];
    data_mid_1_50_imag <= _zz_3178[17 : 0];
    data_mid_1_53_real <= _zz_3195[17 : 0];
    data_mid_1_53_imag <= _zz_3203[17 : 0];
    data_mid_1_52_real <= _zz_3211[17 : 0];
    data_mid_1_52_imag <= _zz_3219[17 : 0];
    data_mid_1_55_real <= _zz_3236[17 : 0];
    data_mid_1_55_imag <= _zz_3244[17 : 0];
    data_mid_1_54_real <= _zz_3252[17 : 0];
    data_mid_1_54_imag <= _zz_3260[17 : 0];
    data_mid_1_57_real <= _zz_3277[17 : 0];
    data_mid_1_57_imag <= _zz_3285[17 : 0];
    data_mid_1_56_real <= _zz_3293[17 : 0];
    data_mid_1_56_imag <= _zz_3301[17 : 0];
    data_mid_1_59_real <= _zz_3318[17 : 0];
    data_mid_1_59_imag <= _zz_3326[17 : 0];
    data_mid_1_58_real <= _zz_3334[17 : 0];
    data_mid_1_58_imag <= _zz_3342[17 : 0];
    data_mid_1_61_real <= _zz_3359[17 : 0];
    data_mid_1_61_imag <= _zz_3367[17 : 0];
    data_mid_1_60_real <= _zz_3375[17 : 0];
    data_mid_1_60_imag <= _zz_3383[17 : 0];
    data_mid_1_63_real <= _zz_3400[17 : 0];
    data_mid_1_63_imag <= _zz_3408[17 : 0];
    data_mid_1_62_real <= _zz_3416[17 : 0];
    data_mid_1_62_imag <= _zz_3424[17 : 0];
    data_mid_2_2_real <= _zz_3441[17 : 0];
    data_mid_2_2_imag <= _zz_3449[17 : 0];
    data_mid_2_0_real <= _zz_3457[17 : 0];
    data_mid_2_0_imag <= _zz_3465[17 : 0];
    data_mid_2_3_real <= _zz_3482[17 : 0];
    data_mid_2_3_imag <= _zz_3490[17 : 0];
    data_mid_2_1_real <= _zz_3498[17 : 0];
    data_mid_2_1_imag <= _zz_3506[17 : 0];
    data_mid_2_6_real <= _zz_3523[17 : 0];
    data_mid_2_6_imag <= _zz_3531[17 : 0];
    data_mid_2_4_real <= _zz_3539[17 : 0];
    data_mid_2_4_imag <= _zz_3547[17 : 0];
    data_mid_2_7_real <= _zz_3564[17 : 0];
    data_mid_2_7_imag <= _zz_3572[17 : 0];
    data_mid_2_5_real <= _zz_3580[17 : 0];
    data_mid_2_5_imag <= _zz_3588[17 : 0];
    data_mid_2_10_real <= _zz_3605[17 : 0];
    data_mid_2_10_imag <= _zz_3613[17 : 0];
    data_mid_2_8_real <= _zz_3621[17 : 0];
    data_mid_2_8_imag <= _zz_3629[17 : 0];
    data_mid_2_11_real <= _zz_3646[17 : 0];
    data_mid_2_11_imag <= _zz_3654[17 : 0];
    data_mid_2_9_real <= _zz_3662[17 : 0];
    data_mid_2_9_imag <= _zz_3670[17 : 0];
    data_mid_2_14_real <= _zz_3687[17 : 0];
    data_mid_2_14_imag <= _zz_3695[17 : 0];
    data_mid_2_12_real <= _zz_3703[17 : 0];
    data_mid_2_12_imag <= _zz_3711[17 : 0];
    data_mid_2_15_real <= _zz_3728[17 : 0];
    data_mid_2_15_imag <= _zz_3736[17 : 0];
    data_mid_2_13_real <= _zz_3744[17 : 0];
    data_mid_2_13_imag <= _zz_3752[17 : 0];
    data_mid_2_18_real <= _zz_3769[17 : 0];
    data_mid_2_18_imag <= _zz_3777[17 : 0];
    data_mid_2_16_real <= _zz_3785[17 : 0];
    data_mid_2_16_imag <= _zz_3793[17 : 0];
    data_mid_2_19_real <= _zz_3810[17 : 0];
    data_mid_2_19_imag <= _zz_3818[17 : 0];
    data_mid_2_17_real <= _zz_3826[17 : 0];
    data_mid_2_17_imag <= _zz_3834[17 : 0];
    data_mid_2_22_real <= _zz_3851[17 : 0];
    data_mid_2_22_imag <= _zz_3859[17 : 0];
    data_mid_2_20_real <= _zz_3867[17 : 0];
    data_mid_2_20_imag <= _zz_3875[17 : 0];
    data_mid_2_23_real <= _zz_3892[17 : 0];
    data_mid_2_23_imag <= _zz_3900[17 : 0];
    data_mid_2_21_real <= _zz_3908[17 : 0];
    data_mid_2_21_imag <= _zz_3916[17 : 0];
    data_mid_2_26_real <= _zz_3933[17 : 0];
    data_mid_2_26_imag <= _zz_3941[17 : 0];
    data_mid_2_24_real <= _zz_3949[17 : 0];
    data_mid_2_24_imag <= _zz_3957[17 : 0];
    data_mid_2_27_real <= _zz_3974[17 : 0];
    data_mid_2_27_imag <= _zz_3982[17 : 0];
    data_mid_2_25_real <= _zz_3990[17 : 0];
    data_mid_2_25_imag <= _zz_3998[17 : 0];
    data_mid_2_30_real <= _zz_4015[17 : 0];
    data_mid_2_30_imag <= _zz_4023[17 : 0];
    data_mid_2_28_real <= _zz_4031[17 : 0];
    data_mid_2_28_imag <= _zz_4039[17 : 0];
    data_mid_2_31_real <= _zz_4056[17 : 0];
    data_mid_2_31_imag <= _zz_4064[17 : 0];
    data_mid_2_29_real <= _zz_4072[17 : 0];
    data_mid_2_29_imag <= _zz_4080[17 : 0];
    data_mid_2_34_real <= _zz_4097[17 : 0];
    data_mid_2_34_imag <= _zz_4105[17 : 0];
    data_mid_2_32_real <= _zz_4113[17 : 0];
    data_mid_2_32_imag <= _zz_4121[17 : 0];
    data_mid_2_35_real <= _zz_4138[17 : 0];
    data_mid_2_35_imag <= _zz_4146[17 : 0];
    data_mid_2_33_real <= _zz_4154[17 : 0];
    data_mid_2_33_imag <= _zz_4162[17 : 0];
    data_mid_2_38_real <= _zz_4179[17 : 0];
    data_mid_2_38_imag <= _zz_4187[17 : 0];
    data_mid_2_36_real <= _zz_4195[17 : 0];
    data_mid_2_36_imag <= _zz_4203[17 : 0];
    data_mid_2_39_real <= _zz_4220[17 : 0];
    data_mid_2_39_imag <= _zz_4228[17 : 0];
    data_mid_2_37_real <= _zz_4236[17 : 0];
    data_mid_2_37_imag <= _zz_4244[17 : 0];
    data_mid_2_42_real <= _zz_4261[17 : 0];
    data_mid_2_42_imag <= _zz_4269[17 : 0];
    data_mid_2_40_real <= _zz_4277[17 : 0];
    data_mid_2_40_imag <= _zz_4285[17 : 0];
    data_mid_2_43_real <= _zz_4302[17 : 0];
    data_mid_2_43_imag <= _zz_4310[17 : 0];
    data_mid_2_41_real <= _zz_4318[17 : 0];
    data_mid_2_41_imag <= _zz_4326[17 : 0];
    data_mid_2_46_real <= _zz_4343[17 : 0];
    data_mid_2_46_imag <= _zz_4351[17 : 0];
    data_mid_2_44_real <= _zz_4359[17 : 0];
    data_mid_2_44_imag <= _zz_4367[17 : 0];
    data_mid_2_47_real <= _zz_4384[17 : 0];
    data_mid_2_47_imag <= _zz_4392[17 : 0];
    data_mid_2_45_real <= _zz_4400[17 : 0];
    data_mid_2_45_imag <= _zz_4408[17 : 0];
    data_mid_2_50_real <= _zz_4425[17 : 0];
    data_mid_2_50_imag <= _zz_4433[17 : 0];
    data_mid_2_48_real <= _zz_4441[17 : 0];
    data_mid_2_48_imag <= _zz_4449[17 : 0];
    data_mid_2_51_real <= _zz_4466[17 : 0];
    data_mid_2_51_imag <= _zz_4474[17 : 0];
    data_mid_2_49_real <= _zz_4482[17 : 0];
    data_mid_2_49_imag <= _zz_4490[17 : 0];
    data_mid_2_54_real <= _zz_4507[17 : 0];
    data_mid_2_54_imag <= _zz_4515[17 : 0];
    data_mid_2_52_real <= _zz_4523[17 : 0];
    data_mid_2_52_imag <= _zz_4531[17 : 0];
    data_mid_2_55_real <= _zz_4548[17 : 0];
    data_mid_2_55_imag <= _zz_4556[17 : 0];
    data_mid_2_53_real <= _zz_4564[17 : 0];
    data_mid_2_53_imag <= _zz_4572[17 : 0];
    data_mid_2_58_real <= _zz_4589[17 : 0];
    data_mid_2_58_imag <= _zz_4597[17 : 0];
    data_mid_2_56_real <= _zz_4605[17 : 0];
    data_mid_2_56_imag <= _zz_4613[17 : 0];
    data_mid_2_59_real <= _zz_4630[17 : 0];
    data_mid_2_59_imag <= _zz_4638[17 : 0];
    data_mid_2_57_real <= _zz_4646[17 : 0];
    data_mid_2_57_imag <= _zz_4654[17 : 0];
    data_mid_2_62_real <= _zz_4671[17 : 0];
    data_mid_2_62_imag <= _zz_4679[17 : 0];
    data_mid_2_60_real <= _zz_4687[17 : 0];
    data_mid_2_60_imag <= _zz_4695[17 : 0];
    data_mid_2_63_real <= _zz_4712[17 : 0];
    data_mid_2_63_imag <= _zz_4720[17 : 0];
    data_mid_2_61_real <= _zz_4728[17 : 0];
    data_mid_2_61_imag <= _zz_4736[17 : 0];
    data_mid_3_4_real <= _zz_4753[17 : 0];
    data_mid_3_4_imag <= _zz_4761[17 : 0];
    data_mid_3_0_real <= _zz_4769[17 : 0];
    data_mid_3_0_imag <= _zz_4777[17 : 0];
    data_mid_3_5_real <= _zz_4794[17 : 0];
    data_mid_3_5_imag <= _zz_4802[17 : 0];
    data_mid_3_1_real <= _zz_4810[17 : 0];
    data_mid_3_1_imag <= _zz_4818[17 : 0];
    data_mid_3_6_real <= _zz_4835[17 : 0];
    data_mid_3_6_imag <= _zz_4843[17 : 0];
    data_mid_3_2_real <= _zz_4851[17 : 0];
    data_mid_3_2_imag <= _zz_4859[17 : 0];
    data_mid_3_7_real <= _zz_4876[17 : 0];
    data_mid_3_7_imag <= _zz_4884[17 : 0];
    data_mid_3_3_real <= _zz_4892[17 : 0];
    data_mid_3_3_imag <= _zz_4900[17 : 0];
    data_mid_3_12_real <= _zz_4917[17 : 0];
    data_mid_3_12_imag <= _zz_4925[17 : 0];
    data_mid_3_8_real <= _zz_4933[17 : 0];
    data_mid_3_8_imag <= _zz_4941[17 : 0];
    data_mid_3_13_real <= _zz_4958[17 : 0];
    data_mid_3_13_imag <= _zz_4966[17 : 0];
    data_mid_3_9_real <= _zz_4974[17 : 0];
    data_mid_3_9_imag <= _zz_4982[17 : 0];
    data_mid_3_14_real <= _zz_4999[17 : 0];
    data_mid_3_14_imag <= _zz_5007[17 : 0];
    data_mid_3_10_real <= _zz_5015[17 : 0];
    data_mid_3_10_imag <= _zz_5023[17 : 0];
    data_mid_3_15_real <= _zz_5040[17 : 0];
    data_mid_3_15_imag <= _zz_5048[17 : 0];
    data_mid_3_11_real <= _zz_5056[17 : 0];
    data_mid_3_11_imag <= _zz_5064[17 : 0];
    data_mid_3_20_real <= _zz_5081[17 : 0];
    data_mid_3_20_imag <= _zz_5089[17 : 0];
    data_mid_3_16_real <= _zz_5097[17 : 0];
    data_mid_3_16_imag <= _zz_5105[17 : 0];
    data_mid_3_21_real <= _zz_5122[17 : 0];
    data_mid_3_21_imag <= _zz_5130[17 : 0];
    data_mid_3_17_real <= _zz_5138[17 : 0];
    data_mid_3_17_imag <= _zz_5146[17 : 0];
    data_mid_3_22_real <= _zz_5163[17 : 0];
    data_mid_3_22_imag <= _zz_5171[17 : 0];
    data_mid_3_18_real <= _zz_5179[17 : 0];
    data_mid_3_18_imag <= _zz_5187[17 : 0];
    data_mid_3_23_real <= _zz_5204[17 : 0];
    data_mid_3_23_imag <= _zz_5212[17 : 0];
    data_mid_3_19_real <= _zz_5220[17 : 0];
    data_mid_3_19_imag <= _zz_5228[17 : 0];
    data_mid_3_28_real <= _zz_5245[17 : 0];
    data_mid_3_28_imag <= _zz_5253[17 : 0];
    data_mid_3_24_real <= _zz_5261[17 : 0];
    data_mid_3_24_imag <= _zz_5269[17 : 0];
    data_mid_3_29_real <= _zz_5286[17 : 0];
    data_mid_3_29_imag <= _zz_5294[17 : 0];
    data_mid_3_25_real <= _zz_5302[17 : 0];
    data_mid_3_25_imag <= _zz_5310[17 : 0];
    data_mid_3_30_real <= _zz_5327[17 : 0];
    data_mid_3_30_imag <= _zz_5335[17 : 0];
    data_mid_3_26_real <= _zz_5343[17 : 0];
    data_mid_3_26_imag <= _zz_5351[17 : 0];
    data_mid_3_31_real <= _zz_5368[17 : 0];
    data_mid_3_31_imag <= _zz_5376[17 : 0];
    data_mid_3_27_real <= _zz_5384[17 : 0];
    data_mid_3_27_imag <= _zz_5392[17 : 0];
    data_mid_3_36_real <= _zz_5409[17 : 0];
    data_mid_3_36_imag <= _zz_5417[17 : 0];
    data_mid_3_32_real <= _zz_5425[17 : 0];
    data_mid_3_32_imag <= _zz_5433[17 : 0];
    data_mid_3_37_real <= _zz_5450[17 : 0];
    data_mid_3_37_imag <= _zz_5458[17 : 0];
    data_mid_3_33_real <= _zz_5466[17 : 0];
    data_mid_3_33_imag <= _zz_5474[17 : 0];
    data_mid_3_38_real <= _zz_5491[17 : 0];
    data_mid_3_38_imag <= _zz_5499[17 : 0];
    data_mid_3_34_real <= _zz_5507[17 : 0];
    data_mid_3_34_imag <= _zz_5515[17 : 0];
    data_mid_3_39_real <= _zz_5532[17 : 0];
    data_mid_3_39_imag <= _zz_5540[17 : 0];
    data_mid_3_35_real <= _zz_5548[17 : 0];
    data_mid_3_35_imag <= _zz_5556[17 : 0];
    data_mid_3_44_real <= _zz_5573[17 : 0];
    data_mid_3_44_imag <= _zz_5581[17 : 0];
    data_mid_3_40_real <= _zz_5589[17 : 0];
    data_mid_3_40_imag <= _zz_5597[17 : 0];
    data_mid_3_45_real <= _zz_5614[17 : 0];
    data_mid_3_45_imag <= _zz_5622[17 : 0];
    data_mid_3_41_real <= _zz_5630[17 : 0];
    data_mid_3_41_imag <= _zz_5638[17 : 0];
    data_mid_3_46_real <= _zz_5655[17 : 0];
    data_mid_3_46_imag <= _zz_5663[17 : 0];
    data_mid_3_42_real <= _zz_5671[17 : 0];
    data_mid_3_42_imag <= _zz_5679[17 : 0];
    data_mid_3_47_real <= _zz_5696[17 : 0];
    data_mid_3_47_imag <= _zz_5704[17 : 0];
    data_mid_3_43_real <= _zz_5712[17 : 0];
    data_mid_3_43_imag <= _zz_5720[17 : 0];
    data_mid_3_52_real <= _zz_5737[17 : 0];
    data_mid_3_52_imag <= _zz_5745[17 : 0];
    data_mid_3_48_real <= _zz_5753[17 : 0];
    data_mid_3_48_imag <= _zz_5761[17 : 0];
    data_mid_3_53_real <= _zz_5778[17 : 0];
    data_mid_3_53_imag <= _zz_5786[17 : 0];
    data_mid_3_49_real <= _zz_5794[17 : 0];
    data_mid_3_49_imag <= _zz_5802[17 : 0];
    data_mid_3_54_real <= _zz_5819[17 : 0];
    data_mid_3_54_imag <= _zz_5827[17 : 0];
    data_mid_3_50_real <= _zz_5835[17 : 0];
    data_mid_3_50_imag <= _zz_5843[17 : 0];
    data_mid_3_55_real <= _zz_5860[17 : 0];
    data_mid_3_55_imag <= _zz_5868[17 : 0];
    data_mid_3_51_real <= _zz_5876[17 : 0];
    data_mid_3_51_imag <= _zz_5884[17 : 0];
    data_mid_3_60_real <= _zz_5901[17 : 0];
    data_mid_3_60_imag <= _zz_5909[17 : 0];
    data_mid_3_56_real <= _zz_5917[17 : 0];
    data_mid_3_56_imag <= _zz_5925[17 : 0];
    data_mid_3_61_real <= _zz_5942[17 : 0];
    data_mid_3_61_imag <= _zz_5950[17 : 0];
    data_mid_3_57_real <= _zz_5958[17 : 0];
    data_mid_3_57_imag <= _zz_5966[17 : 0];
    data_mid_3_62_real <= _zz_5983[17 : 0];
    data_mid_3_62_imag <= _zz_5991[17 : 0];
    data_mid_3_58_real <= _zz_5999[17 : 0];
    data_mid_3_58_imag <= _zz_6007[17 : 0];
    data_mid_3_63_real <= _zz_6024[17 : 0];
    data_mid_3_63_imag <= _zz_6032[17 : 0];
    data_mid_3_59_real <= _zz_6040[17 : 0];
    data_mid_3_59_imag <= _zz_6048[17 : 0];
    data_mid_4_8_real <= _zz_6065[17 : 0];
    data_mid_4_8_imag <= _zz_6073[17 : 0];
    data_mid_4_0_real <= _zz_6081[17 : 0];
    data_mid_4_0_imag <= _zz_6089[17 : 0];
    data_mid_4_9_real <= _zz_6106[17 : 0];
    data_mid_4_9_imag <= _zz_6114[17 : 0];
    data_mid_4_1_real <= _zz_6122[17 : 0];
    data_mid_4_1_imag <= _zz_6130[17 : 0];
    data_mid_4_10_real <= _zz_6147[17 : 0];
    data_mid_4_10_imag <= _zz_6155[17 : 0];
    data_mid_4_2_real <= _zz_6163[17 : 0];
    data_mid_4_2_imag <= _zz_6171[17 : 0];
    data_mid_4_11_real <= _zz_6188[17 : 0];
    data_mid_4_11_imag <= _zz_6196[17 : 0];
    data_mid_4_3_real <= _zz_6204[17 : 0];
    data_mid_4_3_imag <= _zz_6212[17 : 0];
    data_mid_4_12_real <= _zz_6229[17 : 0];
    data_mid_4_12_imag <= _zz_6237[17 : 0];
    data_mid_4_4_real <= _zz_6245[17 : 0];
    data_mid_4_4_imag <= _zz_6253[17 : 0];
    data_mid_4_13_real <= _zz_6270[17 : 0];
    data_mid_4_13_imag <= _zz_6278[17 : 0];
    data_mid_4_5_real <= _zz_6286[17 : 0];
    data_mid_4_5_imag <= _zz_6294[17 : 0];
    data_mid_4_14_real <= _zz_6311[17 : 0];
    data_mid_4_14_imag <= _zz_6319[17 : 0];
    data_mid_4_6_real <= _zz_6327[17 : 0];
    data_mid_4_6_imag <= _zz_6335[17 : 0];
    data_mid_4_15_real <= _zz_6352[17 : 0];
    data_mid_4_15_imag <= _zz_6360[17 : 0];
    data_mid_4_7_real <= _zz_6368[17 : 0];
    data_mid_4_7_imag <= _zz_6376[17 : 0];
    data_mid_4_24_real <= _zz_6393[17 : 0];
    data_mid_4_24_imag <= _zz_6401[17 : 0];
    data_mid_4_16_real <= _zz_6409[17 : 0];
    data_mid_4_16_imag <= _zz_6417[17 : 0];
    data_mid_4_25_real <= _zz_6434[17 : 0];
    data_mid_4_25_imag <= _zz_6442[17 : 0];
    data_mid_4_17_real <= _zz_6450[17 : 0];
    data_mid_4_17_imag <= _zz_6458[17 : 0];
    data_mid_4_26_real <= _zz_6475[17 : 0];
    data_mid_4_26_imag <= _zz_6483[17 : 0];
    data_mid_4_18_real <= _zz_6491[17 : 0];
    data_mid_4_18_imag <= _zz_6499[17 : 0];
    data_mid_4_27_real <= _zz_6516[17 : 0];
    data_mid_4_27_imag <= _zz_6524[17 : 0];
    data_mid_4_19_real <= _zz_6532[17 : 0];
    data_mid_4_19_imag <= _zz_6540[17 : 0];
    data_mid_4_28_real <= _zz_6557[17 : 0];
    data_mid_4_28_imag <= _zz_6565[17 : 0];
    data_mid_4_20_real <= _zz_6573[17 : 0];
    data_mid_4_20_imag <= _zz_6581[17 : 0];
    data_mid_4_29_real <= _zz_6598[17 : 0];
    data_mid_4_29_imag <= _zz_6606[17 : 0];
    data_mid_4_21_real <= _zz_6614[17 : 0];
    data_mid_4_21_imag <= _zz_6622[17 : 0];
    data_mid_4_30_real <= _zz_6639[17 : 0];
    data_mid_4_30_imag <= _zz_6647[17 : 0];
    data_mid_4_22_real <= _zz_6655[17 : 0];
    data_mid_4_22_imag <= _zz_6663[17 : 0];
    data_mid_4_31_real <= _zz_6680[17 : 0];
    data_mid_4_31_imag <= _zz_6688[17 : 0];
    data_mid_4_23_real <= _zz_6696[17 : 0];
    data_mid_4_23_imag <= _zz_6704[17 : 0];
    data_mid_4_40_real <= _zz_6721[17 : 0];
    data_mid_4_40_imag <= _zz_6729[17 : 0];
    data_mid_4_32_real <= _zz_6737[17 : 0];
    data_mid_4_32_imag <= _zz_6745[17 : 0];
    data_mid_4_41_real <= _zz_6762[17 : 0];
    data_mid_4_41_imag <= _zz_6770[17 : 0];
    data_mid_4_33_real <= _zz_6778[17 : 0];
    data_mid_4_33_imag <= _zz_6786[17 : 0];
    data_mid_4_42_real <= _zz_6803[17 : 0];
    data_mid_4_42_imag <= _zz_6811[17 : 0];
    data_mid_4_34_real <= _zz_6819[17 : 0];
    data_mid_4_34_imag <= _zz_6827[17 : 0];
    data_mid_4_43_real <= _zz_6844[17 : 0];
    data_mid_4_43_imag <= _zz_6852[17 : 0];
    data_mid_4_35_real <= _zz_6860[17 : 0];
    data_mid_4_35_imag <= _zz_6868[17 : 0];
    data_mid_4_44_real <= _zz_6885[17 : 0];
    data_mid_4_44_imag <= _zz_6893[17 : 0];
    data_mid_4_36_real <= _zz_6901[17 : 0];
    data_mid_4_36_imag <= _zz_6909[17 : 0];
    data_mid_4_45_real <= _zz_6926[17 : 0];
    data_mid_4_45_imag <= _zz_6934[17 : 0];
    data_mid_4_37_real <= _zz_6942[17 : 0];
    data_mid_4_37_imag <= _zz_6950[17 : 0];
    data_mid_4_46_real <= _zz_6967[17 : 0];
    data_mid_4_46_imag <= _zz_6975[17 : 0];
    data_mid_4_38_real <= _zz_6983[17 : 0];
    data_mid_4_38_imag <= _zz_6991[17 : 0];
    data_mid_4_47_real <= _zz_7008[17 : 0];
    data_mid_4_47_imag <= _zz_7016[17 : 0];
    data_mid_4_39_real <= _zz_7024[17 : 0];
    data_mid_4_39_imag <= _zz_7032[17 : 0];
    data_mid_4_56_real <= _zz_7049[17 : 0];
    data_mid_4_56_imag <= _zz_7057[17 : 0];
    data_mid_4_48_real <= _zz_7065[17 : 0];
    data_mid_4_48_imag <= _zz_7073[17 : 0];
    data_mid_4_57_real <= _zz_7090[17 : 0];
    data_mid_4_57_imag <= _zz_7098[17 : 0];
    data_mid_4_49_real <= _zz_7106[17 : 0];
    data_mid_4_49_imag <= _zz_7114[17 : 0];
    data_mid_4_58_real <= _zz_7131[17 : 0];
    data_mid_4_58_imag <= _zz_7139[17 : 0];
    data_mid_4_50_real <= _zz_7147[17 : 0];
    data_mid_4_50_imag <= _zz_7155[17 : 0];
    data_mid_4_59_real <= _zz_7172[17 : 0];
    data_mid_4_59_imag <= _zz_7180[17 : 0];
    data_mid_4_51_real <= _zz_7188[17 : 0];
    data_mid_4_51_imag <= _zz_7196[17 : 0];
    data_mid_4_60_real <= _zz_7213[17 : 0];
    data_mid_4_60_imag <= _zz_7221[17 : 0];
    data_mid_4_52_real <= _zz_7229[17 : 0];
    data_mid_4_52_imag <= _zz_7237[17 : 0];
    data_mid_4_61_real <= _zz_7254[17 : 0];
    data_mid_4_61_imag <= _zz_7262[17 : 0];
    data_mid_4_53_real <= _zz_7270[17 : 0];
    data_mid_4_53_imag <= _zz_7278[17 : 0];
    data_mid_4_62_real <= _zz_7295[17 : 0];
    data_mid_4_62_imag <= _zz_7303[17 : 0];
    data_mid_4_54_real <= _zz_7311[17 : 0];
    data_mid_4_54_imag <= _zz_7319[17 : 0];
    data_mid_4_63_real <= _zz_7336[17 : 0];
    data_mid_4_63_imag <= _zz_7344[17 : 0];
    data_mid_4_55_real <= _zz_7352[17 : 0];
    data_mid_4_55_imag <= _zz_7360[17 : 0];
    data_mid_5_16_real <= _zz_7377[17 : 0];
    data_mid_5_16_imag <= _zz_7385[17 : 0];
    data_mid_5_0_real <= _zz_7393[17 : 0];
    data_mid_5_0_imag <= _zz_7401[17 : 0];
    data_mid_5_17_real <= _zz_7418[17 : 0];
    data_mid_5_17_imag <= _zz_7426[17 : 0];
    data_mid_5_1_real <= _zz_7434[17 : 0];
    data_mid_5_1_imag <= _zz_7442[17 : 0];
    data_mid_5_18_real <= _zz_7459[17 : 0];
    data_mid_5_18_imag <= _zz_7467[17 : 0];
    data_mid_5_2_real <= _zz_7475[17 : 0];
    data_mid_5_2_imag <= _zz_7483[17 : 0];
    data_mid_5_19_real <= _zz_7500[17 : 0];
    data_mid_5_19_imag <= _zz_7508[17 : 0];
    data_mid_5_3_real <= _zz_7516[17 : 0];
    data_mid_5_3_imag <= _zz_7524[17 : 0];
    data_mid_5_20_real <= _zz_7541[17 : 0];
    data_mid_5_20_imag <= _zz_7549[17 : 0];
    data_mid_5_4_real <= _zz_7557[17 : 0];
    data_mid_5_4_imag <= _zz_7565[17 : 0];
    data_mid_5_21_real <= _zz_7582[17 : 0];
    data_mid_5_21_imag <= _zz_7590[17 : 0];
    data_mid_5_5_real <= _zz_7598[17 : 0];
    data_mid_5_5_imag <= _zz_7606[17 : 0];
    data_mid_5_22_real <= _zz_7623[17 : 0];
    data_mid_5_22_imag <= _zz_7631[17 : 0];
    data_mid_5_6_real <= _zz_7639[17 : 0];
    data_mid_5_6_imag <= _zz_7647[17 : 0];
    data_mid_5_23_real <= _zz_7664[17 : 0];
    data_mid_5_23_imag <= _zz_7672[17 : 0];
    data_mid_5_7_real <= _zz_7680[17 : 0];
    data_mid_5_7_imag <= _zz_7688[17 : 0];
    data_mid_5_24_real <= _zz_7705[17 : 0];
    data_mid_5_24_imag <= _zz_7713[17 : 0];
    data_mid_5_8_real <= _zz_7721[17 : 0];
    data_mid_5_8_imag <= _zz_7729[17 : 0];
    data_mid_5_25_real <= _zz_7746[17 : 0];
    data_mid_5_25_imag <= _zz_7754[17 : 0];
    data_mid_5_9_real <= _zz_7762[17 : 0];
    data_mid_5_9_imag <= _zz_7770[17 : 0];
    data_mid_5_26_real <= _zz_7787[17 : 0];
    data_mid_5_26_imag <= _zz_7795[17 : 0];
    data_mid_5_10_real <= _zz_7803[17 : 0];
    data_mid_5_10_imag <= _zz_7811[17 : 0];
    data_mid_5_27_real <= _zz_7828[17 : 0];
    data_mid_5_27_imag <= _zz_7836[17 : 0];
    data_mid_5_11_real <= _zz_7844[17 : 0];
    data_mid_5_11_imag <= _zz_7852[17 : 0];
    data_mid_5_28_real <= _zz_7869[17 : 0];
    data_mid_5_28_imag <= _zz_7877[17 : 0];
    data_mid_5_12_real <= _zz_7885[17 : 0];
    data_mid_5_12_imag <= _zz_7893[17 : 0];
    data_mid_5_29_real <= _zz_7910[17 : 0];
    data_mid_5_29_imag <= _zz_7918[17 : 0];
    data_mid_5_13_real <= _zz_7926[17 : 0];
    data_mid_5_13_imag <= _zz_7934[17 : 0];
    data_mid_5_30_real <= _zz_7951[17 : 0];
    data_mid_5_30_imag <= _zz_7959[17 : 0];
    data_mid_5_14_real <= _zz_7967[17 : 0];
    data_mid_5_14_imag <= _zz_7975[17 : 0];
    data_mid_5_31_real <= _zz_7992[17 : 0];
    data_mid_5_31_imag <= _zz_8000[17 : 0];
    data_mid_5_15_real <= _zz_8008[17 : 0];
    data_mid_5_15_imag <= _zz_8016[17 : 0];
    data_mid_5_48_real <= _zz_8033[17 : 0];
    data_mid_5_48_imag <= _zz_8041[17 : 0];
    data_mid_5_32_real <= _zz_8049[17 : 0];
    data_mid_5_32_imag <= _zz_8057[17 : 0];
    data_mid_5_49_real <= _zz_8074[17 : 0];
    data_mid_5_49_imag <= _zz_8082[17 : 0];
    data_mid_5_33_real <= _zz_8090[17 : 0];
    data_mid_5_33_imag <= _zz_8098[17 : 0];
    data_mid_5_50_real <= _zz_8115[17 : 0];
    data_mid_5_50_imag <= _zz_8123[17 : 0];
    data_mid_5_34_real <= _zz_8131[17 : 0];
    data_mid_5_34_imag <= _zz_8139[17 : 0];
    data_mid_5_51_real <= _zz_8156[17 : 0];
    data_mid_5_51_imag <= _zz_8164[17 : 0];
    data_mid_5_35_real <= _zz_8172[17 : 0];
    data_mid_5_35_imag <= _zz_8180[17 : 0];
    data_mid_5_52_real <= _zz_8197[17 : 0];
    data_mid_5_52_imag <= _zz_8205[17 : 0];
    data_mid_5_36_real <= _zz_8213[17 : 0];
    data_mid_5_36_imag <= _zz_8221[17 : 0];
    data_mid_5_53_real <= _zz_8238[17 : 0];
    data_mid_5_53_imag <= _zz_8246[17 : 0];
    data_mid_5_37_real <= _zz_8254[17 : 0];
    data_mid_5_37_imag <= _zz_8262[17 : 0];
    data_mid_5_54_real <= _zz_8279[17 : 0];
    data_mid_5_54_imag <= _zz_8287[17 : 0];
    data_mid_5_38_real <= _zz_8295[17 : 0];
    data_mid_5_38_imag <= _zz_8303[17 : 0];
    data_mid_5_55_real <= _zz_8320[17 : 0];
    data_mid_5_55_imag <= _zz_8328[17 : 0];
    data_mid_5_39_real <= _zz_8336[17 : 0];
    data_mid_5_39_imag <= _zz_8344[17 : 0];
    data_mid_5_56_real <= _zz_8361[17 : 0];
    data_mid_5_56_imag <= _zz_8369[17 : 0];
    data_mid_5_40_real <= _zz_8377[17 : 0];
    data_mid_5_40_imag <= _zz_8385[17 : 0];
    data_mid_5_57_real <= _zz_8402[17 : 0];
    data_mid_5_57_imag <= _zz_8410[17 : 0];
    data_mid_5_41_real <= _zz_8418[17 : 0];
    data_mid_5_41_imag <= _zz_8426[17 : 0];
    data_mid_5_58_real <= _zz_8443[17 : 0];
    data_mid_5_58_imag <= _zz_8451[17 : 0];
    data_mid_5_42_real <= _zz_8459[17 : 0];
    data_mid_5_42_imag <= _zz_8467[17 : 0];
    data_mid_5_59_real <= _zz_8484[17 : 0];
    data_mid_5_59_imag <= _zz_8492[17 : 0];
    data_mid_5_43_real <= _zz_8500[17 : 0];
    data_mid_5_43_imag <= _zz_8508[17 : 0];
    data_mid_5_60_real <= _zz_8525[17 : 0];
    data_mid_5_60_imag <= _zz_8533[17 : 0];
    data_mid_5_44_real <= _zz_8541[17 : 0];
    data_mid_5_44_imag <= _zz_8549[17 : 0];
    data_mid_5_61_real <= _zz_8566[17 : 0];
    data_mid_5_61_imag <= _zz_8574[17 : 0];
    data_mid_5_45_real <= _zz_8582[17 : 0];
    data_mid_5_45_imag <= _zz_8590[17 : 0];
    data_mid_5_62_real <= _zz_8607[17 : 0];
    data_mid_5_62_imag <= _zz_8615[17 : 0];
    data_mid_5_46_real <= _zz_8623[17 : 0];
    data_mid_5_46_imag <= _zz_8631[17 : 0];
    data_mid_5_63_real <= _zz_8648[17 : 0];
    data_mid_5_63_imag <= _zz_8656[17 : 0];
    data_mid_5_47_real <= _zz_8664[17 : 0];
    data_mid_5_47_imag <= _zz_8672[17 : 0];
    data_mid_6_32_real <= _zz_8689[17 : 0];
    data_mid_6_32_imag <= _zz_8697[17 : 0];
    data_mid_6_0_real <= _zz_8705[17 : 0];
    data_mid_6_0_imag <= _zz_8713[17 : 0];
    data_mid_6_33_real <= _zz_8730[17 : 0];
    data_mid_6_33_imag <= _zz_8738[17 : 0];
    data_mid_6_1_real <= _zz_8746[17 : 0];
    data_mid_6_1_imag <= _zz_8754[17 : 0];
    data_mid_6_34_real <= _zz_8771[17 : 0];
    data_mid_6_34_imag <= _zz_8779[17 : 0];
    data_mid_6_2_real <= _zz_8787[17 : 0];
    data_mid_6_2_imag <= _zz_8795[17 : 0];
    data_mid_6_35_real <= _zz_8812[17 : 0];
    data_mid_6_35_imag <= _zz_8820[17 : 0];
    data_mid_6_3_real <= _zz_8828[17 : 0];
    data_mid_6_3_imag <= _zz_8836[17 : 0];
    data_mid_6_36_real <= _zz_8853[17 : 0];
    data_mid_6_36_imag <= _zz_8861[17 : 0];
    data_mid_6_4_real <= _zz_8869[17 : 0];
    data_mid_6_4_imag <= _zz_8877[17 : 0];
    data_mid_6_37_real <= _zz_8894[17 : 0];
    data_mid_6_37_imag <= _zz_8902[17 : 0];
    data_mid_6_5_real <= _zz_8910[17 : 0];
    data_mid_6_5_imag <= _zz_8918[17 : 0];
    data_mid_6_38_real <= _zz_8935[17 : 0];
    data_mid_6_38_imag <= _zz_8943[17 : 0];
    data_mid_6_6_real <= _zz_8951[17 : 0];
    data_mid_6_6_imag <= _zz_8959[17 : 0];
    data_mid_6_39_real <= _zz_8976[17 : 0];
    data_mid_6_39_imag <= _zz_8984[17 : 0];
    data_mid_6_7_real <= _zz_8992[17 : 0];
    data_mid_6_7_imag <= _zz_9000[17 : 0];
    data_mid_6_40_real <= _zz_9017[17 : 0];
    data_mid_6_40_imag <= _zz_9025[17 : 0];
    data_mid_6_8_real <= _zz_9033[17 : 0];
    data_mid_6_8_imag <= _zz_9041[17 : 0];
    data_mid_6_41_real <= _zz_9058[17 : 0];
    data_mid_6_41_imag <= _zz_9066[17 : 0];
    data_mid_6_9_real <= _zz_9074[17 : 0];
    data_mid_6_9_imag <= _zz_9082[17 : 0];
    data_mid_6_42_real <= _zz_9099[17 : 0];
    data_mid_6_42_imag <= _zz_9107[17 : 0];
    data_mid_6_10_real <= _zz_9115[17 : 0];
    data_mid_6_10_imag <= _zz_9123[17 : 0];
    data_mid_6_43_real <= _zz_9140[17 : 0];
    data_mid_6_43_imag <= _zz_9148[17 : 0];
    data_mid_6_11_real <= _zz_9156[17 : 0];
    data_mid_6_11_imag <= _zz_9164[17 : 0];
    data_mid_6_44_real <= _zz_9181[17 : 0];
    data_mid_6_44_imag <= _zz_9189[17 : 0];
    data_mid_6_12_real <= _zz_9197[17 : 0];
    data_mid_6_12_imag <= _zz_9205[17 : 0];
    data_mid_6_45_real <= _zz_9222[17 : 0];
    data_mid_6_45_imag <= _zz_9230[17 : 0];
    data_mid_6_13_real <= _zz_9238[17 : 0];
    data_mid_6_13_imag <= _zz_9246[17 : 0];
    data_mid_6_46_real <= _zz_9263[17 : 0];
    data_mid_6_46_imag <= _zz_9271[17 : 0];
    data_mid_6_14_real <= _zz_9279[17 : 0];
    data_mid_6_14_imag <= _zz_9287[17 : 0];
    data_mid_6_47_real <= _zz_9304[17 : 0];
    data_mid_6_47_imag <= _zz_9312[17 : 0];
    data_mid_6_15_real <= _zz_9320[17 : 0];
    data_mid_6_15_imag <= _zz_9328[17 : 0];
    data_mid_6_48_real <= _zz_9345[17 : 0];
    data_mid_6_48_imag <= _zz_9353[17 : 0];
    data_mid_6_16_real <= _zz_9361[17 : 0];
    data_mid_6_16_imag <= _zz_9369[17 : 0];
    data_mid_6_49_real <= _zz_9386[17 : 0];
    data_mid_6_49_imag <= _zz_9394[17 : 0];
    data_mid_6_17_real <= _zz_9402[17 : 0];
    data_mid_6_17_imag <= _zz_9410[17 : 0];
    data_mid_6_50_real <= _zz_9427[17 : 0];
    data_mid_6_50_imag <= _zz_9435[17 : 0];
    data_mid_6_18_real <= _zz_9443[17 : 0];
    data_mid_6_18_imag <= _zz_9451[17 : 0];
    data_mid_6_51_real <= _zz_9468[17 : 0];
    data_mid_6_51_imag <= _zz_9476[17 : 0];
    data_mid_6_19_real <= _zz_9484[17 : 0];
    data_mid_6_19_imag <= _zz_9492[17 : 0];
    data_mid_6_52_real <= _zz_9509[17 : 0];
    data_mid_6_52_imag <= _zz_9517[17 : 0];
    data_mid_6_20_real <= _zz_9525[17 : 0];
    data_mid_6_20_imag <= _zz_9533[17 : 0];
    data_mid_6_53_real <= _zz_9550[17 : 0];
    data_mid_6_53_imag <= _zz_9558[17 : 0];
    data_mid_6_21_real <= _zz_9566[17 : 0];
    data_mid_6_21_imag <= _zz_9574[17 : 0];
    data_mid_6_54_real <= _zz_9591[17 : 0];
    data_mid_6_54_imag <= _zz_9599[17 : 0];
    data_mid_6_22_real <= _zz_9607[17 : 0];
    data_mid_6_22_imag <= _zz_9615[17 : 0];
    data_mid_6_55_real <= _zz_9632[17 : 0];
    data_mid_6_55_imag <= _zz_9640[17 : 0];
    data_mid_6_23_real <= _zz_9648[17 : 0];
    data_mid_6_23_imag <= _zz_9656[17 : 0];
    data_mid_6_56_real <= _zz_9673[17 : 0];
    data_mid_6_56_imag <= _zz_9681[17 : 0];
    data_mid_6_24_real <= _zz_9689[17 : 0];
    data_mid_6_24_imag <= _zz_9697[17 : 0];
    data_mid_6_57_real <= _zz_9714[17 : 0];
    data_mid_6_57_imag <= _zz_9722[17 : 0];
    data_mid_6_25_real <= _zz_9730[17 : 0];
    data_mid_6_25_imag <= _zz_9738[17 : 0];
    data_mid_6_58_real <= _zz_9755[17 : 0];
    data_mid_6_58_imag <= _zz_9763[17 : 0];
    data_mid_6_26_real <= _zz_9771[17 : 0];
    data_mid_6_26_imag <= _zz_9779[17 : 0];
    data_mid_6_59_real <= _zz_9796[17 : 0];
    data_mid_6_59_imag <= _zz_9804[17 : 0];
    data_mid_6_27_real <= _zz_9812[17 : 0];
    data_mid_6_27_imag <= _zz_9820[17 : 0];
    data_mid_6_60_real <= _zz_9837[17 : 0];
    data_mid_6_60_imag <= _zz_9845[17 : 0];
    data_mid_6_28_real <= _zz_9853[17 : 0];
    data_mid_6_28_imag <= _zz_9861[17 : 0];
    data_mid_6_61_real <= _zz_9878[17 : 0];
    data_mid_6_61_imag <= _zz_9886[17 : 0];
    data_mid_6_29_real <= _zz_9894[17 : 0];
    data_mid_6_29_imag <= _zz_9902[17 : 0];
    data_mid_6_62_real <= _zz_9919[17 : 0];
    data_mid_6_62_imag <= _zz_9927[17 : 0];
    data_mid_6_30_real <= _zz_9935[17 : 0];
    data_mid_6_30_imag <= _zz_9943[17 : 0];
    data_mid_6_63_real <= _zz_9960[17 : 0];
    data_mid_6_63_imag <= _zz_9968[17 : 0];
    data_mid_6_31_real <= _zz_9976[17 : 0];
    data_mid_6_31_imag <= _zz_9984[17 : 0];
  end

  always @ (posedge clk or posedge reset) begin
    if (reset) begin
      io_data_in_valid_delay_1 <= 1'b0;
      io_data_in_valid_delay_2 <= 1'b0;
      io_data_in_valid_delay_3 <= 1'b0;
      io_data_in_valid_delay_4 <= 1'b0;
      io_data_in_valid_delay_5 <= 1'b0;
      io_data_in_valid_delay_6 <= 1'b0;
      io_data_in_valid_delay_7 <= 1'b0;
      io_data_in_valid_delay_8 <= 1'b0;
    end else begin
      io_data_in_valid_delay_1 <= io_data_in_valid;
      io_data_in_valid_delay_2 <= io_data_in_valid_delay_1;
      io_data_in_valid_delay_3 <= io_data_in_valid_delay_2;
      io_data_in_valid_delay_4 <= io_data_in_valid_delay_3;
      io_data_in_valid_delay_5 <= io_data_in_valid_delay_4;
      io_data_in_valid_delay_6 <= io_data_in_valid_delay_5;
      io_data_in_valid_delay_7 <= io_data_in_valid_delay_6;
      io_data_in_valid_delay_8 <= io_data_in_valid_delay_7;
    end
  end


endmodule

module MyFFT (
  input               io_data_in_valid,
  input      [17:0]   io_data_in_payload_0_real,
  input      [17:0]   io_data_in_payload_0_imag,
  input      [17:0]   io_data_in_payload_1_real,
  input      [17:0]   io_data_in_payload_1_imag,
  input      [17:0]   io_data_in_payload_2_real,
  input      [17:0]   io_data_in_payload_2_imag,
  input      [17:0]   io_data_in_payload_3_real,
  input      [17:0]   io_data_in_payload_3_imag,
  input      [17:0]   io_data_in_payload_4_real,
  input      [17:0]   io_data_in_payload_4_imag,
  input      [17:0]   io_data_in_payload_5_real,
  input      [17:0]   io_data_in_payload_5_imag,
  input      [17:0]   io_data_in_payload_6_real,
  input      [17:0]   io_data_in_payload_6_imag,
  input      [17:0]   io_data_in_payload_7_real,
  input      [17:0]   io_data_in_payload_7_imag,
  input      [17:0]   io_data_in_payload_8_real,
  input      [17:0]   io_data_in_payload_8_imag,
  input      [17:0]   io_data_in_payload_9_real,
  input      [17:0]   io_data_in_payload_9_imag,
  input      [17:0]   io_data_in_payload_10_real,
  input      [17:0]   io_data_in_payload_10_imag,
  input      [17:0]   io_data_in_payload_11_real,
  input      [17:0]   io_data_in_payload_11_imag,
  input      [17:0]   io_data_in_payload_12_real,
  input      [17:0]   io_data_in_payload_12_imag,
  input      [17:0]   io_data_in_payload_13_real,
  input      [17:0]   io_data_in_payload_13_imag,
  input      [17:0]   io_data_in_payload_14_real,
  input      [17:0]   io_data_in_payload_14_imag,
  input      [17:0]   io_data_in_payload_15_real,
  input      [17:0]   io_data_in_payload_15_imag,
  input      [17:0]   io_data_in_payload_16_real,
  input      [17:0]   io_data_in_payload_16_imag,
  input      [17:0]   io_data_in_payload_17_real,
  input      [17:0]   io_data_in_payload_17_imag,
  input      [17:0]   io_data_in_payload_18_real,
  input      [17:0]   io_data_in_payload_18_imag,
  input      [17:0]   io_data_in_payload_19_real,
  input      [17:0]   io_data_in_payload_19_imag,
  input      [17:0]   io_data_in_payload_20_real,
  input      [17:0]   io_data_in_payload_20_imag,
  input      [17:0]   io_data_in_payload_21_real,
  input      [17:0]   io_data_in_payload_21_imag,
  input      [17:0]   io_data_in_payload_22_real,
  input      [17:0]   io_data_in_payload_22_imag,
  input      [17:0]   io_data_in_payload_23_real,
  input      [17:0]   io_data_in_payload_23_imag,
  input      [17:0]   io_data_in_payload_24_real,
  input      [17:0]   io_data_in_payload_24_imag,
  input      [17:0]   io_data_in_payload_25_real,
  input      [17:0]   io_data_in_payload_25_imag,
  input      [17:0]   io_data_in_payload_26_real,
  input      [17:0]   io_data_in_payload_26_imag,
  input      [17:0]   io_data_in_payload_27_real,
  input      [17:0]   io_data_in_payload_27_imag,
  input      [17:0]   io_data_in_payload_28_real,
  input      [17:0]   io_data_in_payload_28_imag,
  input      [17:0]   io_data_in_payload_29_real,
  input      [17:0]   io_data_in_payload_29_imag,
  input      [17:0]   io_data_in_payload_30_real,
  input      [17:0]   io_data_in_payload_30_imag,
  input      [17:0]   io_data_in_payload_31_real,
  input      [17:0]   io_data_in_payload_31_imag,
  input      [17:0]   io_data_in_payload_32_real,
  input      [17:0]   io_data_in_payload_32_imag,
  input      [17:0]   io_data_in_payload_33_real,
  input      [17:0]   io_data_in_payload_33_imag,
  input      [17:0]   io_data_in_payload_34_real,
  input      [17:0]   io_data_in_payload_34_imag,
  input      [17:0]   io_data_in_payload_35_real,
  input      [17:0]   io_data_in_payload_35_imag,
  input      [17:0]   io_data_in_payload_36_real,
  input      [17:0]   io_data_in_payload_36_imag,
  input      [17:0]   io_data_in_payload_37_real,
  input      [17:0]   io_data_in_payload_37_imag,
  input      [17:0]   io_data_in_payload_38_real,
  input      [17:0]   io_data_in_payload_38_imag,
  input      [17:0]   io_data_in_payload_39_real,
  input      [17:0]   io_data_in_payload_39_imag,
  input      [17:0]   io_data_in_payload_40_real,
  input      [17:0]   io_data_in_payload_40_imag,
  input      [17:0]   io_data_in_payload_41_real,
  input      [17:0]   io_data_in_payload_41_imag,
  input      [17:0]   io_data_in_payload_42_real,
  input      [17:0]   io_data_in_payload_42_imag,
  input      [17:0]   io_data_in_payload_43_real,
  input      [17:0]   io_data_in_payload_43_imag,
  input      [17:0]   io_data_in_payload_44_real,
  input      [17:0]   io_data_in_payload_44_imag,
  input      [17:0]   io_data_in_payload_45_real,
  input      [17:0]   io_data_in_payload_45_imag,
  input      [17:0]   io_data_in_payload_46_real,
  input      [17:0]   io_data_in_payload_46_imag,
  input      [17:0]   io_data_in_payload_47_real,
  input      [17:0]   io_data_in_payload_47_imag,
  input      [17:0]   io_data_in_payload_48_real,
  input      [17:0]   io_data_in_payload_48_imag,
  input      [17:0]   io_data_in_payload_49_real,
  input      [17:0]   io_data_in_payload_49_imag,
  input      [17:0]   io_data_in_payload_50_real,
  input      [17:0]   io_data_in_payload_50_imag,
  input      [17:0]   io_data_in_payload_51_real,
  input      [17:0]   io_data_in_payload_51_imag,
  input      [17:0]   io_data_in_payload_52_real,
  input      [17:0]   io_data_in_payload_52_imag,
  input      [17:0]   io_data_in_payload_53_real,
  input      [17:0]   io_data_in_payload_53_imag,
  input      [17:0]   io_data_in_payload_54_real,
  input      [17:0]   io_data_in_payload_54_imag,
  input      [17:0]   io_data_in_payload_55_real,
  input      [17:0]   io_data_in_payload_55_imag,
  input      [17:0]   io_data_in_payload_56_real,
  input      [17:0]   io_data_in_payload_56_imag,
  input      [17:0]   io_data_in_payload_57_real,
  input      [17:0]   io_data_in_payload_57_imag,
  input      [17:0]   io_data_in_payload_58_real,
  input      [17:0]   io_data_in_payload_58_imag,
  input      [17:0]   io_data_in_payload_59_real,
  input      [17:0]   io_data_in_payload_59_imag,
  input      [17:0]   io_data_in_payload_60_real,
  input      [17:0]   io_data_in_payload_60_imag,
  input      [17:0]   io_data_in_payload_61_real,
  input      [17:0]   io_data_in_payload_61_imag,
  input      [17:0]   io_data_in_payload_62_real,
  input      [17:0]   io_data_in_payload_62_imag,
  input      [17:0]   io_data_in_payload_63_real,
  input      [17:0]   io_data_in_payload_63_imag,
  output              fft_row_valid,
  output     [17:0]   fft_row_payload_0_real,
  output     [17:0]   fft_row_payload_0_imag,
  output     [17:0]   fft_row_payload_1_real,
  output     [17:0]   fft_row_payload_1_imag,
  output     [17:0]   fft_row_payload_2_real,
  output     [17:0]   fft_row_payload_2_imag,
  output     [17:0]   fft_row_payload_3_real,
  output     [17:0]   fft_row_payload_3_imag,
  output     [17:0]   fft_row_payload_4_real,
  output     [17:0]   fft_row_payload_4_imag,
  output     [17:0]   fft_row_payload_5_real,
  output     [17:0]   fft_row_payload_5_imag,
  output     [17:0]   fft_row_payload_6_real,
  output     [17:0]   fft_row_payload_6_imag,
  output     [17:0]   fft_row_payload_7_real,
  output     [17:0]   fft_row_payload_7_imag,
  output     [17:0]   fft_row_payload_8_real,
  output     [17:0]   fft_row_payload_8_imag,
  output     [17:0]   fft_row_payload_9_real,
  output     [17:0]   fft_row_payload_9_imag,
  output     [17:0]   fft_row_payload_10_real,
  output     [17:0]   fft_row_payload_10_imag,
  output     [17:0]   fft_row_payload_11_real,
  output     [17:0]   fft_row_payload_11_imag,
  output     [17:0]   fft_row_payload_12_real,
  output     [17:0]   fft_row_payload_12_imag,
  output     [17:0]   fft_row_payload_13_real,
  output     [17:0]   fft_row_payload_13_imag,
  output     [17:0]   fft_row_payload_14_real,
  output     [17:0]   fft_row_payload_14_imag,
  output     [17:0]   fft_row_payload_15_real,
  output     [17:0]   fft_row_payload_15_imag,
  output     [17:0]   fft_row_payload_16_real,
  output     [17:0]   fft_row_payload_16_imag,
  output     [17:0]   fft_row_payload_17_real,
  output     [17:0]   fft_row_payload_17_imag,
  output     [17:0]   fft_row_payload_18_real,
  output     [17:0]   fft_row_payload_18_imag,
  output     [17:0]   fft_row_payload_19_real,
  output     [17:0]   fft_row_payload_19_imag,
  output     [17:0]   fft_row_payload_20_real,
  output     [17:0]   fft_row_payload_20_imag,
  output     [17:0]   fft_row_payload_21_real,
  output     [17:0]   fft_row_payload_21_imag,
  output     [17:0]   fft_row_payload_22_real,
  output     [17:0]   fft_row_payload_22_imag,
  output     [17:0]   fft_row_payload_23_real,
  output     [17:0]   fft_row_payload_23_imag,
  output     [17:0]   fft_row_payload_24_real,
  output     [17:0]   fft_row_payload_24_imag,
  output     [17:0]   fft_row_payload_25_real,
  output     [17:0]   fft_row_payload_25_imag,
  output     [17:0]   fft_row_payload_26_real,
  output     [17:0]   fft_row_payload_26_imag,
  output     [17:0]   fft_row_payload_27_real,
  output     [17:0]   fft_row_payload_27_imag,
  output     [17:0]   fft_row_payload_28_real,
  output     [17:0]   fft_row_payload_28_imag,
  output     [17:0]   fft_row_payload_29_real,
  output     [17:0]   fft_row_payload_29_imag,
  output     [17:0]   fft_row_payload_30_real,
  output     [17:0]   fft_row_payload_30_imag,
  output     [17:0]   fft_row_payload_31_real,
  output     [17:0]   fft_row_payload_31_imag,
  output     [17:0]   fft_row_payload_32_real,
  output     [17:0]   fft_row_payload_32_imag,
  output     [17:0]   fft_row_payload_33_real,
  output     [17:0]   fft_row_payload_33_imag,
  output     [17:0]   fft_row_payload_34_real,
  output     [17:0]   fft_row_payload_34_imag,
  output     [17:0]   fft_row_payload_35_real,
  output     [17:0]   fft_row_payload_35_imag,
  output     [17:0]   fft_row_payload_36_real,
  output     [17:0]   fft_row_payload_36_imag,
  output     [17:0]   fft_row_payload_37_real,
  output     [17:0]   fft_row_payload_37_imag,
  output     [17:0]   fft_row_payload_38_real,
  output     [17:0]   fft_row_payload_38_imag,
  output     [17:0]   fft_row_payload_39_real,
  output     [17:0]   fft_row_payload_39_imag,
  output     [17:0]   fft_row_payload_40_real,
  output     [17:0]   fft_row_payload_40_imag,
  output     [17:0]   fft_row_payload_41_real,
  output     [17:0]   fft_row_payload_41_imag,
  output     [17:0]   fft_row_payload_42_real,
  output     [17:0]   fft_row_payload_42_imag,
  output     [17:0]   fft_row_payload_43_real,
  output     [17:0]   fft_row_payload_43_imag,
  output     [17:0]   fft_row_payload_44_real,
  output     [17:0]   fft_row_payload_44_imag,
  output     [17:0]   fft_row_payload_45_real,
  output     [17:0]   fft_row_payload_45_imag,
  output     [17:0]   fft_row_payload_46_real,
  output     [17:0]   fft_row_payload_46_imag,
  output     [17:0]   fft_row_payload_47_real,
  output     [17:0]   fft_row_payload_47_imag,
  output     [17:0]   fft_row_payload_48_real,
  output     [17:0]   fft_row_payload_48_imag,
  output     [17:0]   fft_row_payload_49_real,
  output     [17:0]   fft_row_payload_49_imag,
  output     [17:0]   fft_row_payload_50_real,
  output     [17:0]   fft_row_payload_50_imag,
  output     [17:0]   fft_row_payload_51_real,
  output     [17:0]   fft_row_payload_51_imag,
  output     [17:0]   fft_row_payload_52_real,
  output     [17:0]   fft_row_payload_52_imag,
  output     [17:0]   fft_row_payload_53_real,
  output     [17:0]   fft_row_payload_53_imag,
  output     [17:0]   fft_row_payload_54_real,
  output     [17:0]   fft_row_payload_54_imag,
  output     [17:0]   fft_row_payload_55_real,
  output     [17:0]   fft_row_payload_55_imag,
  output     [17:0]   fft_row_payload_56_real,
  output     [17:0]   fft_row_payload_56_imag,
  output     [17:0]   fft_row_payload_57_real,
  output     [17:0]   fft_row_payload_57_imag,
  output     [17:0]   fft_row_payload_58_real,
  output     [17:0]   fft_row_payload_58_imag,
  output     [17:0]   fft_row_payload_59_real,
  output     [17:0]   fft_row_payload_59_imag,
  output     [17:0]   fft_row_payload_60_real,
  output     [17:0]   fft_row_payload_60_imag,
  output     [17:0]   fft_row_payload_61_real,
  output     [17:0]   fft_row_payload_61_imag,
  output     [17:0]   fft_row_payload_62_real,
  output     [17:0]   fft_row_payload_62_imag,
  output     [17:0]   fft_row_payload_63_real,
  output     [17:0]   fft_row_payload_63_imag,
  input               clk,
  input               reset
);
  wire       [35:0]   _zz_961;
  wire       [35:0]   _zz_962;
  wire       [35:0]   _zz_963;
  wire       [35:0]   _zz_964;
  wire       [35:0]   _zz_965;
  wire       [35:0]   _zz_966;
  wire       [35:0]   _zz_967;
  wire       [35:0]   _zz_968;
  wire       [35:0]   _zz_969;
  wire       [35:0]   _zz_970;
  wire       [35:0]   _zz_971;
  wire       [35:0]   _zz_972;
  wire       [35:0]   _zz_973;
  wire       [35:0]   _zz_974;
  wire       [35:0]   _zz_975;
  wire       [35:0]   _zz_976;
  wire       [35:0]   _zz_977;
  wire       [35:0]   _zz_978;
  wire       [35:0]   _zz_979;
  wire       [35:0]   _zz_980;
  wire       [35:0]   _zz_981;
  wire       [35:0]   _zz_982;
  wire       [35:0]   _zz_983;
  wire       [35:0]   _zz_984;
  wire       [35:0]   _zz_985;
  wire       [35:0]   _zz_986;
  wire       [35:0]   _zz_987;
  wire       [35:0]   _zz_988;
  wire       [35:0]   _zz_989;
  wire       [35:0]   _zz_990;
  wire       [35:0]   _zz_991;
  wire       [35:0]   _zz_992;
  wire       [35:0]   _zz_993;
  wire       [35:0]   _zz_994;
  wire       [35:0]   _zz_995;
  wire       [35:0]   _zz_996;
  wire       [35:0]   _zz_997;
  wire       [35:0]   _zz_998;
  wire       [35:0]   _zz_999;
  wire       [35:0]   _zz_1000;
  wire       [35:0]   _zz_1001;
  wire       [35:0]   _zz_1002;
  wire       [35:0]   _zz_1003;
  wire       [35:0]   _zz_1004;
  wire       [35:0]   _zz_1005;
  wire       [35:0]   _zz_1006;
  wire       [35:0]   _zz_1007;
  wire       [35:0]   _zz_1008;
  wire       [35:0]   _zz_1009;
  wire       [35:0]   _zz_1010;
  wire       [35:0]   _zz_1011;
  wire       [35:0]   _zz_1012;
  wire       [35:0]   _zz_1013;
  wire       [35:0]   _zz_1014;
  wire       [35:0]   _zz_1015;
  wire       [35:0]   _zz_1016;
  wire       [35:0]   _zz_1017;
  wire       [35:0]   _zz_1018;
  wire       [35:0]   _zz_1019;
  wire       [35:0]   _zz_1020;
  wire       [35:0]   _zz_1021;
  wire       [35:0]   _zz_1022;
  wire       [35:0]   _zz_1023;
  wire       [35:0]   _zz_1024;
  wire       [35:0]   _zz_1025;
  wire       [35:0]   _zz_1026;
  wire       [35:0]   _zz_1027;
  wire       [35:0]   _zz_1028;
  wire       [35:0]   _zz_1029;
  wire       [35:0]   _zz_1030;
  wire       [35:0]   _zz_1031;
  wire       [35:0]   _zz_1032;
  wire       [35:0]   _zz_1033;
  wire       [35:0]   _zz_1034;
  wire       [35:0]   _zz_1035;
  wire       [35:0]   _zz_1036;
  wire       [35:0]   _zz_1037;
  wire       [35:0]   _zz_1038;
  wire       [35:0]   _zz_1039;
  wire       [35:0]   _zz_1040;
  wire       [35:0]   _zz_1041;
  wire       [35:0]   _zz_1042;
  wire       [35:0]   _zz_1043;
  wire       [35:0]   _zz_1044;
  wire       [35:0]   _zz_1045;
  wire       [35:0]   _zz_1046;
  wire       [35:0]   _zz_1047;
  wire       [35:0]   _zz_1048;
  wire       [35:0]   _zz_1049;
  wire       [35:0]   _zz_1050;
  wire       [35:0]   _zz_1051;
  wire       [35:0]   _zz_1052;
  wire       [35:0]   _zz_1053;
  wire       [35:0]   _zz_1054;
  wire       [35:0]   _zz_1055;
  wire       [35:0]   _zz_1056;
  wire       [35:0]   _zz_1057;
  wire       [35:0]   _zz_1058;
  wire       [35:0]   _zz_1059;
  wire       [35:0]   _zz_1060;
  wire       [35:0]   _zz_1061;
  wire       [35:0]   _zz_1062;
  wire       [35:0]   _zz_1063;
  wire       [35:0]   _zz_1064;
  wire       [35:0]   _zz_1065;
  wire       [35:0]   _zz_1066;
  wire       [35:0]   _zz_1067;
  wire       [35:0]   _zz_1068;
  wire       [35:0]   _zz_1069;
  wire       [35:0]   _zz_1070;
  wire       [35:0]   _zz_1071;
  wire       [35:0]   _zz_1072;
  wire       [35:0]   _zz_1073;
  wire       [35:0]   _zz_1074;
  wire       [35:0]   _zz_1075;
  wire       [35:0]   _zz_1076;
  wire       [35:0]   _zz_1077;
  wire       [35:0]   _zz_1078;
  wire       [35:0]   _zz_1079;
  wire       [35:0]   _zz_1080;
  wire       [35:0]   _zz_1081;
  wire       [35:0]   _zz_1082;
  wire       [35:0]   _zz_1083;
  wire       [35:0]   _zz_1084;
  wire       [35:0]   _zz_1085;
  wire       [35:0]   _zz_1086;
  wire       [35:0]   _zz_1087;
  wire       [35:0]   _zz_1088;
  wire       [35:0]   _zz_1089;
  wire       [35:0]   _zz_1090;
  wire       [35:0]   _zz_1091;
  wire       [35:0]   _zz_1092;
  wire       [35:0]   _zz_1093;
  wire       [35:0]   _zz_1094;
  wire       [35:0]   _zz_1095;
  wire       [35:0]   _zz_1096;
  wire       [35:0]   _zz_1097;
  wire       [35:0]   _zz_1098;
  wire       [35:0]   _zz_1099;
  wire       [35:0]   _zz_1100;
  wire       [35:0]   _zz_1101;
  wire       [35:0]   _zz_1102;
  wire       [35:0]   _zz_1103;
  wire       [35:0]   _zz_1104;
  wire       [35:0]   _zz_1105;
  wire       [35:0]   _zz_1106;
  wire       [35:0]   _zz_1107;
  wire       [35:0]   _zz_1108;
  wire       [35:0]   _zz_1109;
  wire       [35:0]   _zz_1110;
  wire       [35:0]   _zz_1111;
  wire       [35:0]   _zz_1112;
  wire       [35:0]   _zz_1113;
  wire       [35:0]   _zz_1114;
  wire       [35:0]   _zz_1115;
  wire       [35:0]   _zz_1116;
  wire       [35:0]   _zz_1117;
  wire       [35:0]   _zz_1118;
  wire       [35:0]   _zz_1119;
  wire       [35:0]   _zz_1120;
  wire       [35:0]   _zz_1121;
  wire       [35:0]   _zz_1122;
  wire       [35:0]   _zz_1123;
  wire       [35:0]   _zz_1124;
  wire       [35:0]   _zz_1125;
  wire       [35:0]   _zz_1126;
  wire       [35:0]   _zz_1127;
  wire       [35:0]   _zz_1128;
  wire       [35:0]   _zz_1129;
  wire       [35:0]   _zz_1130;
  wire       [35:0]   _zz_1131;
  wire       [35:0]   _zz_1132;
  wire       [35:0]   _zz_1133;
  wire       [35:0]   _zz_1134;
  wire       [35:0]   _zz_1135;
  wire       [35:0]   _zz_1136;
  wire       [35:0]   _zz_1137;
  wire       [35:0]   _zz_1138;
  wire       [35:0]   _zz_1139;
  wire       [35:0]   _zz_1140;
  wire       [35:0]   _zz_1141;
  wire       [35:0]   _zz_1142;
  wire       [35:0]   _zz_1143;
  wire       [35:0]   _zz_1144;
  wire       [35:0]   _zz_1145;
  wire       [35:0]   _zz_1146;
  wire       [35:0]   _zz_1147;
  wire       [35:0]   _zz_1148;
  wire       [35:0]   _zz_1149;
  wire       [35:0]   _zz_1150;
  wire       [35:0]   _zz_1151;
  wire       [35:0]   _zz_1152;
  wire       [35:0]   _zz_1153;
  wire       [35:0]   _zz_1154;
  wire       [35:0]   _zz_1155;
  wire       [35:0]   _zz_1156;
  wire       [35:0]   _zz_1157;
  wire       [35:0]   _zz_1158;
  wire       [35:0]   _zz_1159;
  wire       [35:0]   _zz_1160;
  wire       [35:0]   _zz_1161;
  wire       [35:0]   _zz_1162;
  wire       [35:0]   _zz_1163;
  wire       [35:0]   _zz_1164;
  wire       [35:0]   _zz_1165;
  wire       [35:0]   _zz_1166;
  wire       [35:0]   _zz_1167;
  wire       [35:0]   _zz_1168;
  wire       [35:0]   _zz_1169;
  wire       [35:0]   _zz_1170;
  wire       [35:0]   _zz_1171;
  wire       [35:0]   _zz_1172;
  wire       [35:0]   _zz_1173;
  wire       [35:0]   _zz_1174;
  wire       [35:0]   _zz_1175;
  wire       [35:0]   _zz_1176;
  wire       [35:0]   _zz_1177;
  wire       [35:0]   _zz_1178;
  wire       [35:0]   _zz_1179;
  wire       [35:0]   _zz_1180;
  wire       [35:0]   _zz_1181;
  wire       [35:0]   _zz_1182;
  wire       [35:0]   _zz_1183;
  wire       [35:0]   _zz_1184;
  wire       [35:0]   _zz_1185;
  wire       [35:0]   _zz_1186;
  wire       [35:0]   _zz_1187;
  wire       [35:0]   _zz_1188;
  wire       [35:0]   _zz_1189;
  wire       [35:0]   _zz_1190;
  wire       [35:0]   _zz_1191;
  wire       [35:0]   _zz_1192;
  wire       [35:0]   _zz_1193;
  wire       [35:0]   _zz_1194;
  wire       [35:0]   _zz_1195;
  wire       [35:0]   _zz_1196;
  wire       [35:0]   _zz_1197;
  wire       [35:0]   _zz_1198;
  wire       [35:0]   _zz_1199;
  wire       [35:0]   _zz_1200;
  wire       [35:0]   _zz_1201;
  wire       [35:0]   _zz_1202;
  wire       [35:0]   _zz_1203;
  wire       [35:0]   _zz_1204;
  wire       [35:0]   _zz_1205;
  wire       [35:0]   _zz_1206;
  wire       [35:0]   _zz_1207;
  wire       [35:0]   _zz_1208;
  wire       [35:0]   _zz_1209;
  wire       [35:0]   _zz_1210;
  wire       [35:0]   _zz_1211;
  wire       [35:0]   _zz_1212;
  wire       [35:0]   _zz_1213;
  wire       [35:0]   _zz_1214;
  wire       [35:0]   _zz_1215;
  wire       [35:0]   _zz_1216;
  wire       [35:0]   _zz_1217;
  wire       [35:0]   _zz_1218;
  wire       [35:0]   _zz_1219;
  wire       [35:0]   _zz_1220;
  wire       [35:0]   _zz_1221;
  wire       [35:0]   _zz_1222;
  wire       [35:0]   _zz_1223;
  wire       [35:0]   _zz_1224;
  wire       [35:0]   _zz_1225;
  wire       [35:0]   _zz_1226;
  wire       [35:0]   _zz_1227;
  wire       [35:0]   _zz_1228;
  wire       [35:0]   _zz_1229;
  wire       [35:0]   _zz_1230;
  wire       [35:0]   _zz_1231;
  wire       [35:0]   _zz_1232;
  wire       [35:0]   _zz_1233;
  wire       [35:0]   _zz_1234;
  wire       [35:0]   _zz_1235;
  wire       [35:0]   _zz_1236;
  wire       [35:0]   _zz_1237;
  wire       [35:0]   _zz_1238;
  wire       [35:0]   _zz_1239;
  wire       [35:0]   _zz_1240;
  wire       [35:0]   _zz_1241;
  wire       [35:0]   _zz_1242;
  wire       [35:0]   _zz_1243;
  wire       [35:0]   _zz_1244;
  wire       [35:0]   _zz_1245;
  wire       [35:0]   _zz_1246;
  wire       [35:0]   _zz_1247;
  wire       [35:0]   _zz_1248;
  wire       [35:0]   _zz_1249;
  wire       [35:0]   _zz_1250;
  wire       [35:0]   _zz_1251;
  wire       [35:0]   _zz_1252;
  wire       [35:0]   _zz_1253;
  wire       [35:0]   _zz_1254;
  wire       [35:0]   _zz_1255;
  wire       [35:0]   _zz_1256;
  wire       [35:0]   _zz_1257;
  wire       [35:0]   _zz_1258;
  wire       [35:0]   _zz_1259;
  wire       [35:0]   _zz_1260;
  wire       [35:0]   _zz_1261;
  wire       [35:0]   _zz_1262;
  wire       [35:0]   _zz_1263;
  wire       [35:0]   _zz_1264;
  wire       [35:0]   _zz_1265;
  wire       [35:0]   _zz_1266;
  wire       [35:0]   _zz_1267;
  wire       [35:0]   _zz_1268;
  wire       [35:0]   _zz_1269;
  wire       [35:0]   _zz_1270;
  wire       [35:0]   _zz_1271;
  wire       [35:0]   _zz_1272;
  wire       [35:0]   _zz_1273;
  wire       [35:0]   _zz_1274;
  wire       [35:0]   _zz_1275;
  wire       [35:0]   _zz_1276;
  wire       [35:0]   _zz_1277;
  wire       [35:0]   _zz_1278;
  wire       [35:0]   _zz_1279;
  wire       [35:0]   _zz_1280;
  wire       [35:0]   _zz_1281;
  wire       [35:0]   _zz_1282;
  wire       [35:0]   _zz_1283;
  wire       [35:0]   _zz_1284;
  wire       [35:0]   _zz_1285;
  wire       [35:0]   _zz_1286;
  wire       [35:0]   _zz_1287;
  wire       [35:0]   _zz_1288;
  wire       [35:0]   _zz_1289;
  wire       [35:0]   _zz_1290;
  wire       [35:0]   _zz_1291;
  wire       [35:0]   _zz_1292;
  wire       [35:0]   _zz_1293;
  wire       [35:0]   _zz_1294;
  wire       [35:0]   _zz_1295;
  wire       [35:0]   _zz_1296;
  wire       [35:0]   _zz_1297;
  wire       [35:0]   _zz_1298;
  wire       [35:0]   _zz_1299;
  wire       [35:0]   _zz_1300;
  wire       [35:0]   _zz_1301;
  wire       [35:0]   _zz_1302;
  wire       [35:0]   _zz_1303;
  wire       [35:0]   _zz_1304;
  wire       [35:0]   _zz_1305;
  wire       [35:0]   _zz_1306;
  wire       [35:0]   _zz_1307;
  wire       [35:0]   _zz_1308;
  wire       [35:0]   _zz_1309;
  wire       [35:0]   _zz_1310;
  wire       [35:0]   _zz_1311;
  wire       [35:0]   _zz_1312;
  wire       [35:0]   _zz_1313;
  wire       [35:0]   _zz_1314;
  wire       [35:0]   _zz_1315;
  wire       [35:0]   _zz_1316;
  wire       [35:0]   _zz_1317;
  wire       [35:0]   _zz_1318;
  wire       [35:0]   _zz_1319;
  wire       [35:0]   _zz_1320;
  wire       [35:0]   _zz_1321;
  wire       [35:0]   _zz_1322;
  wire       [35:0]   _zz_1323;
  wire       [35:0]   _zz_1324;
  wire       [35:0]   _zz_1325;
  wire       [35:0]   _zz_1326;
  wire       [35:0]   _zz_1327;
  wire       [35:0]   _zz_1328;
  wire       [35:0]   _zz_1329;
  wire       [35:0]   _zz_1330;
  wire       [35:0]   _zz_1331;
  wire       [35:0]   _zz_1332;
  wire       [35:0]   _zz_1333;
  wire       [35:0]   _zz_1334;
  wire       [35:0]   _zz_1335;
  wire       [35:0]   _zz_1336;
  wire       [35:0]   _zz_1337;
  wire       [35:0]   _zz_1338;
  wire       [35:0]   _zz_1339;
  wire       [35:0]   _zz_1340;
  wire       [35:0]   _zz_1341;
  wire       [35:0]   _zz_1342;
  wire       [35:0]   _zz_1343;
  wire       [35:0]   _zz_1344;
  wire       [35:0]   _zz_1345;
  wire       [35:0]   _zz_1346;
  wire       [35:0]   _zz_1347;
  wire       [35:0]   _zz_1348;
  wire       [35:0]   _zz_1349;
  wire       [35:0]   _zz_1350;
  wire       [35:0]   _zz_1351;
  wire       [35:0]   _zz_1352;
  wire       [35:0]   _zz_1353;
  wire       [35:0]   _zz_1354;
  wire       [35:0]   _zz_1355;
  wire       [35:0]   _zz_1356;
  wire       [35:0]   _zz_1357;
  wire       [35:0]   _zz_1358;
  wire       [35:0]   _zz_1359;
  wire       [35:0]   _zz_1360;
  wire       [35:0]   _zz_1361;
  wire       [35:0]   _zz_1362;
  wire       [35:0]   _zz_1363;
  wire       [35:0]   _zz_1364;
  wire       [35:0]   _zz_1365;
  wire       [35:0]   _zz_1366;
  wire       [35:0]   _zz_1367;
  wire       [35:0]   _zz_1368;
  wire       [35:0]   _zz_1369;
  wire       [35:0]   _zz_1370;
  wire       [35:0]   _zz_1371;
  wire       [35:0]   _zz_1372;
  wire       [35:0]   _zz_1373;
  wire       [35:0]   _zz_1374;
  wire       [35:0]   _zz_1375;
  wire       [35:0]   _zz_1376;
  wire       [35:0]   _zz_1377;
  wire       [35:0]   _zz_1378;
  wire       [35:0]   _zz_1379;
  wire       [35:0]   _zz_1380;
  wire       [35:0]   _zz_1381;
  wire       [35:0]   _zz_1382;
  wire       [35:0]   _zz_1383;
  wire       [35:0]   _zz_1384;
  wire       [35:0]   _zz_1385;
  wire       [35:0]   _zz_1386;
  wire       [35:0]   _zz_1387;
  wire       [35:0]   _zz_1388;
  wire       [35:0]   _zz_1389;
  wire       [35:0]   _zz_1390;
  wire       [35:0]   _zz_1391;
  wire       [35:0]   _zz_1392;
  wire       [35:0]   _zz_1393;
  wire       [35:0]   _zz_1394;
  wire       [35:0]   _zz_1395;
  wire       [35:0]   _zz_1396;
  wire       [35:0]   _zz_1397;
  wire       [35:0]   _zz_1398;
  wire       [35:0]   _zz_1399;
  wire       [35:0]   _zz_1400;
  wire       [35:0]   _zz_1401;
  wire       [35:0]   _zz_1402;
  wire       [35:0]   _zz_1403;
  wire       [35:0]   _zz_1404;
  wire       [35:0]   _zz_1405;
  wire       [35:0]   _zz_1406;
  wire       [35:0]   _zz_1407;
  wire       [35:0]   _zz_1408;
  wire       [35:0]   _zz_1409;
  wire       [35:0]   _zz_1410;
  wire       [35:0]   _zz_1411;
  wire       [35:0]   _zz_1412;
  wire       [35:0]   _zz_1413;
  wire       [35:0]   _zz_1414;
  wire       [35:0]   _zz_1415;
  wire       [35:0]   _zz_1416;
  wire       [35:0]   _zz_1417;
  wire       [35:0]   _zz_1418;
  wire       [35:0]   _zz_1419;
  wire       [35:0]   _zz_1420;
  wire       [35:0]   _zz_1421;
  wire       [35:0]   _zz_1422;
  wire       [35:0]   _zz_1423;
  wire       [35:0]   _zz_1424;
  wire       [35:0]   _zz_1425;
  wire       [35:0]   _zz_1426;
  wire       [35:0]   _zz_1427;
  wire       [35:0]   _zz_1428;
  wire       [35:0]   _zz_1429;
  wire       [35:0]   _zz_1430;
  wire       [35:0]   _zz_1431;
  wire       [35:0]   _zz_1432;
  wire       [35:0]   _zz_1433;
  wire       [35:0]   _zz_1434;
  wire       [35:0]   _zz_1435;
  wire       [35:0]   _zz_1436;
  wire       [35:0]   _zz_1437;
  wire       [35:0]   _zz_1438;
  wire       [35:0]   _zz_1439;
  wire       [35:0]   _zz_1440;
  wire       [35:0]   _zz_1441;
  wire       [35:0]   _zz_1442;
  wire       [35:0]   _zz_1443;
  wire       [35:0]   _zz_1444;
  wire       [35:0]   _zz_1445;
  wire       [35:0]   _zz_1446;
  wire       [35:0]   _zz_1447;
  wire       [35:0]   _zz_1448;
  wire       [35:0]   _zz_1449;
  wire       [35:0]   _zz_1450;
  wire       [35:0]   _zz_1451;
  wire       [35:0]   _zz_1452;
  wire       [35:0]   _zz_1453;
  wire       [35:0]   _zz_1454;
  wire       [35:0]   _zz_1455;
  wire       [35:0]   _zz_1456;
  wire       [35:0]   _zz_1457;
  wire       [35:0]   _zz_1458;
  wire       [35:0]   _zz_1459;
  wire       [35:0]   _zz_1460;
  wire       [35:0]   _zz_1461;
  wire       [35:0]   _zz_1462;
  wire       [35:0]   _zz_1463;
  wire       [35:0]   _zz_1464;
  wire       [35:0]   _zz_1465;
  wire       [35:0]   _zz_1466;
  wire       [35:0]   _zz_1467;
  wire       [35:0]   _zz_1468;
  wire       [35:0]   _zz_1469;
  wire       [35:0]   _zz_1470;
  wire       [35:0]   _zz_1471;
  wire       [35:0]   _zz_1472;
  wire       [35:0]   _zz_1473;
  wire       [35:0]   _zz_1474;
  wire       [35:0]   _zz_1475;
  wire       [35:0]   _zz_1476;
  wire       [35:0]   _zz_1477;
  wire       [35:0]   _zz_1478;
  wire       [35:0]   _zz_1479;
  wire       [35:0]   _zz_1480;
  wire       [35:0]   _zz_1481;
  wire       [35:0]   _zz_1482;
  wire       [35:0]   _zz_1483;
  wire       [35:0]   _zz_1484;
  wire       [35:0]   _zz_1485;
  wire       [35:0]   _zz_1486;
  wire       [35:0]   _zz_1487;
  wire       [35:0]   _zz_1488;
  wire       [35:0]   _zz_1489;
  wire       [35:0]   _zz_1490;
  wire       [35:0]   _zz_1491;
  wire       [35:0]   _zz_1492;
  wire       [35:0]   _zz_1493;
  wire       [35:0]   _zz_1494;
  wire       [35:0]   _zz_1495;
  wire       [35:0]   _zz_1496;
  wire       [35:0]   _zz_1497;
  wire       [35:0]   _zz_1498;
  wire       [35:0]   _zz_1499;
  wire       [35:0]   _zz_1500;
  wire       [35:0]   _zz_1501;
  wire       [35:0]   _zz_1502;
  wire       [35:0]   _zz_1503;
  wire       [35:0]   _zz_1504;
  wire       [35:0]   _zz_1505;
  wire       [35:0]   _zz_1506;
  wire       [35:0]   _zz_1507;
  wire       [35:0]   _zz_1508;
  wire       [35:0]   _zz_1509;
  wire       [35:0]   _zz_1510;
  wire       [35:0]   _zz_1511;
  wire       [35:0]   _zz_1512;
  wire       [35:0]   _zz_1513;
  wire       [35:0]   _zz_1514;
  wire       [35:0]   _zz_1515;
  wire       [35:0]   _zz_1516;
  wire       [35:0]   _zz_1517;
  wire       [35:0]   _zz_1518;
  wire       [35:0]   _zz_1519;
  wire       [35:0]   _zz_1520;
  wire       [35:0]   _zz_1521;
  wire       [35:0]   _zz_1522;
  wire       [35:0]   _zz_1523;
  wire       [35:0]   _zz_1524;
  wire       [35:0]   _zz_1525;
  wire       [35:0]   _zz_1526;
  wire       [35:0]   _zz_1527;
  wire       [35:0]   _zz_1528;
  wire       [35:0]   _zz_1529;
  wire       [35:0]   _zz_1530;
  wire       [35:0]   _zz_1531;
  wire       [35:0]   _zz_1532;
  wire       [35:0]   _zz_1533;
  wire       [35:0]   _zz_1534;
  wire       [35:0]   _zz_1535;
  wire       [35:0]   _zz_1536;
  wire       [35:0]   _zz_1537;
  wire       [35:0]   _zz_1538;
  wire       [35:0]   _zz_1539;
  wire       [35:0]   _zz_1540;
  wire       [35:0]   _zz_1541;
  wire       [35:0]   _zz_1542;
  wire       [35:0]   _zz_1543;
  wire       [35:0]   _zz_1544;
  wire       [35:0]   _zz_1545;
  wire       [35:0]   _zz_1546;
  wire       [35:0]   _zz_1547;
  wire       [35:0]   _zz_1548;
  wire       [35:0]   _zz_1549;
  wire       [35:0]   _zz_1550;
  wire       [35:0]   _zz_1551;
  wire       [35:0]   _zz_1552;
  wire       [35:0]   _zz_1553;
  wire       [35:0]   _zz_1554;
  wire       [35:0]   _zz_1555;
  wire       [35:0]   _zz_1556;
  wire       [35:0]   _zz_1557;
  wire       [35:0]   _zz_1558;
  wire       [35:0]   _zz_1559;
  wire       [35:0]   _zz_1560;
  wire       [35:0]   _zz_1561;
  wire       [35:0]   _zz_1562;
  wire       [35:0]   _zz_1563;
  wire       [35:0]   _zz_1564;
  wire       [35:0]   _zz_1565;
  wire       [35:0]   _zz_1566;
  wire       [35:0]   _zz_1567;
  wire       [35:0]   _zz_1568;
  wire       [35:0]   _zz_1569;
  wire       [35:0]   _zz_1570;
  wire       [35:0]   _zz_1571;
  wire       [35:0]   _zz_1572;
  wire       [35:0]   _zz_1573;
  wire       [35:0]   _zz_1574;
  wire       [35:0]   _zz_1575;
  wire       [35:0]   _zz_1576;
  wire       [35:0]   _zz_1577;
  wire       [35:0]   _zz_1578;
  wire       [35:0]   _zz_1579;
  wire       [35:0]   _zz_1580;
  wire       [35:0]   _zz_1581;
  wire       [35:0]   _zz_1582;
  wire       [35:0]   _zz_1583;
  wire       [35:0]   _zz_1584;
  wire       [35:0]   _zz_1585;
  wire       [35:0]   _zz_1586;
  wire       [35:0]   _zz_1587;
  wire       [35:0]   _zz_1588;
  wire       [35:0]   _zz_1589;
  wire       [35:0]   _zz_1590;
  wire       [35:0]   _zz_1591;
  wire       [35:0]   _zz_1592;
  wire       [35:0]   _zz_1593;
  wire       [35:0]   _zz_1594;
  wire       [35:0]   _zz_1595;
  wire       [35:0]   _zz_1596;
  wire       [35:0]   _zz_1597;
  wire       [35:0]   _zz_1598;
  wire       [35:0]   _zz_1599;
  wire       [35:0]   _zz_1600;
  wire       [35:0]   _zz_1601;
  wire       [35:0]   _zz_1602;
  wire       [35:0]   _zz_1603;
  wire       [35:0]   _zz_1604;
  wire       [35:0]   _zz_1605;
  wire       [35:0]   _zz_1606;
  wire       [35:0]   _zz_1607;
  wire       [35:0]   _zz_1608;
  wire       [35:0]   _zz_1609;
  wire       [35:0]   _zz_1610;
  wire       [35:0]   _zz_1611;
  wire       [35:0]   _zz_1612;
  wire       [35:0]   _zz_1613;
  wire       [35:0]   _zz_1614;
  wire       [35:0]   _zz_1615;
  wire       [35:0]   _zz_1616;
  wire       [35:0]   _zz_1617;
  wire       [35:0]   _zz_1618;
  wire       [35:0]   _zz_1619;
  wire       [35:0]   _zz_1620;
  wire       [35:0]   _zz_1621;
  wire       [35:0]   _zz_1622;
  wire       [35:0]   _zz_1623;
  wire       [35:0]   _zz_1624;
  wire       [35:0]   _zz_1625;
  wire       [35:0]   _zz_1626;
  wire       [35:0]   _zz_1627;
  wire       [35:0]   _zz_1628;
  wire       [35:0]   _zz_1629;
  wire       [35:0]   _zz_1630;
  wire       [35:0]   _zz_1631;
  wire       [35:0]   _zz_1632;
  wire       [35:0]   _zz_1633;
  wire       [35:0]   _zz_1634;
  wire       [35:0]   _zz_1635;
  wire       [35:0]   _zz_1636;
  wire       [35:0]   _zz_1637;
  wire       [35:0]   _zz_1638;
  wire       [35:0]   _zz_1639;
  wire       [35:0]   _zz_1640;
  wire       [35:0]   _zz_1641;
  wire       [35:0]   _zz_1642;
  wire       [35:0]   _zz_1643;
  wire       [35:0]   _zz_1644;
  wire       [35:0]   _zz_1645;
  wire       [35:0]   _zz_1646;
  wire       [35:0]   _zz_1647;
  wire       [35:0]   _zz_1648;
  wire       [35:0]   _zz_1649;
  wire       [35:0]   _zz_1650;
  wire       [35:0]   _zz_1651;
  wire       [35:0]   _zz_1652;
  wire       [35:0]   _zz_1653;
  wire       [35:0]   _zz_1654;
  wire       [35:0]   _zz_1655;
  wire       [35:0]   _zz_1656;
  wire       [35:0]   _zz_1657;
  wire       [35:0]   _zz_1658;
  wire       [35:0]   _zz_1659;
  wire       [35:0]   _zz_1660;
  wire       [35:0]   _zz_1661;
  wire       [35:0]   _zz_1662;
  wire       [35:0]   _zz_1663;
  wire       [35:0]   _zz_1664;
  wire       [35:0]   _zz_1665;
  wire       [35:0]   _zz_1666;
  wire       [35:0]   _zz_1667;
  wire       [35:0]   _zz_1668;
  wire       [35:0]   _zz_1669;
  wire       [35:0]   _zz_1670;
  wire       [35:0]   _zz_1671;
  wire       [35:0]   _zz_1672;
  wire       [35:0]   _zz_1673;
  wire       [35:0]   _zz_1674;
  wire       [35:0]   _zz_1675;
  wire       [35:0]   _zz_1676;
  wire       [35:0]   _zz_1677;
  wire       [35:0]   _zz_1678;
  wire       [35:0]   _zz_1679;
  wire       [35:0]   _zz_1680;
  wire       [35:0]   _zz_1681;
  wire       [35:0]   _zz_1682;
  wire       [35:0]   _zz_1683;
  wire       [35:0]   _zz_1684;
  wire       [35:0]   _zz_1685;
  wire       [35:0]   _zz_1686;
  wire       [35:0]   _zz_1687;
  wire       [35:0]   _zz_1688;
  wire       [35:0]   _zz_1689;
  wire       [35:0]   _zz_1690;
  wire       [35:0]   _zz_1691;
  wire       [35:0]   _zz_1692;
  wire       [35:0]   _zz_1693;
  wire       [35:0]   _zz_1694;
  wire       [35:0]   _zz_1695;
  wire       [35:0]   _zz_1696;
  wire       [35:0]   _zz_1697;
  wire       [35:0]   _zz_1698;
  wire       [35:0]   _zz_1699;
  wire       [35:0]   _zz_1700;
  wire       [35:0]   _zz_1701;
  wire       [35:0]   _zz_1702;
  wire       [35:0]   _zz_1703;
  wire       [35:0]   _zz_1704;
  wire       [35:0]   _zz_1705;
  wire       [35:0]   _zz_1706;
  wire       [35:0]   _zz_1707;
  wire       [35:0]   _zz_1708;
  wire       [35:0]   _zz_1709;
  wire       [35:0]   _zz_1710;
  wire       [35:0]   _zz_1711;
  wire       [35:0]   _zz_1712;
  wire       [35:0]   _zz_1713;
  wire       [35:0]   _zz_1714;
  wire       [35:0]   _zz_1715;
  wire       [35:0]   _zz_1716;
  wire       [35:0]   _zz_1717;
  wire       [35:0]   _zz_1718;
  wire       [35:0]   _zz_1719;
  wire       [35:0]   _zz_1720;
  wire       [35:0]   _zz_1721;
  wire       [35:0]   _zz_1722;
  wire       [35:0]   _zz_1723;
  wire       [35:0]   _zz_1724;
  wire       [35:0]   _zz_1725;
  wire       [35:0]   _zz_1726;
  wire       [35:0]   _zz_1727;
  wire       [35:0]   _zz_1728;
  wire       [35:0]   _zz_1729;
  wire       [35:0]   _zz_1730;
  wire       [35:0]   _zz_1731;
  wire       [35:0]   _zz_1732;
  wire       [35:0]   _zz_1733;
  wire       [35:0]   _zz_1734;
  wire       [35:0]   _zz_1735;
  wire       [35:0]   _zz_1736;
  wire       [35:0]   _zz_1737;
  wire       [35:0]   _zz_1738;
  wire       [35:0]   _zz_1739;
  wire       [35:0]   _zz_1740;
  wire       [35:0]   _zz_1741;
  wire       [35:0]   _zz_1742;
  wire       [35:0]   _zz_1743;
  wire       [35:0]   _zz_1744;
  wire       [35:0]   _zz_1745;
  wire       [35:0]   _zz_1746;
  wire       [35:0]   _zz_1747;
  wire       [35:0]   _zz_1748;
  wire       [35:0]   _zz_1749;
  wire       [35:0]   _zz_1750;
  wire       [35:0]   _zz_1751;
  wire       [35:0]   _zz_1752;
  wire       [35:0]   _zz_1753;
  wire       [35:0]   _zz_1754;
  wire       [35:0]   _zz_1755;
  wire       [35:0]   _zz_1756;
  wire       [35:0]   _zz_1757;
  wire       [35:0]   _zz_1758;
  wire       [35:0]   _zz_1759;
  wire       [35:0]   _zz_1760;
  wire       [35:0]   _zz_1761;
  wire       [35:0]   _zz_1762;
  wire       [35:0]   _zz_1763;
  wire       [35:0]   _zz_1764;
  wire       [35:0]   _zz_1765;
  wire       [35:0]   _zz_1766;
  wire       [35:0]   _zz_1767;
  wire       [35:0]   _zz_1768;
  wire       [35:0]   _zz_1769;
  wire       [35:0]   _zz_1770;
  wire       [35:0]   _zz_1771;
  wire       [35:0]   _zz_1772;
  wire       [35:0]   _zz_1773;
  wire       [35:0]   _zz_1774;
  wire       [35:0]   _zz_1775;
  wire       [35:0]   _zz_1776;
  wire       [35:0]   _zz_1777;
  wire       [35:0]   _zz_1778;
  wire       [35:0]   _zz_1779;
  wire       [35:0]   _zz_1780;
  wire       [35:0]   _zz_1781;
  wire       [35:0]   _zz_1782;
  wire       [35:0]   _zz_1783;
  wire       [35:0]   _zz_1784;
  wire       [35:0]   _zz_1785;
  wire       [35:0]   _zz_1786;
  wire       [35:0]   _zz_1787;
  wire       [35:0]   _zz_1788;
  wire       [35:0]   _zz_1789;
  wire       [35:0]   _zz_1790;
  wire       [35:0]   _zz_1791;
  wire       [35:0]   _zz_1792;
  wire       [35:0]   _zz_1793;
  wire       [35:0]   _zz_1794;
  wire       [35:0]   _zz_1795;
  wire       [35:0]   _zz_1796;
  wire       [35:0]   _zz_1797;
  wire       [35:0]   _zz_1798;
  wire       [35:0]   _zz_1799;
  wire       [35:0]   _zz_1800;
  wire       [35:0]   _zz_1801;
  wire       [35:0]   _zz_1802;
  wire       [35:0]   _zz_1803;
  wire       [35:0]   _zz_1804;
  wire       [35:0]   _zz_1805;
  wire       [35:0]   _zz_1806;
  wire       [35:0]   _zz_1807;
  wire       [35:0]   _zz_1808;
  wire       [35:0]   _zz_1809;
  wire       [35:0]   _zz_1810;
  wire       [35:0]   _zz_1811;
  wire       [35:0]   _zz_1812;
  wire       [35:0]   _zz_1813;
  wire       [35:0]   _zz_1814;
  wire       [35:0]   _zz_1815;
  wire       [35:0]   _zz_1816;
  wire       [35:0]   _zz_1817;
  wire       [35:0]   _zz_1818;
  wire       [35:0]   _zz_1819;
  wire       [35:0]   _zz_1820;
  wire       [35:0]   _zz_1821;
  wire       [35:0]   _zz_1822;
  wire       [35:0]   _zz_1823;
  wire       [35:0]   _zz_1824;
  wire       [35:0]   _zz_1825;
  wire       [35:0]   _zz_1826;
  wire       [35:0]   _zz_1827;
  wire       [35:0]   _zz_1828;
  wire       [35:0]   _zz_1829;
  wire       [35:0]   _zz_1830;
  wire       [35:0]   _zz_1831;
  wire       [35:0]   _zz_1832;
  wire       [35:0]   _zz_1833;
  wire       [35:0]   _zz_1834;
  wire       [35:0]   _zz_1835;
  wire       [35:0]   _zz_1836;
  wire       [35:0]   _zz_1837;
  wire       [35:0]   _zz_1838;
  wire       [35:0]   _zz_1839;
  wire       [35:0]   _zz_1840;
  wire       [35:0]   _zz_1841;
  wire       [35:0]   _zz_1842;
  wire       [35:0]   _zz_1843;
  wire       [35:0]   _zz_1844;
  wire       [35:0]   _zz_1845;
  wire       [35:0]   _zz_1846;
  wire       [35:0]   _zz_1847;
  wire       [35:0]   _zz_1848;
  wire       [35:0]   _zz_1849;
  wire       [35:0]   _zz_1850;
  wire       [35:0]   _zz_1851;
  wire       [35:0]   _zz_1852;
  wire       [35:0]   _zz_1853;
  wire       [35:0]   _zz_1854;
  wire       [35:0]   _zz_1855;
  wire       [35:0]   _zz_1856;
  wire       [35:0]   _zz_1857;
  wire       [35:0]   _zz_1858;
  wire       [35:0]   _zz_1859;
  wire       [35:0]   _zz_1860;
  wire       [35:0]   _zz_1861;
  wire       [35:0]   _zz_1862;
  wire       [35:0]   _zz_1863;
  wire       [35:0]   _zz_1864;
  wire       [35:0]   _zz_1865;
  wire       [35:0]   _zz_1866;
  wire       [35:0]   _zz_1867;
  wire       [35:0]   _zz_1868;
  wire       [35:0]   _zz_1869;
  wire       [35:0]   _zz_1870;
  wire       [35:0]   _zz_1871;
  wire       [35:0]   _zz_1872;
  wire       [35:0]   _zz_1873;
  wire       [35:0]   _zz_1874;
  wire       [35:0]   _zz_1875;
  wire       [35:0]   _zz_1876;
  wire       [35:0]   _zz_1877;
  wire       [35:0]   _zz_1878;
  wire       [35:0]   _zz_1879;
  wire       [35:0]   _zz_1880;
  wire       [35:0]   _zz_1881;
  wire       [35:0]   _zz_1882;
  wire       [35:0]   _zz_1883;
  wire       [35:0]   _zz_1884;
  wire       [35:0]   _zz_1885;
  wire       [35:0]   _zz_1886;
  wire       [35:0]   _zz_1887;
  wire       [35:0]   _zz_1888;
  wire       [35:0]   _zz_1889;
  wire       [35:0]   _zz_1890;
  wire       [35:0]   _zz_1891;
  wire       [35:0]   _zz_1892;
  wire       [35:0]   _zz_1893;
  wire       [35:0]   _zz_1894;
  wire       [35:0]   _zz_1895;
  wire       [35:0]   _zz_1896;
  wire       [35:0]   _zz_1897;
  wire       [35:0]   _zz_1898;
  wire       [35:0]   _zz_1899;
  wire       [35:0]   _zz_1900;
  wire       [35:0]   _zz_1901;
  wire       [35:0]   _zz_1902;
  wire       [35:0]   _zz_1903;
  wire       [35:0]   _zz_1904;
  wire       [35:0]   _zz_1905;
  wire       [35:0]   _zz_1906;
  wire       [35:0]   _zz_1907;
  wire       [35:0]   _zz_1908;
  wire       [35:0]   _zz_1909;
  wire       [35:0]   _zz_1910;
  wire       [35:0]   _zz_1911;
  wire       [35:0]   _zz_1912;
  wire       [35:0]   _zz_1913;
  wire       [35:0]   _zz_1914;
  wire       [35:0]   _zz_1915;
  wire       [35:0]   _zz_1916;
  wire       [35:0]   _zz_1917;
  wire       [35:0]   _zz_1918;
  wire       [35:0]   _zz_1919;
  wire       [35:0]   _zz_1920;
  wire       [35:0]   _zz_1921;
  wire       [35:0]   _zz_1922;
  wire       [35:0]   _zz_1923;
  wire       [35:0]   _zz_1924;
  wire       [35:0]   _zz_1925;
  wire       [35:0]   _zz_1926;
  wire       [35:0]   _zz_1927;
  wire       [35:0]   _zz_1928;
  wire       [35:0]   _zz_1929;
  wire       [35:0]   _zz_1930;
  wire       [35:0]   _zz_1931;
  wire       [35:0]   _zz_1932;
  wire       [35:0]   _zz_1933;
  wire       [35:0]   _zz_1934;
  wire       [35:0]   _zz_1935;
  wire       [35:0]   _zz_1936;
  wire       [35:0]   _zz_1937;
  wire       [35:0]   _zz_1938;
  wire       [35:0]   _zz_1939;
  wire       [35:0]   _zz_1940;
  wire       [35:0]   _zz_1941;
  wire       [35:0]   _zz_1942;
  wire       [35:0]   _zz_1943;
  wire       [35:0]   _zz_1944;
  wire       [35:0]   _zz_1945;
  wire       [35:0]   _zz_1946;
  wire       [35:0]   _zz_1947;
  wire       [35:0]   _zz_1948;
  wire       [35:0]   _zz_1949;
  wire       [35:0]   _zz_1950;
  wire       [35:0]   _zz_1951;
  wire       [35:0]   _zz_1952;
  wire       [35:0]   _zz_1953;
  wire       [35:0]   _zz_1954;
  wire       [35:0]   _zz_1955;
  wire       [35:0]   _zz_1956;
  wire       [35:0]   _zz_1957;
  wire       [35:0]   _zz_1958;
  wire       [35:0]   _zz_1959;
  wire       [35:0]   _zz_1960;
  wire       [35:0]   _zz_1961;
  wire       [35:0]   _zz_1962;
  wire       [35:0]   _zz_1963;
  wire       [35:0]   _zz_1964;
  wire       [35:0]   _zz_1965;
  wire       [35:0]   _zz_1966;
  wire       [35:0]   _zz_1967;
  wire       [35:0]   _zz_1968;
  wire       [35:0]   _zz_1969;
  wire       [35:0]   _zz_1970;
  wire       [35:0]   _zz_1971;
  wire       [35:0]   _zz_1972;
  wire       [35:0]   _zz_1973;
  wire       [35:0]   _zz_1974;
  wire       [35:0]   _zz_1975;
  wire       [35:0]   _zz_1976;
  wire       [35:0]   _zz_1977;
  wire       [35:0]   _zz_1978;
  wire       [35:0]   _zz_1979;
  wire       [35:0]   _zz_1980;
  wire       [35:0]   _zz_1981;
  wire       [35:0]   _zz_1982;
  wire       [35:0]   _zz_1983;
  wire       [35:0]   _zz_1984;
  wire       [35:0]   _zz_1985;
  wire       [35:0]   _zz_1986;
  wire       [35:0]   _zz_1987;
  wire       [35:0]   _zz_1988;
  wire       [35:0]   _zz_1989;
  wire       [35:0]   _zz_1990;
  wire       [35:0]   _zz_1991;
  wire       [35:0]   _zz_1992;
  wire       [35:0]   _zz_1993;
  wire       [35:0]   _zz_1994;
  wire       [35:0]   _zz_1995;
  wire       [35:0]   _zz_1996;
  wire       [35:0]   _zz_1997;
  wire       [35:0]   _zz_1998;
  wire       [35:0]   _zz_1999;
  wire       [35:0]   _zz_2000;
  wire       [35:0]   _zz_2001;
  wire       [35:0]   _zz_2002;
  wire       [35:0]   _zz_2003;
  wire       [35:0]   _zz_2004;
  wire       [35:0]   _zz_2005;
  wire       [35:0]   _zz_2006;
  wire       [35:0]   _zz_2007;
  wire       [35:0]   _zz_2008;
  wire       [35:0]   _zz_2009;
  wire       [35:0]   _zz_2010;
  wire       [35:0]   _zz_2011;
  wire       [35:0]   _zz_2012;
  wire       [35:0]   _zz_2013;
  wire       [35:0]   _zz_2014;
  wire       [35:0]   _zz_2015;
  wire       [35:0]   _zz_2016;
  wire       [35:0]   _zz_2017;
  wire       [35:0]   _zz_2018;
  wire       [35:0]   _zz_2019;
  wire       [35:0]   _zz_2020;
  wire       [35:0]   _zz_2021;
  wire       [35:0]   _zz_2022;
  wire       [35:0]   _zz_2023;
  wire       [35:0]   _zz_2024;
  wire       [35:0]   _zz_2025;
  wire       [35:0]   _zz_2026;
  wire       [35:0]   _zz_2027;
  wire       [35:0]   _zz_2028;
  wire       [35:0]   _zz_2029;
  wire       [35:0]   _zz_2030;
  wire       [35:0]   _zz_2031;
  wire       [35:0]   _zz_2032;
  wire       [35:0]   _zz_2033;
  wire       [35:0]   _zz_2034;
  wire       [35:0]   _zz_2035;
  wire       [35:0]   _zz_2036;
  wire       [35:0]   _zz_2037;
  wire       [35:0]   _zz_2038;
  wire       [35:0]   _zz_2039;
  wire       [35:0]   _zz_2040;
  wire       [35:0]   _zz_2041;
  wire       [35:0]   _zz_2042;
  wire       [35:0]   _zz_2043;
  wire       [35:0]   _zz_2044;
  wire       [35:0]   _zz_2045;
  wire       [35:0]   _zz_2046;
  wire       [35:0]   _zz_2047;
  wire       [35:0]   _zz_2048;
  wire       [35:0]   _zz_2049;
  wire       [35:0]   _zz_2050;
  wire       [35:0]   _zz_2051;
  wire       [35:0]   _zz_2052;
  wire       [35:0]   _zz_2053;
  wire       [35:0]   _zz_2054;
  wire       [35:0]   _zz_2055;
  wire       [35:0]   _zz_2056;
  wire       [35:0]   _zz_2057;
  wire       [35:0]   _zz_2058;
  wire       [35:0]   _zz_2059;
  wire       [35:0]   _zz_2060;
  wire       [35:0]   _zz_2061;
  wire       [35:0]   _zz_2062;
  wire       [35:0]   _zz_2063;
  wire       [35:0]   _zz_2064;
  wire       [35:0]   _zz_2065;
  wire       [35:0]   _zz_2066;
  wire       [35:0]   _zz_2067;
  wire       [35:0]   _zz_2068;
  wire       [35:0]   _zz_2069;
  wire       [35:0]   _zz_2070;
  wire       [35:0]   _zz_2071;
  wire       [35:0]   _zz_2072;
  wire       [35:0]   _zz_2073;
  wire       [35:0]   _zz_2074;
  wire       [35:0]   _zz_2075;
  wire       [35:0]   _zz_2076;
  wire       [35:0]   _zz_2077;
  wire       [35:0]   _zz_2078;
  wire       [35:0]   _zz_2079;
  wire       [35:0]   _zz_2080;
  wire       [35:0]   _zz_2081;
  wire       [35:0]   _zz_2082;
  wire       [35:0]   _zz_2083;
  wire       [35:0]   _zz_2084;
  wire       [35:0]   _zz_2085;
  wire       [35:0]   _zz_2086;
  wire       [35:0]   _zz_2087;
  wire       [35:0]   _zz_2088;
  wire       [35:0]   _zz_2089;
  wire       [35:0]   _zz_2090;
  wire       [35:0]   _zz_2091;
  wire       [35:0]   _zz_2092;
  wire       [35:0]   _zz_2093;
  wire       [35:0]   _zz_2094;
  wire       [35:0]   _zz_2095;
  wire       [35:0]   _zz_2096;
  wire       [35:0]   _zz_2097;
  wire       [35:0]   _zz_2098;
  wire       [35:0]   _zz_2099;
  wire       [35:0]   _zz_2100;
  wire       [35:0]   _zz_2101;
  wire       [35:0]   _zz_2102;
  wire       [35:0]   _zz_2103;
  wire       [35:0]   _zz_2104;
  wire       [35:0]   _zz_2105;
  wire       [35:0]   _zz_2106;
  wire       [35:0]   _zz_2107;
  wire       [35:0]   _zz_2108;
  wire       [35:0]   _zz_2109;
  wire       [35:0]   _zz_2110;
  wire       [35:0]   _zz_2111;
  wire       [35:0]   _zz_2112;
  wire       [35:0]   fixTo_dout;
  wire       [35:0]   fixTo_1_dout;
  wire       [17:0]   fixTo_2_dout;
  wire       [17:0]   fixTo_3_dout;
  wire       [17:0]   fixTo_4_dout;
  wire       [17:0]   fixTo_5_dout;
  wire       [35:0]   fixTo_6_dout;
  wire       [35:0]   fixTo_7_dout;
  wire       [17:0]   fixTo_8_dout;
  wire       [17:0]   fixTo_9_dout;
  wire       [17:0]   fixTo_10_dout;
  wire       [17:0]   fixTo_11_dout;
  wire       [35:0]   fixTo_12_dout;
  wire       [35:0]   fixTo_13_dout;
  wire       [17:0]   fixTo_14_dout;
  wire       [17:0]   fixTo_15_dout;
  wire       [17:0]   fixTo_16_dout;
  wire       [17:0]   fixTo_17_dout;
  wire       [35:0]   fixTo_18_dout;
  wire       [35:0]   fixTo_19_dout;
  wire       [17:0]   fixTo_20_dout;
  wire       [17:0]   fixTo_21_dout;
  wire       [17:0]   fixTo_22_dout;
  wire       [17:0]   fixTo_23_dout;
  wire       [35:0]   fixTo_24_dout;
  wire       [35:0]   fixTo_25_dout;
  wire       [17:0]   fixTo_26_dout;
  wire       [17:0]   fixTo_27_dout;
  wire       [17:0]   fixTo_28_dout;
  wire       [17:0]   fixTo_29_dout;
  wire       [35:0]   fixTo_30_dout;
  wire       [35:0]   fixTo_31_dout;
  wire       [17:0]   fixTo_32_dout;
  wire       [17:0]   fixTo_33_dout;
  wire       [17:0]   fixTo_34_dout;
  wire       [17:0]   fixTo_35_dout;
  wire       [35:0]   fixTo_36_dout;
  wire       [35:0]   fixTo_37_dout;
  wire       [17:0]   fixTo_38_dout;
  wire       [17:0]   fixTo_39_dout;
  wire       [17:0]   fixTo_40_dout;
  wire       [17:0]   fixTo_41_dout;
  wire       [35:0]   fixTo_42_dout;
  wire       [35:0]   fixTo_43_dout;
  wire       [17:0]   fixTo_44_dout;
  wire       [17:0]   fixTo_45_dout;
  wire       [17:0]   fixTo_46_dout;
  wire       [17:0]   fixTo_47_dout;
  wire       [35:0]   fixTo_48_dout;
  wire       [35:0]   fixTo_49_dout;
  wire       [17:0]   fixTo_50_dout;
  wire       [17:0]   fixTo_51_dout;
  wire       [17:0]   fixTo_52_dout;
  wire       [17:0]   fixTo_53_dout;
  wire       [35:0]   fixTo_54_dout;
  wire       [35:0]   fixTo_55_dout;
  wire       [17:0]   fixTo_56_dout;
  wire       [17:0]   fixTo_57_dout;
  wire       [17:0]   fixTo_58_dout;
  wire       [17:0]   fixTo_59_dout;
  wire       [35:0]   fixTo_60_dout;
  wire       [35:0]   fixTo_61_dout;
  wire       [17:0]   fixTo_62_dout;
  wire       [17:0]   fixTo_63_dout;
  wire       [17:0]   fixTo_64_dout;
  wire       [17:0]   fixTo_65_dout;
  wire       [35:0]   fixTo_66_dout;
  wire       [35:0]   fixTo_67_dout;
  wire       [17:0]   fixTo_68_dout;
  wire       [17:0]   fixTo_69_dout;
  wire       [17:0]   fixTo_70_dout;
  wire       [17:0]   fixTo_71_dout;
  wire       [35:0]   fixTo_72_dout;
  wire       [35:0]   fixTo_73_dout;
  wire       [17:0]   fixTo_74_dout;
  wire       [17:0]   fixTo_75_dout;
  wire       [17:0]   fixTo_76_dout;
  wire       [17:0]   fixTo_77_dout;
  wire       [35:0]   fixTo_78_dout;
  wire       [35:0]   fixTo_79_dout;
  wire       [17:0]   fixTo_80_dout;
  wire       [17:0]   fixTo_81_dout;
  wire       [17:0]   fixTo_82_dout;
  wire       [17:0]   fixTo_83_dout;
  wire       [35:0]   fixTo_84_dout;
  wire       [35:0]   fixTo_85_dout;
  wire       [17:0]   fixTo_86_dout;
  wire       [17:0]   fixTo_87_dout;
  wire       [17:0]   fixTo_88_dout;
  wire       [17:0]   fixTo_89_dout;
  wire       [35:0]   fixTo_90_dout;
  wire       [35:0]   fixTo_91_dout;
  wire       [17:0]   fixTo_92_dout;
  wire       [17:0]   fixTo_93_dout;
  wire       [17:0]   fixTo_94_dout;
  wire       [17:0]   fixTo_95_dout;
  wire       [35:0]   fixTo_96_dout;
  wire       [35:0]   fixTo_97_dout;
  wire       [17:0]   fixTo_98_dout;
  wire       [17:0]   fixTo_99_dout;
  wire       [17:0]   fixTo_100_dout;
  wire       [17:0]   fixTo_101_dout;
  wire       [35:0]   fixTo_102_dout;
  wire       [35:0]   fixTo_103_dout;
  wire       [17:0]   fixTo_104_dout;
  wire       [17:0]   fixTo_105_dout;
  wire       [17:0]   fixTo_106_dout;
  wire       [17:0]   fixTo_107_dout;
  wire       [35:0]   fixTo_108_dout;
  wire       [35:0]   fixTo_109_dout;
  wire       [17:0]   fixTo_110_dout;
  wire       [17:0]   fixTo_111_dout;
  wire       [17:0]   fixTo_112_dout;
  wire       [17:0]   fixTo_113_dout;
  wire       [35:0]   fixTo_114_dout;
  wire       [35:0]   fixTo_115_dout;
  wire       [17:0]   fixTo_116_dout;
  wire       [17:0]   fixTo_117_dout;
  wire       [17:0]   fixTo_118_dout;
  wire       [17:0]   fixTo_119_dout;
  wire       [35:0]   fixTo_120_dout;
  wire       [35:0]   fixTo_121_dout;
  wire       [17:0]   fixTo_122_dout;
  wire       [17:0]   fixTo_123_dout;
  wire       [17:0]   fixTo_124_dout;
  wire       [17:0]   fixTo_125_dout;
  wire       [35:0]   fixTo_126_dout;
  wire       [35:0]   fixTo_127_dout;
  wire       [17:0]   fixTo_128_dout;
  wire       [17:0]   fixTo_129_dout;
  wire       [17:0]   fixTo_130_dout;
  wire       [17:0]   fixTo_131_dout;
  wire       [35:0]   fixTo_132_dout;
  wire       [35:0]   fixTo_133_dout;
  wire       [17:0]   fixTo_134_dout;
  wire       [17:0]   fixTo_135_dout;
  wire       [17:0]   fixTo_136_dout;
  wire       [17:0]   fixTo_137_dout;
  wire       [35:0]   fixTo_138_dout;
  wire       [35:0]   fixTo_139_dout;
  wire       [17:0]   fixTo_140_dout;
  wire       [17:0]   fixTo_141_dout;
  wire       [17:0]   fixTo_142_dout;
  wire       [17:0]   fixTo_143_dout;
  wire       [35:0]   fixTo_144_dout;
  wire       [35:0]   fixTo_145_dout;
  wire       [17:0]   fixTo_146_dout;
  wire       [17:0]   fixTo_147_dout;
  wire       [17:0]   fixTo_148_dout;
  wire       [17:0]   fixTo_149_dout;
  wire       [35:0]   fixTo_150_dout;
  wire       [35:0]   fixTo_151_dout;
  wire       [17:0]   fixTo_152_dout;
  wire       [17:0]   fixTo_153_dout;
  wire       [17:0]   fixTo_154_dout;
  wire       [17:0]   fixTo_155_dout;
  wire       [35:0]   fixTo_156_dout;
  wire       [35:0]   fixTo_157_dout;
  wire       [17:0]   fixTo_158_dout;
  wire       [17:0]   fixTo_159_dout;
  wire       [17:0]   fixTo_160_dout;
  wire       [17:0]   fixTo_161_dout;
  wire       [35:0]   fixTo_162_dout;
  wire       [35:0]   fixTo_163_dout;
  wire       [17:0]   fixTo_164_dout;
  wire       [17:0]   fixTo_165_dout;
  wire       [17:0]   fixTo_166_dout;
  wire       [17:0]   fixTo_167_dout;
  wire       [35:0]   fixTo_168_dout;
  wire       [35:0]   fixTo_169_dout;
  wire       [17:0]   fixTo_170_dout;
  wire       [17:0]   fixTo_171_dout;
  wire       [17:0]   fixTo_172_dout;
  wire       [17:0]   fixTo_173_dout;
  wire       [35:0]   fixTo_174_dout;
  wire       [35:0]   fixTo_175_dout;
  wire       [17:0]   fixTo_176_dout;
  wire       [17:0]   fixTo_177_dout;
  wire       [17:0]   fixTo_178_dout;
  wire       [17:0]   fixTo_179_dout;
  wire       [35:0]   fixTo_180_dout;
  wire       [35:0]   fixTo_181_dout;
  wire       [17:0]   fixTo_182_dout;
  wire       [17:0]   fixTo_183_dout;
  wire       [17:0]   fixTo_184_dout;
  wire       [17:0]   fixTo_185_dout;
  wire       [35:0]   fixTo_186_dout;
  wire       [35:0]   fixTo_187_dout;
  wire       [17:0]   fixTo_188_dout;
  wire       [17:0]   fixTo_189_dout;
  wire       [17:0]   fixTo_190_dout;
  wire       [17:0]   fixTo_191_dout;
  wire       [35:0]   fixTo_192_dout;
  wire       [35:0]   fixTo_193_dout;
  wire       [17:0]   fixTo_194_dout;
  wire       [17:0]   fixTo_195_dout;
  wire       [17:0]   fixTo_196_dout;
  wire       [17:0]   fixTo_197_dout;
  wire       [35:0]   fixTo_198_dout;
  wire       [35:0]   fixTo_199_dout;
  wire       [17:0]   fixTo_200_dout;
  wire       [17:0]   fixTo_201_dout;
  wire       [17:0]   fixTo_202_dout;
  wire       [17:0]   fixTo_203_dout;
  wire       [35:0]   fixTo_204_dout;
  wire       [35:0]   fixTo_205_dout;
  wire       [17:0]   fixTo_206_dout;
  wire       [17:0]   fixTo_207_dout;
  wire       [17:0]   fixTo_208_dout;
  wire       [17:0]   fixTo_209_dout;
  wire       [35:0]   fixTo_210_dout;
  wire       [35:0]   fixTo_211_dout;
  wire       [17:0]   fixTo_212_dout;
  wire       [17:0]   fixTo_213_dout;
  wire       [17:0]   fixTo_214_dout;
  wire       [17:0]   fixTo_215_dout;
  wire       [35:0]   fixTo_216_dout;
  wire       [35:0]   fixTo_217_dout;
  wire       [17:0]   fixTo_218_dout;
  wire       [17:0]   fixTo_219_dout;
  wire       [17:0]   fixTo_220_dout;
  wire       [17:0]   fixTo_221_dout;
  wire       [35:0]   fixTo_222_dout;
  wire       [35:0]   fixTo_223_dout;
  wire       [17:0]   fixTo_224_dout;
  wire       [17:0]   fixTo_225_dout;
  wire       [17:0]   fixTo_226_dout;
  wire       [17:0]   fixTo_227_dout;
  wire       [35:0]   fixTo_228_dout;
  wire       [35:0]   fixTo_229_dout;
  wire       [17:0]   fixTo_230_dout;
  wire       [17:0]   fixTo_231_dout;
  wire       [17:0]   fixTo_232_dout;
  wire       [17:0]   fixTo_233_dout;
  wire       [35:0]   fixTo_234_dout;
  wire       [35:0]   fixTo_235_dout;
  wire       [17:0]   fixTo_236_dout;
  wire       [17:0]   fixTo_237_dout;
  wire       [17:0]   fixTo_238_dout;
  wire       [17:0]   fixTo_239_dout;
  wire       [35:0]   fixTo_240_dout;
  wire       [35:0]   fixTo_241_dout;
  wire       [17:0]   fixTo_242_dout;
  wire       [17:0]   fixTo_243_dout;
  wire       [17:0]   fixTo_244_dout;
  wire       [17:0]   fixTo_245_dout;
  wire       [35:0]   fixTo_246_dout;
  wire       [35:0]   fixTo_247_dout;
  wire       [17:0]   fixTo_248_dout;
  wire       [17:0]   fixTo_249_dout;
  wire       [17:0]   fixTo_250_dout;
  wire       [17:0]   fixTo_251_dout;
  wire       [35:0]   fixTo_252_dout;
  wire       [35:0]   fixTo_253_dout;
  wire       [17:0]   fixTo_254_dout;
  wire       [17:0]   fixTo_255_dout;
  wire       [17:0]   fixTo_256_dout;
  wire       [17:0]   fixTo_257_dout;
  wire       [35:0]   fixTo_258_dout;
  wire       [35:0]   fixTo_259_dout;
  wire       [17:0]   fixTo_260_dout;
  wire       [17:0]   fixTo_261_dout;
  wire       [17:0]   fixTo_262_dout;
  wire       [17:0]   fixTo_263_dout;
  wire       [35:0]   fixTo_264_dout;
  wire       [35:0]   fixTo_265_dout;
  wire       [17:0]   fixTo_266_dout;
  wire       [17:0]   fixTo_267_dout;
  wire       [17:0]   fixTo_268_dout;
  wire       [17:0]   fixTo_269_dout;
  wire       [35:0]   fixTo_270_dout;
  wire       [35:0]   fixTo_271_dout;
  wire       [17:0]   fixTo_272_dout;
  wire       [17:0]   fixTo_273_dout;
  wire       [17:0]   fixTo_274_dout;
  wire       [17:0]   fixTo_275_dout;
  wire       [35:0]   fixTo_276_dout;
  wire       [35:0]   fixTo_277_dout;
  wire       [17:0]   fixTo_278_dout;
  wire       [17:0]   fixTo_279_dout;
  wire       [17:0]   fixTo_280_dout;
  wire       [17:0]   fixTo_281_dout;
  wire       [35:0]   fixTo_282_dout;
  wire       [35:0]   fixTo_283_dout;
  wire       [17:0]   fixTo_284_dout;
  wire       [17:0]   fixTo_285_dout;
  wire       [17:0]   fixTo_286_dout;
  wire       [17:0]   fixTo_287_dout;
  wire       [35:0]   fixTo_288_dout;
  wire       [35:0]   fixTo_289_dout;
  wire       [17:0]   fixTo_290_dout;
  wire       [17:0]   fixTo_291_dout;
  wire       [17:0]   fixTo_292_dout;
  wire       [17:0]   fixTo_293_dout;
  wire       [35:0]   fixTo_294_dout;
  wire       [35:0]   fixTo_295_dout;
  wire       [17:0]   fixTo_296_dout;
  wire       [17:0]   fixTo_297_dout;
  wire       [17:0]   fixTo_298_dout;
  wire       [17:0]   fixTo_299_dout;
  wire       [35:0]   fixTo_300_dout;
  wire       [35:0]   fixTo_301_dout;
  wire       [17:0]   fixTo_302_dout;
  wire       [17:0]   fixTo_303_dout;
  wire       [17:0]   fixTo_304_dout;
  wire       [17:0]   fixTo_305_dout;
  wire       [35:0]   fixTo_306_dout;
  wire       [35:0]   fixTo_307_dout;
  wire       [17:0]   fixTo_308_dout;
  wire       [17:0]   fixTo_309_dout;
  wire       [17:0]   fixTo_310_dout;
  wire       [17:0]   fixTo_311_dout;
  wire       [35:0]   fixTo_312_dout;
  wire       [35:0]   fixTo_313_dout;
  wire       [17:0]   fixTo_314_dout;
  wire       [17:0]   fixTo_315_dout;
  wire       [17:0]   fixTo_316_dout;
  wire       [17:0]   fixTo_317_dout;
  wire       [35:0]   fixTo_318_dout;
  wire       [35:0]   fixTo_319_dout;
  wire       [17:0]   fixTo_320_dout;
  wire       [17:0]   fixTo_321_dout;
  wire       [17:0]   fixTo_322_dout;
  wire       [17:0]   fixTo_323_dout;
  wire       [35:0]   fixTo_324_dout;
  wire       [35:0]   fixTo_325_dout;
  wire       [17:0]   fixTo_326_dout;
  wire       [17:0]   fixTo_327_dout;
  wire       [17:0]   fixTo_328_dout;
  wire       [17:0]   fixTo_329_dout;
  wire       [35:0]   fixTo_330_dout;
  wire       [35:0]   fixTo_331_dout;
  wire       [17:0]   fixTo_332_dout;
  wire       [17:0]   fixTo_333_dout;
  wire       [17:0]   fixTo_334_dout;
  wire       [17:0]   fixTo_335_dout;
  wire       [35:0]   fixTo_336_dout;
  wire       [35:0]   fixTo_337_dout;
  wire       [17:0]   fixTo_338_dout;
  wire       [17:0]   fixTo_339_dout;
  wire       [17:0]   fixTo_340_dout;
  wire       [17:0]   fixTo_341_dout;
  wire       [35:0]   fixTo_342_dout;
  wire       [35:0]   fixTo_343_dout;
  wire       [17:0]   fixTo_344_dout;
  wire       [17:0]   fixTo_345_dout;
  wire       [17:0]   fixTo_346_dout;
  wire       [17:0]   fixTo_347_dout;
  wire       [35:0]   fixTo_348_dout;
  wire       [35:0]   fixTo_349_dout;
  wire       [17:0]   fixTo_350_dout;
  wire       [17:0]   fixTo_351_dout;
  wire       [17:0]   fixTo_352_dout;
  wire       [17:0]   fixTo_353_dout;
  wire       [35:0]   fixTo_354_dout;
  wire       [35:0]   fixTo_355_dout;
  wire       [17:0]   fixTo_356_dout;
  wire       [17:0]   fixTo_357_dout;
  wire       [17:0]   fixTo_358_dout;
  wire       [17:0]   fixTo_359_dout;
  wire       [35:0]   fixTo_360_dout;
  wire       [35:0]   fixTo_361_dout;
  wire       [17:0]   fixTo_362_dout;
  wire       [17:0]   fixTo_363_dout;
  wire       [17:0]   fixTo_364_dout;
  wire       [17:0]   fixTo_365_dout;
  wire       [35:0]   fixTo_366_dout;
  wire       [35:0]   fixTo_367_dout;
  wire       [17:0]   fixTo_368_dout;
  wire       [17:0]   fixTo_369_dout;
  wire       [17:0]   fixTo_370_dout;
  wire       [17:0]   fixTo_371_dout;
  wire       [35:0]   fixTo_372_dout;
  wire       [35:0]   fixTo_373_dout;
  wire       [17:0]   fixTo_374_dout;
  wire       [17:0]   fixTo_375_dout;
  wire       [17:0]   fixTo_376_dout;
  wire       [17:0]   fixTo_377_dout;
  wire       [35:0]   fixTo_378_dout;
  wire       [35:0]   fixTo_379_dout;
  wire       [17:0]   fixTo_380_dout;
  wire       [17:0]   fixTo_381_dout;
  wire       [17:0]   fixTo_382_dout;
  wire       [17:0]   fixTo_383_dout;
  wire       [35:0]   fixTo_384_dout;
  wire       [35:0]   fixTo_385_dout;
  wire       [17:0]   fixTo_386_dout;
  wire       [17:0]   fixTo_387_dout;
  wire       [17:0]   fixTo_388_dout;
  wire       [17:0]   fixTo_389_dout;
  wire       [35:0]   fixTo_390_dout;
  wire       [35:0]   fixTo_391_dout;
  wire       [17:0]   fixTo_392_dout;
  wire       [17:0]   fixTo_393_dout;
  wire       [17:0]   fixTo_394_dout;
  wire       [17:0]   fixTo_395_dout;
  wire       [35:0]   fixTo_396_dout;
  wire       [35:0]   fixTo_397_dout;
  wire       [17:0]   fixTo_398_dout;
  wire       [17:0]   fixTo_399_dout;
  wire       [17:0]   fixTo_400_dout;
  wire       [17:0]   fixTo_401_dout;
  wire       [35:0]   fixTo_402_dout;
  wire       [35:0]   fixTo_403_dout;
  wire       [17:0]   fixTo_404_dout;
  wire       [17:0]   fixTo_405_dout;
  wire       [17:0]   fixTo_406_dout;
  wire       [17:0]   fixTo_407_dout;
  wire       [35:0]   fixTo_408_dout;
  wire       [35:0]   fixTo_409_dout;
  wire       [17:0]   fixTo_410_dout;
  wire       [17:0]   fixTo_411_dout;
  wire       [17:0]   fixTo_412_dout;
  wire       [17:0]   fixTo_413_dout;
  wire       [35:0]   fixTo_414_dout;
  wire       [35:0]   fixTo_415_dout;
  wire       [17:0]   fixTo_416_dout;
  wire       [17:0]   fixTo_417_dout;
  wire       [17:0]   fixTo_418_dout;
  wire       [17:0]   fixTo_419_dout;
  wire       [35:0]   fixTo_420_dout;
  wire       [35:0]   fixTo_421_dout;
  wire       [17:0]   fixTo_422_dout;
  wire       [17:0]   fixTo_423_dout;
  wire       [17:0]   fixTo_424_dout;
  wire       [17:0]   fixTo_425_dout;
  wire       [35:0]   fixTo_426_dout;
  wire       [35:0]   fixTo_427_dout;
  wire       [17:0]   fixTo_428_dout;
  wire       [17:0]   fixTo_429_dout;
  wire       [17:0]   fixTo_430_dout;
  wire       [17:0]   fixTo_431_dout;
  wire       [35:0]   fixTo_432_dout;
  wire       [35:0]   fixTo_433_dout;
  wire       [17:0]   fixTo_434_dout;
  wire       [17:0]   fixTo_435_dout;
  wire       [17:0]   fixTo_436_dout;
  wire       [17:0]   fixTo_437_dout;
  wire       [35:0]   fixTo_438_dout;
  wire       [35:0]   fixTo_439_dout;
  wire       [17:0]   fixTo_440_dout;
  wire       [17:0]   fixTo_441_dout;
  wire       [17:0]   fixTo_442_dout;
  wire       [17:0]   fixTo_443_dout;
  wire       [35:0]   fixTo_444_dout;
  wire       [35:0]   fixTo_445_dout;
  wire       [17:0]   fixTo_446_dout;
  wire       [17:0]   fixTo_447_dout;
  wire       [17:0]   fixTo_448_dout;
  wire       [17:0]   fixTo_449_dout;
  wire       [35:0]   fixTo_450_dout;
  wire       [35:0]   fixTo_451_dout;
  wire       [17:0]   fixTo_452_dout;
  wire       [17:0]   fixTo_453_dout;
  wire       [17:0]   fixTo_454_dout;
  wire       [17:0]   fixTo_455_dout;
  wire       [35:0]   fixTo_456_dout;
  wire       [35:0]   fixTo_457_dout;
  wire       [17:0]   fixTo_458_dout;
  wire       [17:0]   fixTo_459_dout;
  wire       [17:0]   fixTo_460_dout;
  wire       [17:0]   fixTo_461_dout;
  wire       [35:0]   fixTo_462_dout;
  wire       [35:0]   fixTo_463_dout;
  wire       [17:0]   fixTo_464_dout;
  wire       [17:0]   fixTo_465_dout;
  wire       [17:0]   fixTo_466_dout;
  wire       [17:0]   fixTo_467_dout;
  wire       [35:0]   fixTo_468_dout;
  wire       [35:0]   fixTo_469_dout;
  wire       [17:0]   fixTo_470_dout;
  wire       [17:0]   fixTo_471_dout;
  wire       [17:0]   fixTo_472_dout;
  wire       [17:0]   fixTo_473_dout;
  wire       [35:0]   fixTo_474_dout;
  wire       [35:0]   fixTo_475_dout;
  wire       [17:0]   fixTo_476_dout;
  wire       [17:0]   fixTo_477_dout;
  wire       [17:0]   fixTo_478_dout;
  wire       [17:0]   fixTo_479_dout;
  wire       [35:0]   fixTo_480_dout;
  wire       [35:0]   fixTo_481_dout;
  wire       [17:0]   fixTo_482_dout;
  wire       [17:0]   fixTo_483_dout;
  wire       [17:0]   fixTo_484_dout;
  wire       [17:0]   fixTo_485_dout;
  wire       [35:0]   fixTo_486_dout;
  wire       [35:0]   fixTo_487_dout;
  wire       [17:0]   fixTo_488_dout;
  wire       [17:0]   fixTo_489_dout;
  wire       [17:0]   fixTo_490_dout;
  wire       [17:0]   fixTo_491_dout;
  wire       [35:0]   fixTo_492_dout;
  wire       [35:0]   fixTo_493_dout;
  wire       [17:0]   fixTo_494_dout;
  wire       [17:0]   fixTo_495_dout;
  wire       [17:0]   fixTo_496_dout;
  wire       [17:0]   fixTo_497_dout;
  wire       [35:0]   fixTo_498_dout;
  wire       [35:0]   fixTo_499_dout;
  wire       [17:0]   fixTo_500_dout;
  wire       [17:0]   fixTo_501_dout;
  wire       [17:0]   fixTo_502_dout;
  wire       [17:0]   fixTo_503_dout;
  wire       [35:0]   fixTo_504_dout;
  wire       [35:0]   fixTo_505_dout;
  wire       [17:0]   fixTo_506_dout;
  wire       [17:0]   fixTo_507_dout;
  wire       [17:0]   fixTo_508_dout;
  wire       [17:0]   fixTo_509_dout;
  wire       [35:0]   fixTo_510_dout;
  wire       [35:0]   fixTo_511_dout;
  wire       [17:0]   fixTo_512_dout;
  wire       [17:0]   fixTo_513_dout;
  wire       [17:0]   fixTo_514_dout;
  wire       [17:0]   fixTo_515_dout;
  wire       [35:0]   fixTo_516_dout;
  wire       [35:0]   fixTo_517_dout;
  wire       [17:0]   fixTo_518_dout;
  wire       [17:0]   fixTo_519_dout;
  wire       [17:0]   fixTo_520_dout;
  wire       [17:0]   fixTo_521_dout;
  wire       [35:0]   fixTo_522_dout;
  wire       [35:0]   fixTo_523_dout;
  wire       [17:0]   fixTo_524_dout;
  wire       [17:0]   fixTo_525_dout;
  wire       [17:0]   fixTo_526_dout;
  wire       [17:0]   fixTo_527_dout;
  wire       [35:0]   fixTo_528_dout;
  wire       [35:0]   fixTo_529_dout;
  wire       [17:0]   fixTo_530_dout;
  wire       [17:0]   fixTo_531_dout;
  wire       [17:0]   fixTo_532_dout;
  wire       [17:0]   fixTo_533_dout;
  wire       [35:0]   fixTo_534_dout;
  wire       [35:0]   fixTo_535_dout;
  wire       [17:0]   fixTo_536_dout;
  wire       [17:0]   fixTo_537_dout;
  wire       [17:0]   fixTo_538_dout;
  wire       [17:0]   fixTo_539_dout;
  wire       [35:0]   fixTo_540_dout;
  wire       [35:0]   fixTo_541_dout;
  wire       [17:0]   fixTo_542_dout;
  wire       [17:0]   fixTo_543_dout;
  wire       [17:0]   fixTo_544_dout;
  wire       [17:0]   fixTo_545_dout;
  wire       [35:0]   fixTo_546_dout;
  wire       [35:0]   fixTo_547_dout;
  wire       [17:0]   fixTo_548_dout;
  wire       [17:0]   fixTo_549_dout;
  wire       [17:0]   fixTo_550_dout;
  wire       [17:0]   fixTo_551_dout;
  wire       [35:0]   fixTo_552_dout;
  wire       [35:0]   fixTo_553_dout;
  wire       [17:0]   fixTo_554_dout;
  wire       [17:0]   fixTo_555_dout;
  wire       [17:0]   fixTo_556_dout;
  wire       [17:0]   fixTo_557_dout;
  wire       [35:0]   fixTo_558_dout;
  wire       [35:0]   fixTo_559_dout;
  wire       [17:0]   fixTo_560_dout;
  wire       [17:0]   fixTo_561_dout;
  wire       [17:0]   fixTo_562_dout;
  wire       [17:0]   fixTo_563_dout;
  wire       [35:0]   fixTo_564_dout;
  wire       [35:0]   fixTo_565_dout;
  wire       [17:0]   fixTo_566_dout;
  wire       [17:0]   fixTo_567_dout;
  wire       [17:0]   fixTo_568_dout;
  wire       [17:0]   fixTo_569_dout;
  wire       [35:0]   fixTo_570_dout;
  wire       [35:0]   fixTo_571_dout;
  wire       [17:0]   fixTo_572_dout;
  wire       [17:0]   fixTo_573_dout;
  wire       [17:0]   fixTo_574_dout;
  wire       [17:0]   fixTo_575_dout;
  wire       [35:0]   fixTo_576_dout;
  wire       [35:0]   fixTo_577_dout;
  wire       [17:0]   fixTo_578_dout;
  wire       [17:0]   fixTo_579_dout;
  wire       [17:0]   fixTo_580_dout;
  wire       [17:0]   fixTo_581_dout;
  wire       [35:0]   fixTo_582_dout;
  wire       [35:0]   fixTo_583_dout;
  wire       [17:0]   fixTo_584_dout;
  wire       [17:0]   fixTo_585_dout;
  wire       [17:0]   fixTo_586_dout;
  wire       [17:0]   fixTo_587_dout;
  wire       [35:0]   fixTo_588_dout;
  wire       [35:0]   fixTo_589_dout;
  wire       [17:0]   fixTo_590_dout;
  wire       [17:0]   fixTo_591_dout;
  wire       [17:0]   fixTo_592_dout;
  wire       [17:0]   fixTo_593_dout;
  wire       [35:0]   fixTo_594_dout;
  wire       [35:0]   fixTo_595_dout;
  wire       [17:0]   fixTo_596_dout;
  wire       [17:0]   fixTo_597_dout;
  wire       [17:0]   fixTo_598_dout;
  wire       [17:0]   fixTo_599_dout;
  wire       [35:0]   fixTo_600_dout;
  wire       [35:0]   fixTo_601_dout;
  wire       [17:0]   fixTo_602_dout;
  wire       [17:0]   fixTo_603_dout;
  wire       [17:0]   fixTo_604_dout;
  wire       [17:0]   fixTo_605_dout;
  wire       [35:0]   fixTo_606_dout;
  wire       [35:0]   fixTo_607_dout;
  wire       [17:0]   fixTo_608_dout;
  wire       [17:0]   fixTo_609_dout;
  wire       [17:0]   fixTo_610_dout;
  wire       [17:0]   fixTo_611_dout;
  wire       [35:0]   fixTo_612_dout;
  wire       [35:0]   fixTo_613_dout;
  wire       [17:0]   fixTo_614_dout;
  wire       [17:0]   fixTo_615_dout;
  wire       [17:0]   fixTo_616_dout;
  wire       [17:0]   fixTo_617_dout;
  wire       [35:0]   fixTo_618_dout;
  wire       [35:0]   fixTo_619_dout;
  wire       [17:0]   fixTo_620_dout;
  wire       [17:0]   fixTo_621_dout;
  wire       [17:0]   fixTo_622_dout;
  wire       [17:0]   fixTo_623_dout;
  wire       [35:0]   fixTo_624_dout;
  wire       [35:0]   fixTo_625_dout;
  wire       [17:0]   fixTo_626_dout;
  wire       [17:0]   fixTo_627_dout;
  wire       [17:0]   fixTo_628_dout;
  wire       [17:0]   fixTo_629_dout;
  wire       [35:0]   fixTo_630_dout;
  wire       [35:0]   fixTo_631_dout;
  wire       [17:0]   fixTo_632_dout;
  wire       [17:0]   fixTo_633_dout;
  wire       [17:0]   fixTo_634_dout;
  wire       [17:0]   fixTo_635_dout;
  wire       [35:0]   fixTo_636_dout;
  wire       [35:0]   fixTo_637_dout;
  wire       [17:0]   fixTo_638_dout;
  wire       [17:0]   fixTo_639_dout;
  wire       [17:0]   fixTo_640_dout;
  wire       [17:0]   fixTo_641_dout;
  wire       [35:0]   fixTo_642_dout;
  wire       [35:0]   fixTo_643_dout;
  wire       [17:0]   fixTo_644_dout;
  wire       [17:0]   fixTo_645_dout;
  wire       [17:0]   fixTo_646_dout;
  wire       [17:0]   fixTo_647_dout;
  wire       [35:0]   fixTo_648_dout;
  wire       [35:0]   fixTo_649_dout;
  wire       [17:0]   fixTo_650_dout;
  wire       [17:0]   fixTo_651_dout;
  wire       [17:0]   fixTo_652_dout;
  wire       [17:0]   fixTo_653_dout;
  wire       [35:0]   fixTo_654_dout;
  wire       [35:0]   fixTo_655_dout;
  wire       [17:0]   fixTo_656_dout;
  wire       [17:0]   fixTo_657_dout;
  wire       [17:0]   fixTo_658_dout;
  wire       [17:0]   fixTo_659_dout;
  wire       [35:0]   fixTo_660_dout;
  wire       [35:0]   fixTo_661_dout;
  wire       [17:0]   fixTo_662_dout;
  wire       [17:0]   fixTo_663_dout;
  wire       [17:0]   fixTo_664_dout;
  wire       [17:0]   fixTo_665_dout;
  wire       [35:0]   fixTo_666_dout;
  wire       [35:0]   fixTo_667_dout;
  wire       [17:0]   fixTo_668_dout;
  wire       [17:0]   fixTo_669_dout;
  wire       [17:0]   fixTo_670_dout;
  wire       [17:0]   fixTo_671_dout;
  wire       [35:0]   fixTo_672_dout;
  wire       [35:0]   fixTo_673_dout;
  wire       [17:0]   fixTo_674_dout;
  wire       [17:0]   fixTo_675_dout;
  wire       [17:0]   fixTo_676_dout;
  wire       [17:0]   fixTo_677_dout;
  wire       [35:0]   fixTo_678_dout;
  wire       [35:0]   fixTo_679_dout;
  wire       [17:0]   fixTo_680_dout;
  wire       [17:0]   fixTo_681_dout;
  wire       [17:0]   fixTo_682_dout;
  wire       [17:0]   fixTo_683_dout;
  wire       [35:0]   fixTo_684_dout;
  wire       [35:0]   fixTo_685_dout;
  wire       [17:0]   fixTo_686_dout;
  wire       [17:0]   fixTo_687_dout;
  wire       [17:0]   fixTo_688_dout;
  wire       [17:0]   fixTo_689_dout;
  wire       [35:0]   fixTo_690_dout;
  wire       [35:0]   fixTo_691_dout;
  wire       [17:0]   fixTo_692_dout;
  wire       [17:0]   fixTo_693_dout;
  wire       [17:0]   fixTo_694_dout;
  wire       [17:0]   fixTo_695_dout;
  wire       [35:0]   fixTo_696_dout;
  wire       [35:0]   fixTo_697_dout;
  wire       [17:0]   fixTo_698_dout;
  wire       [17:0]   fixTo_699_dout;
  wire       [17:0]   fixTo_700_dout;
  wire       [17:0]   fixTo_701_dout;
  wire       [35:0]   fixTo_702_dout;
  wire       [35:0]   fixTo_703_dout;
  wire       [17:0]   fixTo_704_dout;
  wire       [17:0]   fixTo_705_dout;
  wire       [17:0]   fixTo_706_dout;
  wire       [17:0]   fixTo_707_dout;
  wire       [35:0]   fixTo_708_dout;
  wire       [35:0]   fixTo_709_dout;
  wire       [17:0]   fixTo_710_dout;
  wire       [17:0]   fixTo_711_dout;
  wire       [17:0]   fixTo_712_dout;
  wire       [17:0]   fixTo_713_dout;
  wire       [35:0]   fixTo_714_dout;
  wire       [35:0]   fixTo_715_dout;
  wire       [17:0]   fixTo_716_dout;
  wire       [17:0]   fixTo_717_dout;
  wire       [17:0]   fixTo_718_dout;
  wire       [17:0]   fixTo_719_dout;
  wire       [35:0]   fixTo_720_dout;
  wire       [35:0]   fixTo_721_dout;
  wire       [17:0]   fixTo_722_dout;
  wire       [17:0]   fixTo_723_dout;
  wire       [17:0]   fixTo_724_dout;
  wire       [17:0]   fixTo_725_dout;
  wire       [35:0]   fixTo_726_dout;
  wire       [35:0]   fixTo_727_dout;
  wire       [17:0]   fixTo_728_dout;
  wire       [17:0]   fixTo_729_dout;
  wire       [17:0]   fixTo_730_dout;
  wire       [17:0]   fixTo_731_dout;
  wire       [35:0]   fixTo_732_dout;
  wire       [35:0]   fixTo_733_dout;
  wire       [17:0]   fixTo_734_dout;
  wire       [17:0]   fixTo_735_dout;
  wire       [17:0]   fixTo_736_dout;
  wire       [17:0]   fixTo_737_dout;
  wire       [35:0]   fixTo_738_dout;
  wire       [35:0]   fixTo_739_dout;
  wire       [17:0]   fixTo_740_dout;
  wire       [17:0]   fixTo_741_dout;
  wire       [17:0]   fixTo_742_dout;
  wire       [17:0]   fixTo_743_dout;
  wire       [35:0]   fixTo_744_dout;
  wire       [35:0]   fixTo_745_dout;
  wire       [17:0]   fixTo_746_dout;
  wire       [17:0]   fixTo_747_dout;
  wire       [17:0]   fixTo_748_dout;
  wire       [17:0]   fixTo_749_dout;
  wire       [35:0]   fixTo_750_dout;
  wire       [35:0]   fixTo_751_dout;
  wire       [17:0]   fixTo_752_dout;
  wire       [17:0]   fixTo_753_dout;
  wire       [17:0]   fixTo_754_dout;
  wire       [17:0]   fixTo_755_dout;
  wire       [35:0]   fixTo_756_dout;
  wire       [35:0]   fixTo_757_dout;
  wire       [17:0]   fixTo_758_dout;
  wire       [17:0]   fixTo_759_dout;
  wire       [17:0]   fixTo_760_dout;
  wire       [17:0]   fixTo_761_dout;
  wire       [35:0]   fixTo_762_dout;
  wire       [35:0]   fixTo_763_dout;
  wire       [17:0]   fixTo_764_dout;
  wire       [17:0]   fixTo_765_dout;
  wire       [17:0]   fixTo_766_dout;
  wire       [17:0]   fixTo_767_dout;
  wire       [35:0]   fixTo_768_dout;
  wire       [35:0]   fixTo_769_dout;
  wire       [17:0]   fixTo_770_dout;
  wire       [17:0]   fixTo_771_dout;
  wire       [17:0]   fixTo_772_dout;
  wire       [17:0]   fixTo_773_dout;
  wire       [35:0]   fixTo_774_dout;
  wire       [35:0]   fixTo_775_dout;
  wire       [17:0]   fixTo_776_dout;
  wire       [17:0]   fixTo_777_dout;
  wire       [17:0]   fixTo_778_dout;
  wire       [17:0]   fixTo_779_dout;
  wire       [35:0]   fixTo_780_dout;
  wire       [35:0]   fixTo_781_dout;
  wire       [17:0]   fixTo_782_dout;
  wire       [17:0]   fixTo_783_dout;
  wire       [17:0]   fixTo_784_dout;
  wire       [17:0]   fixTo_785_dout;
  wire       [35:0]   fixTo_786_dout;
  wire       [35:0]   fixTo_787_dout;
  wire       [17:0]   fixTo_788_dout;
  wire       [17:0]   fixTo_789_dout;
  wire       [17:0]   fixTo_790_dout;
  wire       [17:0]   fixTo_791_dout;
  wire       [35:0]   fixTo_792_dout;
  wire       [35:0]   fixTo_793_dout;
  wire       [17:0]   fixTo_794_dout;
  wire       [17:0]   fixTo_795_dout;
  wire       [17:0]   fixTo_796_dout;
  wire       [17:0]   fixTo_797_dout;
  wire       [35:0]   fixTo_798_dout;
  wire       [35:0]   fixTo_799_dout;
  wire       [17:0]   fixTo_800_dout;
  wire       [17:0]   fixTo_801_dout;
  wire       [17:0]   fixTo_802_dout;
  wire       [17:0]   fixTo_803_dout;
  wire       [35:0]   fixTo_804_dout;
  wire       [35:0]   fixTo_805_dout;
  wire       [17:0]   fixTo_806_dout;
  wire       [17:0]   fixTo_807_dout;
  wire       [17:0]   fixTo_808_dout;
  wire       [17:0]   fixTo_809_dout;
  wire       [35:0]   fixTo_810_dout;
  wire       [35:0]   fixTo_811_dout;
  wire       [17:0]   fixTo_812_dout;
  wire       [17:0]   fixTo_813_dout;
  wire       [17:0]   fixTo_814_dout;
  wire       [17:0]   fixTo_815_dout;
  wire       [35:0]   fixTo_816_dout;
  wire       [35:0]   fixTo_817_dout;
  wire       [17:0]   fixTo_818_dout;
  wire       [17:0]   fixTo_819_dout;
  wire       [17:0]   fixTo_820_dout;
  wire       [17:0]   fixTo_821_dout;
  wire       [35:0]   fixTo_822_dout;
  wire       [35:0]   fixTo_823_dout;
  wire       [17:0]   fixTo_824_dout;
  wire       [17:0]   fixTo_825_dout;
  wire       [17:0]   fixTo_826_dout;
  wire       [17:0]   fixTo_827_dout;
  wire       [35:0]   fixTo_828_dout;
  wire       [35:0]   fixTo_829_dout;
  wire       [17:0]   fixTo_830_dout;
  wire       [17:0]   fixTo_831_dout;
  wire       [17:0]   fixTo_832_dout;
  wire       [17:0]   fixTo_833_dout;
  wire       [35:0]   fixTo_834_dout;
  wire       [35:0]   fixTo_835_dout;
  wire       [17:0]   fixTo_836_dout;
  wire       [17:0]   fixTo_837_dout;
  wire       [17:0]   fixTo_838_dout;
  wire       [17:0]   fixTo_839_dout;
  wire       [35:0]   fixTo_840_dout;
  wire       [35:0]   fixTo_841_dout;
  wire       [17:0]   fixTo_842_dout;
  wire       [17:0]   fixTo_843_dout;
  wire       [17:0]   fixTo_844_dout;
  wire       [17:0]   fixTo_845_dout;
  wire       [35:0]   fixTo_846_dout;
  wire       [35:0]   fixTo_847_dout;
  wire       [17:0]   fixTo_848_dout;
  wire       [17:0]   fixTo_849_dout;
  wire       [17:0]   fixTo_850_dout;
  wire       [17:0]   fixTo_851_dout;
  wire       [35:0]   fixTo_852_dout;
  wire       [35:0]   fixTo_853_dout;
  wire       [17:0]   fixTo_854_dout;
  wire       [17:0]   fixTo_855_dout;
  wire       [17:0]   fixTo_856_dout;
  wire       [17:0]   fixTo_857_dout;
  wire       [35:0]   fixTo_858_dout;
  wire       [35:0]   fixTo_859_dout;
  wire       [17:0]   fixTo_860_dout;
  wire       [17:0]   fixTo_861_dout;
  wire       [17:0]   fixTo_862_dout;
  wire       [17:0]   fixTo_863_dout;
  wire       [35:0]   fixTo_864_dout;
  wire       [35:0]   fixTo_865_dout;
  wire       [17:0]   fixTo_866_dout;
  wire       [17:0]   fixTo_867_dout;
  wire       [17:0]   fixTo_868_dout;
  wire       [17:0]   fixTo_869_dout;
  wire       [35:0]   fixTo_870_dout;
  wire       [35:0]   fixTo_871_dout;
  wire       [17:0]   fixTo_872_dout;
  wire       [17:0]   fixTo_873_dout;
  wire       [17:0]   fixTo_874_dout;
  wire       [17:0]   fixTo_875_dout;
  wire       [35:0]   fixTo_876_dout;
  wire       [35:0]   fixTo_877_dout;
  wire       [17:0]   fixTo_878_dout;
  wire       [17:0]   fixTo_879_dout;
  wire       [17:0]   fixTo_880_dout;
  wire       [17:0]   fixTo_881_dout;
  wire       [35:0]   fixTo_882_dout;
  wire       [35:0]   fixTo_883_dout;
  wire       [17:0]   fixTo_884_dout;
  wire       [17:0]   fixTo_885_dout;
  wire       [17:0]   fixTo_886_dout;
  wire       [17:0]   fixTo_887_dout;
  wire       [35:0]   fixTo_888_dout;
  wire       [35:0]   fixTo_889_dout;
  wire       [17:0]   fixTo_890_dout;
  wire       [17:0]   fixTo_891_dout;
  wire       [17:0]   fixTo_892_dout;
  wire       [17:0]   fixTo_893_dout;
  wire       [35:0]   fixTo_894_dout;
  wire       [35:0]   fixTo_895_dout;
  wire       [17:0]   fixTo_896_dout;
  wire       [17:0]   fixTo_897_dout;
  wire       [17:0]   fixTo_898_dout;
  wire       [17:0]   fixTo_899_dout;
  wire       [35:0]   fixTo_900_dout;
  wire       [35:0]   fixTo_901_dout;
  wire       [17:0]   fixTo_902_dout;
  wire       [17:0]   fixTo_903_dout;
  wire       [17:0]   fixTo_904_dout;
  wire       [17:0]   fixTo_905_dout;
  wire       [35:0]   fixTo_906_dout;
  wire       [35:0]   fixTo_907_dout;
  wire       [17:0]   fixTo_908_dout;
  wire       [17:0]   fixTo_909_dout;
  wire       [17:0]   fixTo_910_dout;
  wire       [17:0]   fixTo_911_dout;
  wire       [35:0]   fixTo_912_dout;
  wire       [35:0]   fixTo_913_dout;
  wire       [17:0]   fixTo_914_dout;
  wire       [17:0]   fixTo_915_dout;
  wire       [17:0]   fixTo_916_dout;
  wire       [17:0]   fixTo_917_dout;
  wire       [35:0]   fixTo_918_dout;
  wire       [35:0]   fixTo_919_dout;
  wire       [17:0]   fixTo_920_dout;
  wire       [17:0]   fixTo_921_dout;
  wire       [17:0]   fixTo_922_dout;
  wire       [17:0]   fixTo_923_dout;
  wire       [35:0]   fixTo_924_dout;
  wire       [35:0]   fixTo_925_dout;
  wire       [17:0]   fixTo_926_dout;
  wire       [17:0]   fixTo_927_dout;
  wire       [17:0]   fixTo_928_dout;
  wire       [17:0]   fixTo_929_dout;
  wire       [35:0]   fixTo_930_dout;
  wire       [35:0]   fixTo_931_dout;
  wire       [17:0]   fixTo_932_dout;
  wire       [17:0]   fixTo_933_dout;
  wire       [17:0]   fixTo_934_dout;
  wire       [17:0]   fixTo_935_dout;
  wire       [35:0]   fixTo_936_dout;
  wire       [35:0]   fixTo_937_dout;
  wire       [17:0]   fixTo_938_dout;
  wire       [17:0]   fixTo_939_dout;
  wire       [17:0]   fixTo_940_dout;
  wire       [17:0]   fixTo_941_dout;
  wire       [35:0]   fixTo_942_dout;
  wire       [35:0]   fixTo_943_dout;
  wire       [17:0]   fixTo_944_dout;
  wire       [17:0]   fixTo_945_dout;
  wire       [17:0]   fixTo_946_dout;
  wire       [17:0]   fixTo_947_dout;
  wire       [35:0]   fixTo_948_dout;
  wire       [35:0]   fixTo_949_dout;
  wire       [17:0]   fixTo_950_dout;
  wire       [17:0]   fixTo_951_dout;
  wire       [17:0]   fixTo_952_dout;
  wire       [17:0]   fixTo_953_dout;
  wire       [35:0]   fixTo_954_dout;
  wire       [35:0]   fixTo_955_dout;
  wire       [17:0]   fixTo_956_dout;
  wire       [17:0]   fixTo_957_dout;
  wire       [17:0]   fixTo_958_dout;
  wire       [17:0]   fixTo_959_dout;
  wire       [35:0]   fixTo_960_dout;
  wire       [35:0]   fixTo_961_dout;
  wire       [17:0]   fixTo_962_dout;
  wire       [17:0]   fixTo_963_dout;
  wire       [17:0]   fixTo_964_dout;
  wire       [17:0]   fixTo_965_dout;
  wire       [35:0]   fixTo_966_dout;
  wire       [35:0]   fixTo_967_dout;
  wire       [17:0]   fixTo_968_dout;
  wire       [17:0]   fixTo_969_dout;
  wire       [17:0]   fixTo_970_dout;
  wire       [17:0]   fixTo_971_dout;
  wire       [35:0]   fixTo_972_dout;
  wire       [35:0]   fixTo_973_dout;
  wire       [17:0]   fixTo_974_dout;
  wire       [17:0]   fixTo_975_dout;
  wire       [17:0]   fixTo_976_dout;
  wire       [17:0]   fixTo_977_dout;
  wire       [35:0]   fixTo_978_dout;
  wire       [35:0]   fixTo_979_dout;
  wire       [17:0]   fixTo_980_dout;
  wire       [17:0]   fixTo_981_dout;
  wire       [17:0]   fixTo_982_dout;
  wire       [17:0]   fixTo_983_dout;
  wire       [35:0]   fixTo_984_dout;
  wire       [35:0]   fixTo_985_dout;
  wire       [17:0]   fixTo_986_dout;
  wire       [17:0]   fixTo_987_dout;
  wire       [17:0]   fixTo_988_dout;
  wire       [17:0]   fixTo_989_dout;
  wire       [35:0]   fixTo_990_dout;
  wire       [35:0]   fixTo_991_dout;
  wire       [17:0]   fixTo_992_dout;
  wire       [17:0]   fixTo_993_dout;
  wire       [17:0]   fixTo_994_dout;
  wire       [17:0]   fixTo_995_dout;
  wire       [35:0]   fixTo_996_dout;
  wire       [35:0]   fixTo_997_dout;
  wire       [17:0]   fixTo_998_dout;
  wire       [17:0]   fixTo_999_dout;
  wire       [17:0]   fixTo_1000_dout;
  wire       [17:0]   fixTo_1001_dout;
  wire       [35:0]   fixTo_1002_dout;
  wire       [35:0]   fixTo_1003_dout;
  wire       [17:0]   fixTo_1004_dout;
  wire       [17:0]   fixTo_1005_dout;
  wire       [17:0]   fixTo_1006_dout;
  wire       [17:0]   fixTo_1007_dout;
  wire       [35:0]   fixTo_1008_dout;
  wire       [35:0]   fixTo_1009_dout;
  wire       [17:0]   fixTo_1010_dout;
  wire       [17:0]   fixTo_1011_dout;
  wire       [17:0]   fixTo_1012_dout;
  wire       [17:0]   fixTo_1013_dout;
  wire       [35:0]   fixTo_1014_dout;
  wire       [35:0]   fixTo_1015_dout;
  wire       [17:0]   fixTo_1016_dout;
  wire       [17:0]   fixTo_1017_dout;
  wire       [17:0]   fixTo_1018_dout;
  wire       [17:0]   fixTo_1019_dout;
  wire       [35:0]   fixTo_1020_dout;
  wire       [35:0]   fixTo_1021_dout;
  wire       [17:0]   fixTo_1022_dout;
  wire       [17:0]   fixTo_1023_dout;
  wire       [17:0]   fixTo_1024_dout;
  wire       [17:0]   fixTo_1025_dout;
  wire       [35:0]   fixTo_1026_dout;
  wire       [35:0]   fixTo_1027_dout;
  wire       [17:0]   fixTo_1028_dout;
  wire       [17:0]   fixTo_1029_dout;
  wire       [17:0]   fixTo_1030_dout;
  wire       [17:0]   fixTo_1031_dout;
  wire       [35:0]   fixTo_1032_dout;
  wire       [35:0]   fixTo_1033_dout;
  wire       [17:0]   fixTo_1034_dout;
  wire       [17:0]   fixTo_1035_dout;
  wire       [17:0]   fixTo_1036_dout;
  wire       [17:0]   fixTo_1037_dout;
  wire       [35:0]   fixTo_1038_dout;
  wire       [35:0]   fixTo_1039_dout;
  wire       [17:0]   fixTo_1040_dout;
  wire       [17:0]   fixTo_1041_dout;
  wire       [17:0]   fixTo_1042_dout;
  wire       [17:0]   fixTo_1043_dout;
  wire       [35:0]   fixTo_1044_dout;
  wire       [35:0]   fixTo_1045_dout;
  wire       [17:0]   fixTo_1046_dout;
  wire       [17:0]   fixTo_1047_dout;
  wire       [17:0]   fixTo_1048_dout;
  wire       [17:0]   fixTo_1049_dout;
  wire       [35:0]   fixTo_1050_dout;
  wire       [35:0]   fixTo_1051_dout;
  wire       [17:0]   fixTo_1052_dout;
  wire       [17:0]   fixTo_1053_dout;
  wire       [17:0]   fixTo_1054_dout;
  wire       [17:0]   fixTo_1055_dout;
  wire       [35:0]   fixTo_1056_dout;
  wire       [35:0]   fixTo_1057_dout;
  wire       [17:0]   fixTo_1058_dout;
  wire       [17:0]   fixTo_1059_dout;
  wire       [17:0]   fixTo_1060_dout;
  wire       [17:0]   fixTo_1061_dout;
  wire       [35:0]   fixTo_1062_dout;
  wire       [35:0]   fixTo_1063_dout;
  wire       [17:0]   fixTo_1064_dout;
  wire       [17:0]   fixTo_1065_dout;
  wire       [17:0]   fixTo_1066_dout;
  wire       [17:0]   fixTo_1067_dout;
  wire       [35:0]   fixTo_1068_dout;
  wire       [35:0]   fixTo_1069_dout;
  wire       [17:0]   fixTo_1070_dout;
  wire       [17:0]   fixTo_1071_dout;
  wire       [17:0]   fixTo_1072_dout;
  wire       [17:0]   fixTo_1073_dout;
  wire       [35:0]   fixTo_1074_dout;
  wire       [35:0]   fixTo_1075_dout;
  wire       [17:0]   fixTo_1076_dout;
  wire       [17:0]   fixTo_1077_dout;
  wire       [17:0]   fixTo_1078_dout;
  wire       [17:0]   fixTo_1079_dout;
  wire       [35:0]   fixTo_1080_dout;
  wire       [35:0]   fixTo_1081_dout;
  wire       [17:0]   fixTo_1082_dout;
  wire       [17:0]   fixTo_1083_dout;
  wire       [17:0]   fixTo_1084_dout;
  wire       [17:0]   fixTo_1085_dout;
  wire       [35:0]   fixTo_1086_dout;
  wire       [35:0]   fixTo_1087_dout;
  wire       [17:0]   fixTo_1088_dout;
  wire       [17:0]   fixTo_1089_dout;
  wire       [17:0]   fixTo_1090_dout;
  wire       [17:0]   fixTo_1091_dout;
  wire       [35:0]   fixTo_1092_dout;
  wire       [35:0]   fixTo_1093_dout;
  wire       [17:0]   fixTo_1094_dout;
  wire       [17:0]   fixTo_1095_dout;
  wire       [17:0]   fixTo_1096_dout;
  wire       [17:0]   fixTo_1097_dout;
  wire       [35:0]   fixTo_1098_dout;
  wire       [35:0]   fixTo_1099_dout;
  wire       [17:0]   fixTo_1100_dout;
  wire       [17:0]   fixTo_1101_dout;
  wire       [17:0]   fixTo_1102_dout;
  wire       [17:0]   fixTo_1103_dout;
  wire       [35:0]   fixTo_1104_dout;
  wire       [35:0]   fixTo_1105_dout;
  wire       [17:0]   fixTo_1106_dout;
  wire       [17:0]   fixTo_1107_dout;
  wire       [17:0]   fixTo_1108_dout;
  wire       [17:0]   fixTo_1109_dout;
  wire       [35:0]   fixTo_1110_dout;
  wire       [35:0]   fixTo_1111_dout;
  wire       [17:0]   fixTo_1112_dout;
  wire       [17:0]   fixTo_1113_dout;
  wire       [17:0]   fixTo_1114_dout;
  wire       [17:0]   fixTo_1115_dout;
  wire       [35:0]   fixTo_1116_dout;
  wire       [35:0]   fixTo_1117_dout;
  wire       [17:0]   fixTo_1118_dout;
  wire       [17:0]   fixTo_1119_dout;
  wire       [17:0]   fixTo_1120_dout;
  wire       [17:0]   fixTo_1121_dout;
  wire       [35:0]   fixTo_1122_dout;
  wire       [35:0]   fixTo_1123_dout;
  wire       [17:0]   fixTo_1124_dout;
  wire       [17:0]   fixTo_1125_dout;
  wire       [17:0]   fixTo_1126_dout;
  wire       [17:0]   fixTo_1127_dout;
  wire       [35:0]   fixTo_1128_dout;
  wire       [35:0]   fixTo_1129_dout;
  wire       [17:0]   fixTo_1130_dout;
  wire       [17:0]   fixTo_1131_dout;
  wire       [17:0]   fixTo_1132_dout;
  wire       [17:0]   fixTo_1133_dout;
  wire       [35:0]   fixTo_1134_dout;
  wire       [35:0]   fixTo_1135_dout;
  wire       [17:0]   fixTo_1136_dout;
  wire       [17:0]   fixTo_1137_dout;
  wire       [17:0]   fixTo_1138_dout;
  wire       [17:0]   fixTo_1139_dout;
  wire       [35:0]   fixTo_1140_dout;
  wire       [35:0]   fixTo_1141_dout;
  wire       [17:0]   fixTo_1142_dout;
  wire       [17:0]   fixTo_1143_dout;
  wire       [17:0]   fixTo_1144_dout;
  wire       [17:0]   fixTo_1145_dout;
  wire       [35:0]   fixTo_1146_dout;
  wire       [35:0]   fixTo_1147_dout;
  wire       [17:0]   fixTo_1148_dout;
  wire       [17:0]   fixTo_1149_dout;
  wire       [17:0]   fixTo_1150_dout;
  wire       [17:0]   fixTo_1151_dout;
  wire       [17:0]   _zz_2113;
  wire       [35:0]   _zz_2114;
  wire       [35:0]   _zz_2115;
  wire       [17:0]   _zz_2116;
  wire       [35:0]   _zz_2117;
  wire       [35:0]   _zz_2118;
  wire       [35:0]   _zz_2119;
  wire       [17:0]   _zz_2120;
  wire       [35:0]   _zz_2121;
  wire       [35:0]   _zz_2122;
  wire       [35:0]   _zz_2123;
  wire       [35:0]   _zz_2124;
  wire       [35:0]   _zz_2125;
  wire       [35:0]   _zz_2126;
  wire       [26:0]   _zz_2127;
  wire       [35:0]   _zz_2128;
  wire       [17:0]   _zz_2129;
  wire       [35:0]   _zz_2130;
  wire       [35:0]   _zz_2131;
  wire       [35:0]   _zz_2132;
  wire       [35:0]   _zz_2133;
  wire       [35:0]   _zz_2134;
  wire       [26:0]   _zz_2135;
  wire       [35:0]   _zz_2136;
  wire       [17:0]   _zz_2137;
  wire       [35:0]   _zz_2138;
  wire       [35:0]   _zz_2139;
  wire       [35:0]   _zz_2140;
  wire       [35:0]   _zz_2141;
  wire       [35:0]   _zz_2142;
  wire       [26:0]   _zz_2143;
  wire       [35:0]   _zz_2144;
  wire       [17:0]   _zz_2145;
  wire       [35:0]   _zz_2146;
  wire       [35:0]   _zz_2147;
  wire       [35:0]   _zz_2148;
  wire       [35:0]   _zz_2149;
  wire       [35:0]   _zz_2150;
  wire       [26:0]   _zz_2151;
  wire       [35:0]   _zz_2152;
  wire       [17:0]   _zz_2153;
  wire       [17:0]   _zz_2154;
  wire       [35:0]   _zz_2155;
  wire       [35:0]   _zz_2156;
  wire       [17:0]   _zz_2157;
  wire       [35:0]   _zz_2158;
  wire       [35:0]   _zz_2159;
  wire       [35:0]   _zz_2160;
  wire       [17:0]   _zz_2161;
  wire       [35:0]   _zz_2162;
  wire       [35:0]   _zz_2163;
  wire       [35:0]   _zz_2164;
  wire       [35:0]   _zz_2165;
  wire       [35:0]   _zz_2166;
  wire       [35:0]   _zz_2167;
  wire       [26:0]   _zz_2168;
  wire       [35:0]   _zz_2169;
  wire       [17:0]   _zz_2170;
  wire       [35:0]   _zz_2171;
  wire       [35:0]   _zz_2172;
  wire       [35:0]   _zz_2173;
  wire       [35:0]   _zz_2174;
  wire       [35:0]   _zz_2175;
  wire       [26:0]   _zz_2176;
  wire       [35:0]   _zz_2177;
  wire       [17:0]   _zz_2178;
  wire       [35:0]   _zz_2179;
  wire       [35:0]   _zz_2180;
  wire       [35:0]   _zz_2181;
  wire       [35:0]   _zz_2182;
  wire       [35:0]   _zz_2183;
  wire       [26:0]   _zz_2184;
  wire       [35:0]   _zz_2185;
  wire       [17:0]   _zz_2186;
  wire       [35:0]   _zz_2187;
  wire       [35:0]   _zz_2188;
  wire       [35:0]   _zz_2189;
  wire       [35:0]   _zz_2190;
  wire       [35:0]   _zz_2191;
  wire       [26:0]   _zz_2192;
  wire       [35:0]   _zz_2193;
  wire       [17:0]   _zz_2194;
  wire       [17:0]   _zz_2195;
  wire       [35:0]   _zz_2196;
  wire       [35:0]   _zz_2197;
  wire       [17:0]   _zz_2198;
  wire       [35:0]   _zz_2199;
  wire       [35:0]   _zz_2200;
  wire       [35:0]   _zz_2201;
  wire       [17:0]   _zz_2202;
  wire       [35:0]   _zz_2203;
  wire       [35:0]   _zz_2204;
  wire       [35:0]   _zz_2205;
  wire       [35:0]   _zz_2206;
  wire       [35:0]   _zz_2207;
  wire       [35:0]   _zz_2208;
  wire       [26:0]   _zz_2209;
  wire       [35:0]   _zz_2210;
  wire       [17:0]   _zz_2211;
  wire       [35:0]   _zz_2212;
  wire       [35:0]   _zz_2213;
  wire       [35:0]   _zz_2214;
  wire       [35:0]   _zz_2215;
  wire       [35:0]   _zz_2216;
  wire       [26:0]   _zz_2217;
  wire       [35:0]   _zz_2218;
  wire       [17:0]   _zz_2219;
  wire       [35:0]   _zz_2220;
  wire       [35:0]   _zz_2221;
  wire       [35:0]   _zz_2222;
  wire       [35:0]   _zz_2223;
  wire       [35:0]   _zz_2224;
  wire       [26:0]   _zz_2225;
  wire       [35:0]   _zz_2226;
  wire       [17:0]   _zz_2227;
  wire       [35:0]   _zz_2228;
  wire       [35:0]   _zz_2229;
  wire       [35:0]   _zz_2230;
  wire       [35:0]   _zz_2231;
  wire       [35:0]   _zz_2232;
  wire       [26:0]   _zz_2233;
  wire       [35:0]   _zz_2234;
  wire       [17:0]   _zz_2235;
  wire       [17:0]   _zz_2236;
  wire       [35:0]   _zz_2237;
  wire       [35:0]   _zz_2238;
  wire       [17:0]   _zz_2239;
  wire       [35:0]   _zz_2240;
  wire       [35:0]   _zz_2241;
  wire       [35:0]   _zz_2242;
  wire       [17:0]   _zz_2243;
  wire       [35:0]   _zz_2244;
  wire       [35:0]   _zz_2245;
  wire       [35:0]   _zz_2246;
  wire       [35:0]   _zz_2247;
  wire       [35:0]   _zz_2248;
  wire       [35:0]   _zz_2249;
  wire       [26:0]   _zz_2250;
  wire       [35:0]   _zz_2251;
  wire       [17:0]   _zz_2252;
  wire       [35:0]   _zz_2253;
  wire       [35:0]   _zz_2254;
  wire       [35:0]   _zz_2255;
  wire       [35:0]   _zz_2256;
  wire       [35:0]   _zz_2257;
  wire       [26:0]   _zz_2258;
  wire       [35:0]   _zz_2259;
  wire       [17:0]   _zz_2260;
  wire       [35:0]   _zz_2261;
  wire       [35:0]   _zz_2262;
  wire       [35:0]   _zz_2263;
  wire       [35:0]   _zz_2264;
  wire       [35:0]   _zz_2265;
  wire       [26:0]   _zz_2266;
  wire       [35:0]   _zz_2267;
  wire       [17:0]   _zz_2268;
  wire       [35:0]   _zz_2269;
  wire       [35:0]   _zz_2270;
  wire       [35:0]   _zz_2271;
  wire       [35:0]   _zz_2272;
  wire       [35:0]   _zz_2273;
  wire       [26:0]   _zz_2274;
  wire       [35:0]   _zz_2275;
  wire       [17:0]   _zz_2276;
  wire       [17:0]   _zz_2277;
  wire       [35:0]   _zz_2278;
  wire       [35:0]   _zz_2279;
  wire       [17:0]   _zz_2280;
  wire       [35:0]   _zz_2281;
  wire       [35:0]   _zz_2282;
  wire       [35:0]   _zz_2283;
  wire       [17:0]   _zz_2284;
  wire       [35:0]   _zz_2285;
  wire       [35:0]   _zz_2286;
  wire       [35:0]   _zz_2287;
  wire       [35:0]   _zz_2288;
  wire       [35:0]   _zz_2289;
  wire       [35:0]   _zz_2290;
  wire       [26:0]   _zz_2291;
  wire       [35:0]   _zz_2292;
  wire       [17:0]   _zz_2293;
  wire       [35:0]   _zz_2294;
  wire       [35:0]   _zz_2295;
  wire       [35:0]   _zz_2296;
  wire       [35:0]   _zz_2297;
  wire       [35:0]   _zz_2298;
  wire       [26:0]   _zz_2299;
  wire       [35:0]   _zz_2300;
  wire       [17:0]   _zz_2301;
  wire       [35:0]   _zz_2302;
  wire       [35:0]   _zz_2303;
  wire       [35:0]   _zz_2304;
  wire       [35:0]   _zz_2305;
  wire       [35:0]   _zz_2306;
  wire       [26:0]   _zz_2307;
  wire       [35:0]   _zz_2308;
  wire       [17:0]   _zz_2309;
  wire       [35:0]   _zz_2310;
  wire       [35:0]   _zz_2311;
  wire       [35:0]   _zz_2312;
  wire       [35:0]   _zz_2313;
  wire       [35:0]   _zz_2314;
  wire       [26:0]   _zz_2315;
  wire       [35:0]   _zz_2316;
  wire       [17:0]   _zz_2317;
  wire       [17:0]   _zz_2318;
  wire       [35:0]   _zz_2319;
  wire       [35:0]   _zz_2320;
  wire       [17:0]   _zz_2321;
  wire       [35:0]   _zz_2322;
  wire       [35:0]   _zz_2323;
  wire       [35:0]   _zz_2324;
  wire       [17:0]   _zz_2325;
  wire       [35:0]   _zz_2326;
  wire       [35:0]   _zz_2327;
  wire       [35:0]   _zz_2328;
  wire       [35:0]   _zz_2329;
  wire       [35:0]   _zz_2330;
  wire       [35:0]   _zz_2331;
  wire       [26:0]   _zz_2332;
  wire       [35:0]   _zz_2333;
  wire       [17:0]   _zz_2334;
  wire       [35:0]   _zz_2335;
  wire       [35:0]   _zz_2336;
  wire       [35:0]   _zz_2337;
  wire       [35:0]   _zz_2338;
  wire       [35:0]   _zz_2339;
  wire       [26:0]   _zz_2340;
  wire       [35:0]   _zz_2341;
  wire       [17:0]   _zz_2342;
  wire       [35:0]   _zz_2343;
  wire       [35:0]   _zz_2344;
  wire       [35:0]   _zz_2345;
  wire       [35:0]   _zz_2346;
  wire       [35:0]   _zz_2347;
  wire       [26:0]   _zz_2348;
  wire       [35:0]   _zz_2349;
  wire       [17:0]   _zz_2350;
  wire       [35:0]   _zz_2351;
  wire       [35:0]   _zz_2352;
  wire       [35:0]   _zz_2353;
  wire       [35:0]   _zz_2354;
  wire       [35:0]   _zz_2355;
  wire       [26:0]   _zz_2356;
  wire       [35:0]   _zz_2357;
  wire       [17:0]   _zz_2358;
  wire       [17:0]   _zz_2359;
  wire       [35:0]   _zz_2360;
  wire       [35:0]   _zz_2361;
  wire       [17:0]   _zz_2362;
  wire       [35:0]   _zz_2363;
  wire       [35:0]   _zz_2364;
  wire       [35:0]   _zz_2365;
  wire       [17:0]   _zz_2366;
  wire       [35:0]   _zz_2367;
  wire       [35:0]   _zz_2368;
  wire       [35:0]   _zz_2369;
  wire       [35:0]   _zz_2370;
  wire       [35:0]   _zz_2371;
  wire       [35:0]   _zz_2372;
  wire       [26:0]   _zz_2373;
  wire       [35:0]   _zz_2374;
  wire       [17:0]   _zz_2375;
  wire       [35:0]   _zz_2376;
  wire       [35:0]   _zz_2377;
  wire       [35:0]   _zz_2378;
  wire       [35:0]   _zz_2379;
  wire       [35:0]   _zz_2380;
  wire       [26:0]   _zz_2381;
  wire       [35:0]   _zz_2382;
  wire       [17:0]   _zz_2383;
  wire       [35:0]   _zz_2384;
  wire       [35:0]   _zz_2385;
  wire       [35:0]   _zz_2386;
  wire       [35:0]   _zz_2387;
  wire       [35:0]   _zz_2388;
  wire       [26:0]   _zz_2389;
  wire       [35:0]   _zz_2390;
  wire       [17:0]   _zz_2391;
  wire       [35:0]   _zz_2392;
  wire       [35:0]   _zz_2393;
  wire       [35:0]   _zz_2394;
  wire       [35:0]   _zz_2395;
  wire       [35:0]   _zz_2396;
  wire       [26:0]   _zz_2397;
  wire       [35:0]   _zz_2398;
  wire       [17:0]   _zz_2399;
  wire       [17:0]   _zz_2400;
  wire       [35:0]   _zz_2401;
  wire       [35:0]   _zz_2402;
  wire       [17:0]   _zz_2403;
  wire       [35:0]   _zz_2404;
  wire       [35:0]   _zz_2405;
  wire       [35:0]   _zz_2406;
  wire       [17:0]   _zz_2407;
  wire       [35:0]   _zz_2408;
  wire       [35:0]   _zz_2409;
  wire       [35:0]   _zz_2410;
  wire       [35:0]   _zz_2411;
  wire       [35:0]   _zz_2412;
  wire       [35:0]   _zz_2413;
  wire       [26:0]   _zz_2414;
  wire       [35:0]   _zz_2415;
  wire       [17:0]   _zz_2416;
  wire       [35:0]   _zz_2417;
  wire       [35:0]   _zz_2418;
  wire       [35:0]   _zz_2419;
  wire       [35:0]   _zz_2420;
  wire       [35:0]   _zz_2421;
  wire       [26:0]   _zz_2422;
  wire       [35:0]   _zz_2423;
  wire       [17:0]   _zz_2424;
  wire       [35:0]   _zz_2425;
  wire       [35:0]   _zz_2426;
  wire       [35:0]   _zz_2427;
  wire       [35:0]   _zz_2428;
  wire       [35:0]   _zz_2429;
  wire       [26:0]   _zz_2430;
  wire       [35:0]   _zz_2431;
  wire       [17:0]   _zz_2432;
  wire       [35:0]   _zz_2433;
  wire       [35:0]   _zz_2434;
  wire       [35:0]   _zz_2435;
  wire       [35:0]   _zz_2436;
  wire       [35:0]   _zz_2437;
  wire       [26:0]   _zz_2438;
  wire       [35:0]   _zz_2439;
  wire       [17:0]   _zz_2440;
  wire       [17:0]   _zz_2441;
  wire       [35:0]   _zz_2442;
  wire       [35:0]   _zz_2443;
  wire       [17:0]   _zz_2444;
  wire       [35:0]   _zz_2445;
  wire       [35:0]   _zz_2446;
  wire       [35:0]   _zz_2447;
  wire       [17:0]   _zz_2448;
  wire       [35:0]   _zz_2449;
  wire       [35:0]   _zz_2450;
  wire       [35:0]   _zz_2451;
  wire       [35:0]   _zz_2452;
  wire       [35:0]   _zz_2453;
  wire       [35:0]   _zz_2454;
  wire       [26:0]   _zz_2455;
  wire       [35:0]   _zz_2456;
  wire       [17:0]   _zz_2457;
  wire       [35:0]   _zz_2458;
  wire       [35:0]   _zz_2459;
  wire       [35:0]   _zz_2460;
  wire       [35:0]   _zz_2461;
  wire       [35:0]   _zz_2462;
  wire       [26:0]   _zz_2463;
  wire       [35:0]   _zz_2464;
  wire       [17:0]   _zz_2465;
  wire       [35:0]   _zz_2466;
  wire       [35:0]   _zz_2467;
  wire       [35:0]   _zz_2468;
  wire       [35:0]   _zz_2469;
  wire       [35:0]   _zz_2470;
  wire       [26:0]   _zz_2471;
  wire       [35:0]   _zz_2472;
  wire       [17:0]   _zz_2473;
  wire       [35:0]   _zz_2474;
  wire       [35:0]   _zz_2475;
  wire       [35:0]   _zz_2476;
  wire       [35:0]   _zz_2477;
  wire       [35:0]   _zz_2478;
  wire       [26:0]   _zz_2479;
  wire       [35:0]   _zz_2480;
  wire       [17:0]   _zz_2481;
  wire       [17:0]   _zz_2482;
  wire       [35:0]   _zz_2483;
  wire       [35:0]   _zz_2484;
  wire       [17:0]   _zz_2485;
  wire       [35:0]   _zz_2486;
  wire       [35:0]   _zz_2487;
  wire       [35:0]   _zz_2488;
  wire       [17:0]   _zz_2489;
  wire       [35:0]   _zz_2490;
  wire       [35:0]   _zz_2491;
  wire       [35:0]   _zz_2492;
  wire       [35:0]   _zz_2493;
  wire       [35:0]   _zz_2494;
  wire       [35:0]   _zz_2495;
  wire       [26:0]   _zz_2496;
  wire       [35:0]   _zz_2497;
  wire       [17:0]   _zz_2498;
  wire       [35:0]   _zz_2499;
  wire       [35:0]   _zz_2500;
  wire       [35:0]   _zz_2501;
  wire       [35:0]   _zz_2502;
  wire       [35:0]   _zz_2503;
  wire       [26:0]   _zz_2504;
  wire       [35:0]   _zz_2505;
  wire       [17:0]   _zz_2506;
  wire       [35:0]   _zz_2507;
  wire       [35:0]   _zz_2508;
  wire       [35:0]   _zz_2509;
  wire       [35:0]   _zz_2510;
  wire       [35:0]   _zz_2511;
  wire       [26:0]   _zz_2512;
  wire       [35:0]   _zz_2513;
  wire       [17:0]   _zz_2514;
  wire       [35:0]   _zz_2515;
  wire       [35:0]   _zz_2516;
  wire       [35:0]   _zz_2517;
  wire       [35:0]   _zz_2518;
  wire       [35:0]   _zz_2519;
  wire       [26:0]   _zz_2520;
  wire       [35:0]   _zz_2521;
  wire       [17:0]   _zz_2522;
  wire       [17:0]   _zz_2523;
  wire       [35:0]   _zz_2524;
  wire       [35:0]   _zz_2525;
  wire       [17:0]   _zz_2526;
  wire       [35:0]   _zz_2527;
  wire       [35:0]   _zz_2528;
  wire       [35:0]   _zz_2529;
  wire       [17:0]   _zz_2530;
  wire       [35:0]   _zz_2531;
  wire       [35:0]   _zz_2532;
  wire       [35:0]   _zz_2533;
  wire       [35:0]   _zz_2534;
  wire       [35:0]   _zz_2535;
  wire       [35:0]   _zz_2536;
  wire       [26:0]   _zz_2537;
  wire       [35:0]   _zz_2538;
  wire       [17:0]   _zz_2539;
  wire       [35:0]   _zz_2540;
  wire       [35:0]   _zz_2541;
  wire       [35:0]   _zz_2542;
  wire       [35:0]   _zz_2543;
  wire       [35:0]   _zz_2544;
  wire       [26:0]   _zz_2545;
  wire       [35:0]   _zz_2546;
  wire       [17:0]   _zz_2547;
  wire       [35:0]   _zz_2548;
  wire       [35:0]   _zz_2549;
  wire       [35:0]   _zz_2550;
  wire       [35:0]   _zz_2551;
  wire       [35:0]   _zz_2552;
  wire       [26:0]   _zz_2553;
  wire       [35:0]   _zz_2554;
  wire       [17:0]   _zz_2555;
  wire       [35:0]   _zz_2556;
  wire       [35:0]   _zz_2557;
  wire       [35:0]   _zz_2558;
  wire       [35:0]   _zz_2559;
  wire       [35:0]   _zz_2560;
  wire       [26:0]   _zz_2561;
  wire       [35:0]   _zz_2562;
  wire       [17:0]   _zz_2563;
  wire       [17:0]   _zz_2564;
  wire       [35:0]   _zz_2565;
  wire       [35:0]   _zz_2566;
  wire       [17:0]   _zz_2567;
  wire       [35:0]   _zz_2568;
  wire       [35:0]   _zz_2569;
  wire       [35:0]   _zz_2570;
  wire       [17:0]   _zz_2571;
  wire       [35:0]   _zz_2572;
  wire       [35:0]   _zz_2573;
  wire       [35:0]   _zz_2574;
  wire       [35:0]   _zz_2575;
  wire       [35:0]   _zz_2576;
  wire       [35:0]   _zz_2577;
  wire       [26:0]   _zz_2578;
  wire       [35:0]   _zz_2579;
  wire       [17:0]   _zz_2580;
  wire       [35:0]   _zz_2581;
  wire       [35:0]   _zz_2582;
  wire       [35:0]   _zz_2583;
  wire       [35:0]   _zz_2584;
  wire       [35:0]   _zz_2585;
  wire       [26:0]   _zz_2586;
  wire       [35:0]   _zz_2587;
  wire       [17:0]   _zz_2588;
  wire       [35:0]   _zz_2589;
  wire       [35:0]   _zz_2590;
  wire       [35:0]   _zz_2591;
  wire       [35:0]   _zz_2592;
  wire       [35:0]   _zz_2593;
  wire       [26:0]   _zz_2594;
  wire       [35:0]   _zz_2595;
  wire       [17:0]   _zz_2596;
  wire       [35:0]   _zz_2597;
  wire       [35:0]   _zz_2598;
  wire       [35:0]   _zz_2599;
  wire       [35:0]   _zz_2600;
  wire       [35:0]   _zz_2601;
  wire       [26:0]   _zz_2602;
  wire       [35:0]   _zz_2603;
  wire       [17:0]   _zz_2604;
  wire       [17:0]   _zz_2605;
  wire       [35:0]   _zz_2606;
  wire       [35:0]   _zz_2607;
  wire       [17:0]   _zz_2608;
  wire       [35:0]   _zz_2609;
  wire       [35:0]   _zz_2610;
  wire       [35:0]   _zz_2611;
  wire       [17:0]   _zz_2612;
  wire       [35:0]   _zz_2613;
  wire       [35:0]   _zz_2614;
  wire       [35:0]   _zz_2615;
  wire       [35:0]   _zz_2616;
  wire       [35:0]   _zz_2617;
  wire       [35:0]   _zz_2618;
  wire       [26:0]   _zz_2619;
  wire       [35:0]   _zz_2620;
  wire       [17:0]   _zz_2621;
  wire       [35:0]   _zz_2622;
  wire       [35:0]   _zz_2623;
  wire       [35:0]   _zz_2624;
  wire       [35:0]   _zz_2625;
  wire       [35:0]   _zz_2626;
  wire       [26:0]   _zz_2627;
  wire       [35:0]   _zz_2628;
  wire       [17:0]   _zz_2629;
  wire       [35:0]   _zz_2630;
  wire       [35:0]   _zz_2631;
  wire       [35:0]   _zz_2632;
  wire       [35:0]   _zz_2633;
  wire       [35:0]   _zz_2634;
  wire       [26:0]   _zz_2635;
  wire       [35:0]   _zz_2636;
  wire       [17:0]   _zz_2637;
  wire       [35:0]   _zz_2638;
  wire       [35:0]   _zz_2639;
  wire       [35:0]   _zz_2640;
  wire       [35:0]   _zz_2641;
  wire       [35:0]   _zz_2642;
  wire       [26:0]   _zz_2643;
  wire       [35:0]   _zz_2644;
  wire       [17:0]   _zz_2645;
  wire       [17:0]   _zz_2646;
  wire       [35:0]   _zz_2647;
  wire       [35:0]   _zz_2648;
  wire       [17:0]   _zz_2649;
  wire       [35:0]   _zz_2650;
  wire       [35:0]   _zz_2651;
  wire       [35:0]   _zz_2652;
  wire       [17:0]   _zz_2653;
  wire       [35:0]   _zz_2654;
  wire       [35:0]   _zz_2655;
  wire       [35:0]   _zz_2656;
  wire       [35:0]   _zz_2657;
  wire       [35:0]   _zz_2658;
  wire       [35:0]   _zz_2659;
  wire       [26:0]   _zz_2660;
  wire       [35:0]   _zz_2661;
  wire       [17:0]   _zz_2662;
  wire       [35:0]   _zz_2663;
  wire       [35:0]   _zz_2664;
  wire       [35:0]   _zz_2665;
  wire       [35:0]   _zz_2666;
  wire       [35:0]   _zz_2667;
  wire       [26:0]   _zz_2668;
  wire       [35:0]   _zz_2669;
  wire       [17:0]   _zz_2670;
  wire       [35:0]   _zz_2671;
  wire       [35:0]   _zz_2672;
  wire       [35:0]   _zz_2673;
  wire       [35:0]   _zz_2674;
  wire       [35:0]   _zz_2675;
  wire       [26:0]   _zz_2676;
  wire       [35:0]   _zz_2677;
  wire       [17:0]   _zz_2678;
  wire       [35:0]   _zz_2679;
  wire       [35:0]   _zz_2680;
  wire       [35:0]   _zz_2681;
  wire       [35:0]   _zz_2682;
  wire       [35:0]   _zz_2683;
  wire       [26:0]   _zz_2684;
  wire       [35:0]   _zz_2685;
  wire       [17:0]   _zz_2686;
  wire       [17:0]   _zz_2687;
  wire       [35:0]   _zz_2688;
  wire       [35:0]   _zz_2689;
  wire       [17:0]   _zz_2690;
  wire       [35:0]   _zz_2691;
  wire       [35:0]   _zz_2692;
  wire       [35:0]   _zz_2693;
  wire       [17:0]   _zz_2694;
  wire       [35:0]   _zz_2695;
  wire       [35:0]   _zz_2696;
  wire       [35:0]   _zz_2697;
  wire       [35:0]   _zz_2698;
  wire       [35:0]   _zz_2699;
  wire       [35:0]   _zz_2700;
  wire       [26:0]   _zz_2701;
  wire       [35:0]   _zz_2702;
  wire       [17:0]   _zz_2703;
  wire       [35:0]   _zz_2704;
  wire       [35:0]   _zz_2705;
  wire       [35:0]   _zz_2706;
  wire       [35:0]   _zz_2707;
  wire       [35:0]   _zz_2708;
  wire       [26:0]   _zz_2709;
  wire       [35:0]   _zz_2710;
  wire       [17:0]   _zz_2711;
  wire       [35:0]   _zz_2712;
  wire       [35:0]   _zz_2713;
  wire       [35:0]   _zz_2714;
  wire       [35:0]   _zz_2715;
  wire       [35:0]   _zz_2716;
  wire       [26:0]   _zz_2717;
  wire       [35:0]   _zz_2718;
  wire       [17:0]   _zz_2719;
  wire       [35:0]   _zz_2720;
  wire       [35:0]   _zz_2721;
  wire       [35:0]   _zz_2722;
  wire       [35:0]   _zz_2723;
  wire       [35:0]   _zz_2724;
  wire       [26:0]   _zz_2725;
  wire       [35:0]   _zz_2726;
  wire       [17:0]   _zz_2727;
  wire       [17:0]   _zz_2728;
  wire       [35:0]   _zz_2729;
  wire       [35:0]   _zz_2730;
  wire       [17:0]   _zz_2731;
  wire       [35:0]   _zz_2732;
  wire       [35:0]   _zz_2733;
  wire       [35:0]   _zz_2734;
  wire       [17:0]   _zz_2735;
  wire       [35:0]   _zz_2736;
  wire       [35:0]   _zz_2737;
  wire       [35:0]   _zz_2738;
  wire       [35:0]   _zz_2739;
  wire       [35:0]   _zz_2740;
  wire       [35:0]   _zz_2741;
  wire       [26:0]   _zz_2742;
  wire       [35:0]   _zz_2743;
  wire       [17:0]   _zz_2744;
  wire       [35:0]   _zz_2745;
  wire       [35:0]   _zz_2746;
  wire       [35:0]   _zz_2747;
  wire       [35:0]   _zz_2748;
  wire       [35:0]   _zz_2749;
  wire       [26:0]   _zz_2750;
  wire       [35:0]   _zz_2751;
  wire       [17:0]   _zz_2752;
  wire       [35:0]   _zz_2753;
  wire       [35:0]   _zz_2754;
  wire       [35:0]   _zz_2755;
  wire       [35:0]   _zz_2756;
  wire       [35:0]   _zz_2757;
  wire       [26:0]   _zz_2758;
  wire       [35:0]   _zz_2759;
  wire       [17:0]   _zz_2760;
  wire       [35:0]   _zz_2761;
  wire       [35:0]   _zz_2762;
  wire       [35:0]   _zz_2763;
  wire       [35:0]   _zz_2764;
  wire       [35:0]   _zz_2765;
  wire       [26:0]   _zz_2766;
  wire       [35:0]   _zz_2767;
  wire       [17:0]   _zz_2768;
  wire       [17:0]   _zz_2769;
  wire       [35:0]   _zz_2770;
  wire       [35:0]   _zz_2771;
  wire       [17:0]   _zz_2772;
  wire       [35:0]   _zz_2773;
  wire       [35:0]   _zz_2774;
  wire       [35:0]   _zz_2775;
  wire       [17:0]   _zz_2776;
  wire       [35:0]   _zz_2777;
  wire       [35:0]   _zz_2778;
  wire       [35:0]   _zz_2779;
  wire       [35:0]   _zz_2780;
  wire       [35:0]   _zz_2781;
  wire       [35:0]   _zz_2782;
  wire       [26:0]   _zz_2783;
  wire       [35:0]   _zz_2784;
  wire       [17:0]   _zz_2785;
  wire       [35:0]   _zz_2786;
  wire       [35:0]   _zz_2787;
  wire       [35:0]   _zz_2788;
  wire       [35:0]   _zz_2789;
  wire       [35:0]   _zz_2790;
  wire       [26:0]   _zz_2791;
  wire       [35:0]   _zz_2792;
  wire       [17:0]   _zz_2793;
  wire       [35:0]   _zz_2794;
  wire       [35:0]   _zz_2795;
  wire       [35:0]   _zz_2796;
  wire       [35:0]   _zz_2797;
  wire       [35:0]   _zz_2798;
  wire       [26:0]   _zz_2799;
  wire       [35:0]   _zz_2800;
  wire       [17:0]   _zz_2801;
  wire       [35:0]   _zz_2802;
  wire       [35:0]   _zz_2803;
  wire       [35:0]   _zz_2804;
  wire       [35:0]   _zz_2805;
  wire       [35:0]   _zz_2806;
  wire       [26:0]   _zz_2807;
  wire       [35:0]   _zz_2808;
  wire       [17:0]   _zz_2809;
  wire       [17:0]   _zz_2810;
  wire       [35:0]   _zz_2811;
  wire       [35:0]   _zz_2812;
  wire       [17:0]   _zz_2813;
  wire       [35:0]   _zz_2814;
  wire       [35:0]   _zz_2815;
  wire       [35:0]   _zz_2816;
  wire       [17:0]   _zz_2817;
  wire       [35:0]   _zz_2818;
  wire       [35:0]   _zz_2819;
  wire       [35:0]   _zz_2820;
  wire       [35:0]   _zz_2821;
  wire       [35:0]   _zz_2822;
  wire       [35:0]   _zz_2823;
  wire       [26:0]   _zz_2824;
  wire       [35:0]   _zz_2825;
  wire       [17:0]   _zz_2826;
  wire       [35:0]   _zz_2827;
  wire       [35:0]   _zz_2828;
  wire       [35:0]   _zz_2829;
  wire       [35:0]   _zz_2830;
  wire       [35:0]   _zz_2831;
  wire       [26:0]   _zz_2832;
  wire       [35:0]   _zz_2833;
  wire       [17:0]   _zz_2834;
  wire       [35:0]   _zz_2835;
  wire       [35:0]   _zz_2836;
  wire       [35:0]   _zz_2837;
  wire       [35:0]   _zz_2838;
  wire       [35:0]   _zz_2839;
  wire       [26:0]   _zz_2840;
  wire       [35:0]   _zz_2841;
  wire       [17:0]   _zz_2842;
  wire       [35:0]   _zz_2843;
  wire       [35:0]   _zz_2844;
  wire       [35:0]   _zz_2845;
  wire       [35:0]   _zz_2846;
  wire       [35:0]   _zz_2847;
  wire       [26:0]   _zz_2848;
  wire       [35:0]   _zz_2849;
  wire       [17:0]   _zz_2850;
  wire       [17:0]   _zz_2851;
  wire       [35:0]   _zz_2852;
  wire       [35:0]   _zz_2853;
  wire       [17:0]   _zz_2854;
  wire       [35:0]   _zz_2855;
  wire       [35:0]   _zz_2856;
  wire       [35:0]   _zz_2857;
  wire       [17:0]   _zz_2858;
  wire       [35:0]   _zz_2859;
  wire       [35:0]   _zz_2860;
  wire       [35:0]   _zz_2861;
  wire       [35:0]   _zz_2862;
  wire       [35:0]   _zz_2863;
  wire       [35:0]   _zz_2864;
  wire       [26:0]   _zz_2865;
  wire       [35:0]   _zz_2866;
  wire       [17:0]   _zz_2867;
  wire       [35:0]   _zz_2868;
  wire       [35:0]   _zz_2869;
  wire       [35:0]   _zz_2870;
  wire       [35:0]   _zz_2871;
  wire       [35:0]   _zz_2872;
  wire       [26:0]   _zz_2873;
  wire       [35:0]   _zz_2874;
  wire       [17:0]   _zz_2875;
  wire       [35:0]   _zz_2876;
  wire       [35:0]   _zz_2877;
  wire       [35:0]   _zz_2878;
  wire       [35:0]   _zz_2879;
  wire       [35:0]   _zz_2880;
  wire       [26:0]   _zz_2881;
  wire       [35:0]   _zz_2882;
  wire       [17:0]   _zz_2883;
  wire       [35:0]   _zz_2884;
  wire       [35:0]   _zz_2885;
  wire       [35:0]   _zz_2886;
  wire       [35:0]   _zz_2887;
  wire       [35:0]   _zz_2888;
  wire       [26:0]   _zz_2889;
  wire       [35:0]   _zz_2890;
  wire       [17:0]   _zz_2891;
  wire       [17:0]   _zz_2892;
  wire       [35:0]   _zz_2893;
  wire       [35:0]   _zz_2894;
  wire       [17:0]   _zz_2895;
  wire       [35:0]   _zz_2896;
  wire       [35:0]   _zz_2897;
  wire       [35:0]   _zz_2898;
  wire       [17:0]   _zz_2899;
  wire       [35:0]   _zz_2900;
  wire       [35:0]   _zz_2901;
  wire       [35:0]   _zz_2902;
  wire       [35:0]   _zz_2903;
  wire       [35:0]   _zz_2904;
  wire       [35:0]   _zz_2905;
  wire       [26:0]   _zz_2906;
  wire       [35:0]   _zz_2907;
  wire       [17:0]   _zz_2908;
  wire       [35:0]   _zz_2909;
  wire       [35:0]   _zz_2910;
  wire       [35:0]   _zz_2911;
  wire       [35:0]   _zz_2912;
  wire       [35:0]   _zz_2913;
  wire       [26:0]   _zz_2914;
  wire       [35:0]   _zz_2915;
  wire       [17:0]   _zz_2916;
  wire       [35:0]   _zz_2917;
  wire       [35:0]   _zz_2918;
  wire       [35:0]   _zz_2919;
  wire       [35:0]   _zz_2920;
  wire       [35:0]   _zz_2921;
  wire       [26:0]   _zz_2922;
  wire       [35:0]   _zz_2923;
  wire       [17:0]   _zz_2924;
  wire       [35:0]   _zz_2925;
  wire       [35:0]   _zz_2926;
  wire       [35:0]   _zz_2927;
  wire       [35:0]   _zz_2928;
  wire       [35:0]   _zz_2929;
  wire       [26:0]   _zz_2930;
  wire       [35:0]   _zz_2931;
  wire       [17:0]   _zz_2932;
  wire       [17:0]   _zz_2933;
  wire       [35:0]   _zz_2934;
  wire       [35:0]   _zz_2935;
  wire       [17:0]   _zz_2936;
  wire       [35:0]   _zz_2937;
  wire       [35:0]   _zz_2938;
  wire       [35:0]   _zz_2939;
  wire       [17:0]   _zz_2940;
  wire       [35:0]   _zz_2941;
  wire       [35:0]   _zz_2942;
  wire       [35:0]   _zz_2943;
  wire       [35:0]   _zz_2944;
  wire       [35:0]   _zz_2945;
  wire       [35:0]   _zz_2946;
  wire       [26:0]   _zz_2947;
  wire       [35:0]   _zz_2948;
  wire       [17:0]   _zz_2949;
  wire       [35:0]   _zz_2950;
  wire       [35:0]   _zz_2951;
  wire       [35:0]   _zz_2952;
  wire       [35:0]   _zz_2953;
  wire       [35:0]   _zz_2954;
  wire       [26:0]   _zz_2955;
  wire       [35:0]   _zz_2956;
  wire       [17:0]   _zz_2957;
  wire       [35:0]   _zz_2958;
  wire       [35:0]   _zz_2959;
  wire       [35:0]   _zz_2960;
  wire       [35:0]   _zz_2961;
  wire       [35:0]   _zz_2962;
  wire       [26:0]   _zz_2963;
  wire       [35:0]   _zz_2964;
  wire       [17:0]   _zz_2965;
  wire       [35:0]   _zz_2966;
  wire       [35:0]   _zz_2967;
  wire       [35:0]   _zz_2968;
  wire       [35:0]   _zz_2969;
  wire       [35:0]   _zz_2970;
  wire       [26:0]   _zz_2971;
  wire       [35:0]   _zz_2972;
  wire       [17:0]   _zz_2973;
  wire       [17:0]   _zz_2974;
  wire       [35:0]   _zz_2975;
  wire       [35:0]   _zz_2976;
  wire       [17:0]   _zz_2977;
  wire       [35:0]   _zz_2978;
  wire       [35:0]   _zz_2979;
  wire       [35:0]   _zz_2980;
  wire       [17:0]   _zz_2981;
  wire       [35:0]   _zz_2982;
  wire       [35:0]   _zz_2983;
  wire       [35:0]   _zz_2984;
  wire       [35:0]   _zz_2985;
  wire       [35:0]   _zz_2986;
  wire       [35:0]   _zz_2987;
  wire       [26:0]   _zz_2988;
  wire       [35:0]   _zz_2989;
  wire       [17:0]   _zz_2990;
  wire       [35:0]   _zz_2991;
  wire       [35:0]   _zz_2992;
  wire       [35:0]   _zz_2993;
  wire       [35:0]   _zz_2994;
  wire       [35:0]   _zz_2995;
  wire       [26:0]   _zz_2996;
  wire       [35:0]   _zz_2997;
  wire       [17:0]   _zz_2998;
  wire       [35:0]   _zz_2999;
  wire       [35:0]   _zz_3000;
  wire       [35:0]   _zz_3001;
  wire       [35:0]   _zz_3002;
  wire       [35:0]   _zz_3003;
  wire       [26:0]   _zz_3004;
  wire       [35:0]   _zz_3005;
  wire       [17:0]   _zz_3006;
  wire       [35:0]   _zz_3007;
  wire       [35:0]   _zz_3008;
  wire       [35:0]   _zz_3009;
  wire       [35:0]   _zz_3010;
  wire       [35:0]   _zz_3011;
  wire       [26:0]   _zz_3012;
  wire       [35:0]   _zz_3013;
  wire       [17:0]   _zz_3014;
  wire       [17:0]   _zz_3015;
  wire       [35:0]   _zz_3016;
  wire       [35:0]   _zz_3017;
  wire       [17:0]   _zz_3018;
  wire       [35:0]   _zz_3019;
  wire       [35:0]   _zz_3020;
  wire       [35:0]   _zz_3021;
  wire       [17:0]   _zz_3022;
  wire       [35:0]   _zz_3023;
  wire       [35:0]   _zz_3024;
  wire       [35:0]   _zz_3025;
  wire       [35:0]   _zz_3026;
  wire       [35:0]   _zz_3027;
  wire       [35:0]   _zz_3028;
  wire       [26:0]   _zz_3029;
  wire       [35:0]   _zz_3030;
  wire       [17:0]   _zz_3031;
  wire       [35:0]   _zz_3032;
  wire       [35:0]   _zz_3033;
  wire       [35:0]   _zz_3034;
  wire       [35:0]   _zz_3035;
  wire       [35:0]   _zz_3036;
  wire       [26:0]   _zz_3037;
  wire       [35:0]   _zz_3038;
  wire       [17:0]   _zz_3039;
  wire       [35:0]   _zz_3040;
  wire       [35:0]   _zz_3041;
  wire       [35:0]   _zz_3042;
  wire       [35:0]   _zz_3043;
  wire       [35:0]   _zz_3044;
  wire       [26:0]   _zz_3045;
  wire       [35:0]   _zz_3046;
  wire       [17:0]   _zz_3047;
  wire       [35:0]   _zz_3048;
  wire       [35:0]   _zz_3049;
  wire       [35:0]   _zz_3050;
  wire       [35:0]   _zz_3051;
  wire       [35:0]   _zz_3052;
  wire       [26:0]   _zz_3053;
  wire       [35:0]   _zz_3054;
  wire       [17:0]   _zz_3055;
  wire       [17:0]   _zz_3056;
  wire       [35:0]   _zz_3057;
  wire       [35:0]   _zz_3058;
  wire       [17:0]   _zz_3059;
  wire       [35:0]   _zz_3060;
  wire       [35:0]   _zz_3061;
  wire       [35:0]   _zz_3062;
  wire       [17:0]   _zz_3063;
  wire       [35:0]   _zz_3064;
  wire       [35:0]   _zz_3065;
  wire       [35:0]   _zz_3066;
  wire       [35:0]   _zz_3067;
  wire       [35:0]   _zz_3068;
  wire       [35:0]   _zz_3069;
  wire       [26:0]   _zz_3070;
  wire       [35:0]   _zz_3071;
  wire       [17:0]   _zz_3072;
  wire       [35:0]   _zz_3073;
  wire       [35:0]   _zz_3074;
  wire       [35:0]   _zz_3075;
  wire       [35:0]   _zz_3076;
  wire       [35:0]   _zz_3077;
  wire       [26:0]   _zz_3078;
  wire       [35:0]   _zz_3079;
  wire       [17:0]   _zz_3080;
  wire       [35:0]   _zz_3081;
  wire       [35:0]   _zz_3082;
  wire       [35:0]   _zz_3083;
  wire       [35:0]   _zz_3084;
  wire       [35:0]   _zz_3085;
  wire       [26:0]   _zz_3086;
  wire       [35:0]   _zz_3087;
  wire       [17:0]   _zz_3088;
  wire       [35:0]   _zz_3089;
  wire       [35:0]   _zz_3090;
  wire       [35:0]   _zz_3091;
  wire       [35:0]   _zz_3092;
  wire       [35:0]   _zz_3093;
  wire       [26:0]   _zz_3094;
  wire       [35:0]   _zz_3095;
  wire       [17:0]   _zz_3096;
  wire       [17:0]   _zz_3097;
  wire       [35:0]   _zz_3098;
  wire       [35:0]   _zz_3099;
  wire       [17:0]   _zz_3100;
  wire       [35:0]   _zz_3101;
  wire       [35:0]   _zz_3102;
  wire       [35:0]   _zz_3103;
  wire       [17:0]   _zz_3104;
  wire       [35:0]   _zz_3105;
  wire       [35:0]   _zz_3106;
  wire       [35:0]   _zz_3107;
  wire       [35:0]   _zz_3108;
  wire       [35:0]   _zz_3109;
  wire       [35:0]   _zz_3110;
  wire       [26:0]   _zz_3111;
  wire       [35:0]   _zz_3112;
  wire       [17:0]   _zz_3113;
  wire       [35:0]   _zz_3114;
  wire       [35:0]   _zz_3115;
  wire       [35:0]   _zz_3116;
  wire       [35:0]   _zz_3117;
  wire       [35:0]   _zz_3118;
  wire       [26:0]   _zz_3119;
  wire       [35:0]   _zz_3120;
  wire       [17:0]   _zz_3121;
  wire       [35:0]   _zz_3122;
  wire       [35:0]   _zz_3123;
  wire       [35:0]   _zz_3124;
  wire       [35:0]   _zz_3125;
  wire       [35:0]   _zz_3126;
  wire       [26:0]   _zz_3127;
  wire       [35:0]   _zz_3128;
  wire       [17:0]   _zz_3129;
  wire       [35:0]   _zz_3130;
  wire       [35:0]   _zz_3131;
  wire       [35:0]   _zz_3132;
  wire       [35:0]   _zz_3133;
  wire       [35:0]   _zz_3134;
  wire       [26:0]   _zz_3135;
  wire       [35:0]   _zz_3136;
  wire       [17:0]   _zz_3137;
  wire       [17:0]   _zz_3138;
  wire       [35:0]   _zz_3139;
  wire       [35:0]   _zz_3140;
  wire       [17:0]   _zz_3141;
  wire       [35:0]   _zz_3142;
  wire       [35:0]   _zz_3143;
  wire       [35:0]   _zz_3144;
  wire       [17:0]   _zz_3145;
  wire       [35:0]   _zz_3146;
  wire       [35:0]   _zz_3147;
  wire       [35:0]   _zz_3148;
  wire       [35:0]   _zz_3149;
  wire       [35:0]   _zz_3150;
  wire       [35:0]   _zz_3151;
  wire       [26:0]   _zz_3152;
  wire       [35:0]   _zz_3153;
  wire       [17:0]   _zz_3154;
  wire       [35:0]   _zz_3155;
  wire       [35:0]   _zz_3156;
  wire       [35:0]   _zz_3157;
  wire       [35:0]   _zz_3158;
  wire       [35:0]   _zz_3159;
  wire       [26:0]   _zz_3160;
  wire       [35:0]   _zz_3161;
  wire       [17:0]   _zz_3162;
  wire       [35:0]   _zz_3163;
  wire       [35:0]   _zz_3164;
  wire       [35:0]   _zz_3165;
  wire       [35:0]   _zz_3166;
  wire       [35:0]   _zz_3167;
  wire       [26:0]   _zz_3168;
  wire       [35:0]   _zz_3169;
  wire       [17:0]   _zz_3170;
  wire       [35:0]   _zz_3171;
  wire       [35:0]   _zz_3172;
  wire       [35:0]   _zz_3173;
  wire       [35:0]   _zz_3174;
  wire       [35:0]   _zz_3175;
  wire       [26:0]   _zz_3176;
  wire       [35:0]   _zz_3177;
  wire       [17:0]   _zz_3178;
  wire       [17:0]   _zz_3179;
  wire       [35:0]   _zz_3180;
  wire       [35:0]   _zz_3181;
  wire       [17:0]   _zz_3182;
  wire       [35:0]   _zz_3183;
  wire       [35:0]   _zz_3184;
  wire       [35:0]   _zz_3185;
  wire       [17:0]   _zz_3186;
  wire       [35:0]   _zz_3187;
  wire       [35:0]   _zz_3188;
  wire       [35:0]   _zz_3189;
  wire       [35:0]   _zz_3190;
  wire       [35:0]   _zz_3191;
  wire       [35:0]   _zz_3192;
  wire       [26:0]   _zz_3193;
  wire       [35:0]   _zz_3194;
  wire       [17:0]   _zz_3195;
  wire       [35:0]   _zz_3196;
  wire       [35:0]   _zz_3197;
  wire       [35:0]   _zz_3198;
  wire       [35:0]   _zz_3199;
  wire       [35:0]   _zz_3200;
  wire       [26:0]   _zz_3201;
  wire       [35:0]   _zz_3202;
  wire       [17:0]   _zz_3203;
  wire       [35:0]   _zz_3204;
  wire       [35:0]   _zz_3205;
  wire       [35:0]   _zz_3206;
  wire       [35:0]   _zz_3207;
  wire       [35:0]   _zz_3208;
  wire       [26:0]   _zz_3209;
  wire       [35:0]   _zz_3210;
  wire       [17:0]   _zz_3211;
  wire       [35:0]   _zz_3212;
  wire       [35:0]   _zz_3213;
  wire       [35:0]   _zz_3214;
  wire       [35:0]   _zz_3215;
  wire       [35:0]   _zz_3216;
  wire       [26:0]   _zz_3217;
  wire       [35:0]   _zz_3218;
  wire       [17:0]   _zz_3219;
  wire       [17:0]   _zz_3220;
  wire       [35:0]   _zz_3221;
  wire       [35:0]   _zz_3222;
  wire       [17:0]   _zz_3223;
  wire       [35:0]   _zz_3224;
  wire       [35:0]   _zz_3225;
  wire       [35:0]   _zz_3226;
  wire       [17:0]   _zz_3227;
  wire       [35:0]   _zz_3228;
  wire       [35:0]   _zz_3229;
  wire       [35:0]   _zz_3230;
  wire       [35:0]   _zz_3231;
  wire       [35:0]   _zz_3232;
  wire       [35:0]   _zz_3233;
  wire       [26:0]   _zz_3234;
  wire       [35:0]   _zz_3235;
  wire       [17:0]   _zz_3236;
  wire       [35:0]   _zz_3237;
  wire       [35:0]   _zz_3238;
  wire       [35:0]   _zz_3239;
  wire       [35:0]   _zz_3240;
  wire       [35:0]   _zz_3241;
  wire       [26:0]   _zz_3242;
  wire       [35:0]   _zz_3243;
  wire       [17:0]   _zz_3244;
  wire       [35:0]   _zz_3245;
  wire       [35:0]   _zz_3246;
  wire       [35:0]   _zz_3247;
  wire       [35:0]   _zz_3248;
  wire       [35:0]   _zz_3249;
  wire       [26:0]   _zz_3250;
  wire       [35:0]   _zz_3251;
  wire       [17:0]   _zz_3252;
  wire       [35:0]   _zz_3253;
  wire       [35:0]   _zz_3254;
  wire       [35:0]   _zz_3255;
  wire       [35:0]   _zz_3256;
  wire       [35:0]   _zz_3257;
  wire       [26:0]   _zz_3258;
  wire       [35:0]   _zz_3259;
  wire       [17:0]   _zz_3260;
  wire       [17:0]   _zz_3261;
  wire       [35:0]   _zz_3262;
  wire       [35:0]   _zz_3263;
  wire       [17:0]   _zz_3264;
  wire       [35:0]   _zz_3265;
  wire       [35:0]   _zz_3266;
  wire       [35:0]   _zz_3267;
  wire       [17:0]   _zz_3268;
  wire       [35:0]   _zz_3269;
  wire       [35:0]   _zz_3270;
  wire       [35:0]   _zz_3271;
  wire       [35:0]   _zz_3272;
  wire       [35:0]   _zz_3273;
  wire       [35:0]   _zz_3274;
  wire       [26:0]   _zz_3275;
  wire       [35:0]   _zz_3276;
  wire       [17:0]   _zz_3277;
  wire       [35:0]   _zz_3278;
  wire       [35:0]   _zz_3279;
  wire       [35:0]   _zz_3280;
  wire       [35:0]   _zz_3281;
  wire       [35:0]   _zz_3282;
  wire       [26:0]   _zz_3283;
  wire       [35:0]   _zz_3284;
  wire       [17:0]   _zz_3285;
  wire       [35:0]   _zz_3286;
  wire       [35:0]   _zz_3287;
  wire       [35:0]   _zz_3288;
  wire       [35:0]   _zz_3289;
  wire       [35:0]   _zz_3290;
  wire       [26:0]   _zz_3291;
  wire       [35:0]   _zz_3292;
  wire       [17:0]   _zz_3293;
  wire       [35:0]   _zz_3294;
  wire       [35:0]   _zz_3295;
  wire       [35:0]   _zz_3296;
  wire       [35:0]   _zz_3297;
  wire       [35:0]   _zz_3298;
  wire       [26:0]   _zz_3299;
  wire       [35:0]   _zz_3300;
  wire       [17:0]   _zz_3301;
  wire       [17:0]   _zz_3302;
  wire       [35:0]   _zz_3303;
  wire       [35:0]   _zz_3304;
  wire       [17:0]   _zz_3305;
  wire       [35:0]   _zz_3306;
  wire       [35:0]   _zz_3307;
  wire       [35:0]   _zz_3308;
  wire       [17:0]   _zz_3309;
  wire       [35:0]   _zz_3310;
  wire       [35:0]   _zz_3311;
  wire       [35:0]   _zz_3312;
  wire       [35:0]   _zz_3313;
  wire       [35:0]   _zz_3314;
  wire       [35:0]   _zz_3315;
  wire       [26:0]   _zz_3316;
  wire       [35:0]   _zz_3317;
  wire       [17:0]   _zz_3318;
  wire       [35:0]   _zz_3319;
  wire       [35:0]   _zz_3320;
  wire       [35:0]   _zz_3321;
  wire       [35:0]   _zz_3322;
  wire       [35:0]   _zz_3323;
  wire       [26:0]   _zz_3324;
  wire       [35:0]   _zz_3325;
  wire       [17:0]   _zz_3326;
  wire       [35:0]   _zz_3327;
  wire       [35:0]   _zz_3328;
  wire       [35:0]   _zz_3329;
  wire       [35:0]   _zz_3330;
  wire       [35:0]   _zz_3331;
  wire       [26:0]   _zz_3332;
  wire       [35:0]   _zz_3333;
  wire       [17:0]   _zz_3334;
  wire       [35:0]   _zz_3335;
  wire       [35:0]   _zz_3336;
  wire       [35:0]   _zz_3337;
  wire       [35:0]   _zz_3338;
  wire       [35:0]   _zz_3339;
  wire       [26:0]   _zz_3340;
  wire       [35:0]   _zz_3341;
  wire       [17:0]   _zz_3342;
  wire       [17:0]   _zz_3343;
  wire       [35:0]   _zz_3344;
  wire       [35:0]   _zz_3345;
  wire       [17:0]   _zz_3346;
  wire       [35:0]   _zz_3347;
  wire       [35:0]   _zz_3348;
  wire       [35:0]   _zz_3349;
  wire       [17:0]   _zz_3350;
  wire       [35:0]   _zz_3351;
  wire       [35:0]   _zz_3352;
  wire       [35:0]   _zz_3353;
  wire       [35:0]   _zz_3354;
  wire       [35:0]   _zz_3355;
  wire       [35:0]   _zz_3356;
  wire       [26:0]   _zz_3357;
  wire       [35:0]   _zz_3358;
  wire       [17:0]   _zz_3359;
  wire       [35:0]   _zz_3360;
  wire       [35:0]   _zz_3361;
  wire       [35:0]   _zz_3362;
  wire       [35:0]   _zz_3363;
  wire       [35:0]   _zz_3364;
  wire       [26:0]   _zz_3365;
  wire       [35:0]   _zz_3366;
  wire       [17:0]   _zz_3367;
  wire       [35:0]   _zz_3368;
  wire       [35:0]   _zz_3369;
  wire       [35:0]   _zz_3370;
  wire       [35:0]   _zz_3371;
  wire       [35:0]   _zz_3372;
  wire       [26:0]   _zz_3373;
  wire       [35:0]   _zz_3374;
  wire       [17:0]   _zz_3375;
  wire       [35:0]   _zz_3376;
  wire       [35:0]   _zz_3377;
  wire       [35:0]   _zz_3378;
  wire       [35:0]   _zz_3379;
  wire       [35:0]   _zz_3380;
  wire       [26:0]   _zz_3381;
  wire       [35:0]   _zz_3382;
  wire       [17:0]   _zz_3383;
  wire       [17:0]   _zz_3384;
  wire       [35:0]   _zz_3385;
  wire       [35:0]   _zz_3386;
  wire       [17:0]   _zz_3387;
  wire       [35:0]   _zz_3388;
  wire       [35:0]   _zz_3389;
  wire       [35:0]   _zz_3390;
  wire       [17:0]   _zz_3391;
  wire       [35:0]   _zz_3392;
  wire       [35:0]   _zz_3393;
  wire       [35:0]   _zz_3394;
  wire       [35:0]   _zz_3395;
  wire       [35:0]   _zz_3396;
  wire       [35:0]   _zz_3397;
  wire       [26:0]   _zz_3398;
  wire       [35:0]   _zz_3399;
  wire       [17:0]   _zz_3400;
  wire       [35:0]   _zz_3401;
  wire       [35:0]   _zz_3402;
  wire       [35:0]   _zz_3403;
  wire       [35:0]   _zz_3404;
  wire       [35:0]   _zz_3405;
  wire       [26:0]   _zz_3406;
  wire       [35:0]   _zz_3407;
  wire       [17:0]   _zz_3408;
  wire       [35:0]   _zz_3409;
  wire       [35:0]   _zz_3410;
  wire       [35:0]   _zz_3411;
  wire       [35:0]   _zz_3412;
  wire       [35:0]   _zz_3413;
  wire       [26:0]   _zz_3414;
  wire       [35:0]   _zz_3415;
  wire       [17:0]   _zz_3416;
  wire       [35:0]   _zz_3417;
  wire       [35:0]   _zz_3418;
  wire       [35:0]   _zz_3419;
  wire       [35:0]   _zz_3420;
  wire       [35:0]   _zz_3421;
  wire       [26:0]   _zz_3422;
  wire       [35:0]   _zz_3423;
  wire       [17:0]   _zz_3424;
  wire       [17:0]   _zz_3425;
  wire       [35:0]   _zz_3426;
  wire       [35:0]   _zz_3427;
  wire       [17:0]   _zz_3428;
  wire       [35:0]   _zz_3429;
  wire       [35:0]   _zz_3430;
  wire       [35:0]   _zz_3431;
  wire       [17:0]   _zz_3432;
  wire       [35:0]   _zz_3433;
  wire       [35:0]   _zz_3434;
  wire       [35:0]   _zz_3435;
  wire       [35:0]   _zz_3436;
  wire       [35:0]   _zz_3437;
  wire       [35:0]   _zz_3438;
  wire       [26:0]   _zz_3439;
  wire       [35:0]   _zz_3440;
  wire       [17:0]   _zz_3441;
  wire       [35:0]   _zz_3442;
  wire       [35:0]   _zz_3443;
  wire       [35:0]   _zz_3444;
  wire       [35:0]   _zz_3445;
  wire       [35:0]   _zz_3446;
  wire       [26:0]   _zz_3447;
  wire       [35:0]   _zz_3448;
  wire       [17:0]   _zz_3449;
  wire       [35:0]   _zz_3450;
  wire       [35:0]   _zz_3451;
  wire       [35:0]   _zz_3452;
  wire       [35:0]   _zz_3453;
  wire       [35:0]   _zz_3454;
  wire       [26:0]   _zz_3455;
  wire       [35:0]   _zz_3456;
  wire       [17:0]   _zz_3457;
  wire       [35:0]   _zz_3458;
  wire       [35:0]   _zz_3459;
  wire       [35:0]   _zz_3460;
  wire       [35:0]   _zz_3461;
  wire       [35:0]   _zz_3462;
  wire       [26:0]   _zz_3463;
  wire       [35:0]   _zz_3464;
  wire       [17:0]   _zz_3465;
  wire       [17:0]   _zz_3466;
  wire       [35:0]   _zz_3467;
  wire       [35:0]   _zz_3468;
  wire       [17:0]   _zz_3469;
  wire       [35:0]   _zz_3470;
  wire       [35:0]   _zz_3471;
  wire       [35:0]   _zz_3472;
  wire       [17:0]   _zz_3473;
  wire       [35:0]   _zz_3474;
  wire       [35:0]   _zz_3475;
  wire       [35:0]   _zz_3476;
  wire       [35:0]   _zz_3477;
  wire       [35:0]   _zz_3478;
  wire       [35:0]   _zz_3479;
  wire       [26:0]   _zz_3480;
  wire       [35:0]   _zz_3481;
  wire       [17:0]   _zz_3482;
  wire       [35:0]   _zz_3483;
  wire       [35:0]   _zz_3484;
  wire       [35:0]   _zz_3485;
  wire       [35:0]   _zz_3486;
  wire       [35:0]   _zz_3487;
  wire       [26:0]   _zz_3488;
  wire       [35:0]   _zz_3489;
  wire       [17:0]   _zz_3490;
  wire       [35:0]   _zz_3491;
  wire       [35:0]   _zz_3492;
  wire       [35:0]   _zz_3493;
  wire       [35:0]   _zz_3494;
  wire       [35:0]   _zz_3495;
  wire       [26:0]   _zz_3496;
  wire       [35:0]   _zz_3497;
  wire       [17:0]   _zz_3498;
  wire       [35:0]   _zz_3499;
  wire       [35:0]   _zz_3500;
  wire       [35:0]   _zz_3501;
  wire       [35:0]   _zz_3502;
  wire       [35:0]   _zz_3503;
  wire       [26:0]   _zz_3504;
  wire       [35:0]   _zz_3505;
  wire       [17:0]   _zz_3506;
  wire       [17:0]   _zz_3507;
  wire       [35:0]   _zz_3508;
  wire       [35:0]   _zz_3509;
  wire       [17:0]   _zz_3510;
  wire       [35:0]   _zz_3511;
  wire       [35:0]   _zz_3512;
  wire       [35:0]   _zz_3513;
  wire       [17:0]   _zz_3514;
  wire       [35:0]   _zz_3515;
  wire       [35:0]   _zz_3516;
  wire       [35:0]   _zz_3517;
  wire       [35:0]   _zz_3518;
  wire       [35:0]   _zz_3519;
  wire       [35:0]   _zz_3520;
  wire       [26:0]   _zz_3521;
  wire       [35:0]   _zz_3522;
  wire       [17:0]   _zz_3523;
  wire       [35:0]   _zz_3524;
  wire       [35:0]   _zz_3525;
  wire       [35:0]   _zz_3526;
  wire       [35:0]   _zz_3527;
  wire       [35:0]   _zz_3528;
  wire       [26:0]   _zz_3529;
  wire       [35:0]   _zz_3530;
  wire       [17:0]   _zz_3531;
  wire       [35:0]   _zz_3532;
  wire       [35:0]   _zz_3533;
  wire       [35:0]   _zz_3534;
  wire       [35:0]   _zz_3535;
  wire       [35:0]   _zz_3536;
  wire       [26:0]   _zz_3537;
  wire       [35:0]   _zz_3538;
  wire       [17:0]   _zz_3539;
  wire       [35:0]   _zz_3540;
  wire       [35:0]   _zz_3541;
  wire       [35:0]   _zz_3542;
  wire       [35:0]   _zz_3543;
  wire       [35:0]   _zz_3544;
  wire       [26:0]   _zz_3545;
  wire       [35:0]   _zz_3546;
  wire       [17:0]   _zz_3547;
  wire       [17:0]   _zz_3548;
  wire       [35:0]   _zz_3549;
  wire       [35:0]   _zz_3550;
  wire       [17:0]   _zz_3551;
  wire       [35:0]   _zz_3552;
  wire       [35:0]   _zz_3553;
  wire       [35:0]   _zz_3554;
  wire       [17:0]   _zz_3555;
  wire       [35:0]   _zz_3556;
  wire       [35:0]   _zz_3557;
  wire       [35:0]   _zz_3558;
  wire       [35:0]   _zz_3559;
  wire       [35:0]   _zz_3560;
  wire       [35:0]   _zz_3561;
  wire       [26:0]   _zz_3562;
  wire       [35:0]   _zz_3563;
  wire       [17:0]   _zz_3564;
  wire       [35:0]   _zz_3565;
  wire       [35:0]   _zz_3566;
  wire       [35:0]   _zz_3567;
  wire       [35:0]   _zz_3568;
  wire       [35:0]   _zz_3569;
  wire       [26:0]   _zz_3570;
  wire       [35:0]   _zz_3571;
  wire       [17:0]   _zz_3572;
  wire       [35:0]   _zz_3573;
  wire       [35:0]   _zz_3574;
  wire       [35:0]   _zz_3575;
  wire       [35:0]   _zz_3576;
  wire       [35:0]   _zz_3577;
  wire       [26:0]   _zz_3578;
  wire       [35:0]   _zz_3579;
  wire       [17:0]   _zz_3580;
  wire       [35:0]   _zz_3581;
  wire       [35:0]   _zz_3582;
  wire       [35:0]   _zz_3583;
  wire       [35:0]   _zz_3584;
  wire       [35:0]   _zz_3585;
  wire       [26:0]   _zz_3586;
  wire       [35:0]   _zz_3587;
  wire       [17:0]   _zz_3588;
  wire       [17:0]   _zz_3589;
  wire       [35:0]   _zz_3590;
  wire       [35:0]   _zz_3591;
  wire       [17:0]   _zz_3592;
  wire       [35:0]   _zz_3593;
  wire       [35:0]   _zz_3594;
  wire       [35:0]   _zz_3595;
  wire       [17:0]   _zz_3596;
  wire       [35:0]   _zz_3597;
  wire       [35:0]   _zz_3598;
  wire       [35:0]   _zz_3599;
  wire       [35:0]   _zz_3600;
  wire       [35:0]   _zz_3601;
  wire       [35:0]   _zz_3602;
  wire       [26:0]   _zz_3603;
  wire       [35:0]   _zz_3604;
  wire       [17:0]   _zz_3605;
  wire       [35:0]   _zz_3606;
  wire       [35:0]   _zz_3607;
  wire       [35:0]   _zz_3608;
  wire       [35:0]   _zz_3609;
  wire       [35:0]   _zz_3610;
  wire       [26:0]   _zz_3611;
  wire       [35:0]   _zz_3612;
  wire       [17:0]   _zz_3613;
  wire       [35:0]   _zz_3614;
  wire       [35:0]   _zz_3615;
  wire       [35:0]   _zz_3616;
  wire       [35:0]   _zz_3617;
  wire       [35:0]   _zz_3618;
  wire       [26:0]   _zz_3619;
  wire       [35:0]   _zz_3620;
  wire       [17:0]   _zz_3621;
  wire       [35:0]   _zz_3622;
  wire       [35:0]   _zz_3623;
  wire       [35:0]   _zz_3624;
  wire       [35:0]   _zz_3625;
  wire       [35:0]   _zz_3626;
  wire       [26:0]   _zz_3627;
  wire       [35:0]   _zz_3628;
  wire       [17:0]   _zz_3629;
  wire       [17:0]   _zz_3630;
  wire       [35:0]   _zz_3631;
  wire       [35:0]   _zz_3632;
  wire       [17:0]   _zz_3633;
  wire       [35:0]   _zz_3634;
  wire       [35:0]   _zz_3635;
  wire       [35:0]   _zz_3636;
  wire       [17:0]   _zz_3637;
  wire       [35:0]   _zz_3638;
  wire       [35:0]   _zz_3639;
  wire       [35:0]   _zz_3640;
  wire       [35:0]   _zz_3641;
  wire       [35:0]   _zz_3642;
  wire       [35:0]   _zz_3643;
  wire       [26:0]   _zz_3644;
  wire       [35:0]   _zz_3645;
  wire       [17:0]   _zz_3646;
  wire       [35:0]   _zz_3647;
  wire       [35:0]   _zz_3648;
  wire       [35:0]   _zz_3649;
  wire       [35:0]   _zz_3650;
  wire       [35:0]   _zz_3651;
  wire       [26:0]   _zz_3652;
  wire       [35:0]   _zz_3653;
  wire       [17:0]   _zz_3654;
  wire       [35:0]   _zz_3655;
  wire       [35:0]   _zz_3656;
  wire       [35:0]   _zz_3657;
  wire       [35:0]   _zz_3658;
  wire       [35:0]   _zz_3659;
  wire       [26:0]   _zz_3660;
  wire       [35:0]   _zz_3661;
  wire       [17:0]   _zz_3662;
  wire       [35:0]   _zz_3663;
  wire       [35:0]   _zz_3664;
  wire       [35:0]   _zz_3665;
  wire       [35:0]   _zz_3666;
  wire       [35:0]   _zz_3667;
  wire       [26:0]   _zz_3668;
  wire       [35:0]   _zz_3669;
  wire       [17:0]   _zz_3670;
  wire       [17:0]   _zz_3671;
  wire       [35:0]   _zz_3672;
  wire       [35:0]   _zz_3673;
  wire       [17:0]   _zz_3674;
  wire       [35:0]   _zz_3675;
  wire       [35:0]   _zz_3676;
  wire       [35:0]   _zz_3677;
  wire       [17:0]   _zz_3678;
  wire       [35:0]   _zz_3679;
  wire       [35:0]   _zz_3680;
  wire       [35:0]   _zz_3681;
  wire       [35:0]   _zz_3682;
  wire       [35:0]   _zz_3683;
  wire       [35:0]   _zz_3684;
  wire       [26:0]   _zz_3685;
  wire       [35:0]   _zz_3686;
  wire       [17:0]   _zz_3687;
  wire       [35:0]   _zz_3688;
  wire       [35:0]   _zz_3689;
  wire       [35:0]   _zz_3690;
  wire       [35:0]   _zz_3691;
  wire       [35:0]   _zz_3692;
  wire       [26:0]   _zz_3693;
  wire       [35:0]   _zz_3694;
  wire       [17:0]   _zz_3695;
  wire       [35:0]   _zz_3696;
  wire       [35:0]   _zz_3697;
  wire       [35:0]   _zz_3698;
  wire       [35:0]   _zz_3699;
  wire       [35:0]   _zz_3700;
  wire       [26:0]   _zz_3701;
  wire       [35:0]   _zz_3702;
  wire       [17:0]   _zz_3703;
  wire       [35:0]   _zz_3704;
  wire       [35:0]   _zz_3705;
  wire       [35:0]   _zz_3706;
  wire       [35:0]   _zz_3707;
  wire       [35:0]   _zz_3708;
  wire       [26:0]   _zz_3709;
  wire       [35:0]   _zz_3710;
  wire       [17:0]   _zz_3711;
  wire       [17:0]   _zz_3712;
  wire       [35:0]   _zz_3713;
  wire       [35:0]   _zz_3714;
  wire       [17:0]   _zz_3715;
  wire       [35:0]   _zz_3716;
  wire       [35:0]   _zz_3717;
  wire       [35:0]   _zz_3718;
  wire       [17:0]   _zz_3719;
  wire       [35:0]   _zz_3720;
  wire       [35:0]   _zz_3721;
  wire       [35:0]   _zz_3722;
  wire       [35:0]   _zz_3723;
  wire       [35:0]   _zz_3724;
  wire       [35:0]   _zz_3725;
  wire       [26:0]   _zz_3726;
  wire       [35:0]   _zz_3727;
  wire       [17:0]   _zz_3728;
  wire       [35:0]   _zz_3729;
  wire       [35:0]   _zz_3730;
  wire       [35:0]   _zz_3731;
  wire       [35:0]   _zz_3732;
  wire       [35:0]   _zz_3733;
  wire       [26:0]   _zz_3734;
  wire       [35:0]   _zz_3735;
  wire       [17:0]   _zz_3736;
  wire       [35:0]   _zz_3737;
  wire       [35:0]   _zz_3738;
  wire       [35:0]   _zz_3739;
  wire       [35:0]   _zz_3740;
  wire       [35:0]   _zz_3741;
  wire       [26:0]   _zz_3742;
  wire       [35:0]   _zz_3743;
  wire       [17:0]   _zz_3744;
  wire       [35:0]   _zz_3745;
  wire       [35:0]   _zz_3746;
  wire       [35:0]   _zz_3747;
  wire       [35:0]   _zz_3748;
  wire       [35:0]   _zz_3749;
  wire       [26:0]   _zz_3750;
  wire       [35:0]   _zz_3751;
  wire       [17:0]   _zz_3752;
  wire       [17:0]   _zz_3753;
  wire       [35:0]   _zz_3754;
  wire       [35:0]   _zz_3755;
  wire       [17:0]   _zz_3756;
  wire       [35:0]   _zz_3757;
  wire       [35:0]   _zz_3758;
  wire       [35:0]   _zz_3759;
  wire       [17:0]   _zz_3760;
  wire       [35:0]   _zz_3761;
  wire       [35:0]   _zz_3762;
  wire       [35:0]   _zz_3763;
  wire       [35:0]   _zz_3764;
  wire       [35:0]   _zz_3765;
  wire       [35:0]   _zz_3766;
  wire       [26:0]   _zz_3767;
  wire       [35:0]   _zz_3768;
  wire       [17:0]   _zz_3769;
  wire       [35:0]   _zz_3770;
  wire       [35:0]   _zz_3771;
  wire       [35:0]   _zz_3772;
  wire       [35:0]   _zz_3773;
  wire       [35:0]   _zz_3774;
  wire       [26:0]   _zz_3775;
  wire       [35:0]   _zz_3776;
  wire       [17:0]   _zz_3777;
  wire       [35:0]   _zz_3778;
  wire       [35:0]   _zz_3779;
  wire       [35:0]   _zz_3780;
  wire       [35:0]   _zz_3781;
  wire       [35:0]   _zz_3782;
  wire       [26:0]   _zz_3783;
  wire       [35:0]   _zz_3784;
  wire       [17:0]   _zz_3785;
  wire       [35:0]   _zz_3786;
  wire       [35:0]   _zz_3787;
  wire       [35:0]   _zz_3788;
  wire       [35:0]   _zz_3789;
  wire       [35:0]   _zz_3790;
  wire       [26:0]   _zz_3791;
  wire       [35:0]   _zz_3792;
  wire       [17:0]   _zz_3793;
  wire       [17:0]   _zz_3794;
  wire       [35:0]   _zz_3795;
  wire       [35:0]   _zz_3796;
  wire       [17:0]   _zz_3797;
  wire       [35:0]   _zz_3798;
  wire       [35:0]   _zz_3799;
  wire       [35:0]   _zz_3800;
  wire       [17:0]   _zz_3801;
  wire       [35:0]   _zz_3802;
  wire       [35:0]   _zz_3803;
  wire       [35:0]   _zz_3804;
  wire       [35:0]   _zz_3805;
  wire       [35:0]   _zz_3806;
  wire       [35:0]   _zz_3807;
  wire       [26:0]   _zz_3808;
  wire       [35:0]   _zz_3809;
  wire       [17:0]   _zz_3810;
  wire       [35:0]   _zz_3811;
  wire       [35:0]   _zz_3812;
  wire       [35:0]   _zz_3813;
  wire       [35:0]   _zz_3814;
  wire       [35:0]   _zz_3815;
  wire       [26:0]   _zz_3816;
  wire       [35:0]   _zz_3817;
  wire       [17:0]   _zz_3818;
  wire       [35:0]   _zz_3819;
  wire       [35:0]   _zz_3820;
  wire       [35:0]   _zz_3821;
  wire       [35:0]   _zz_3822;
  wire       [35:0]   _zz_3823;
  wire       [26:0]   _zz_3824;
  wire       [35:0]   _zz_3825;
  wire       [17:0]   _zz_3826;
  wire       [35:0]   _zz_3827;
  wire       [35:0]   _zz_3828;
  wire       [35:0]   _zz_3829;
  wire       [35:0]   _zz_3830;
  wire       [35:0]   _zz_3831;
  wire       [26:0]   _zz_3832;
  wire       [35:0]   _zz_3833;
  wire       [17:0]   _zz_3834;
  wire       [17:0]   _zz_3835;
  wire       [35:0]   _zz_3836;
  wire       [35:0]   _zz_3837;
  wire       [17:0]   _zz_3838;
  wire       [35:0]   _zz_3839;
  wire       [35:0]   _zz_3840;
  wire       [35:0]   _zz_3841;
  wire       [17:0]   _zz_3842;
  wire       [35:0]   _zz_3843;
  wire       [35:0]   _zz_3844;
  wire       [35:0]   _zz_3845;
  wire       [35:0]   _zz_3846;
  wire       [35:0]   _zz_3847;
  wire       [35:0]   _zz_3848;
  wire       [26:0]   _zz_3849;
  wire       [35:0]   _zz_3850;
  wire       [17:0]   _zz_3851;
  wire       [35:0]   _zz_3852;
  wire       [35:0]   _zz_3853;
  wire       [35:0]   _zz_3854;
  wire       [35:0]   _zz_3855;
  wire       [35:0]   _zz_3856;
  wire       [26:0]   _zz_3857;
  wire       [35:0]   _zz_3858;
  wire       [17:0]   _zz_3859;
  wire       [35:0]   _zz_3860;
  wire       [35:0]   _zz_3861;
  wire       [35:0]   _zz_3862;
  wire       [35:0]   _zz_3863;
  wire       [35:0]   _zz_3864;
  wire       [26:0]   _zz_3865;
  wire       [35:0]   _zz_3866;
  wire       [17:0]   _zz_3867;
  wire       [35:0]   _zz_3868;
  wire       [35:0]   _zz_3869;
  wire       [35:0]   _zz_3870;
  wire       [35:0]   _zz_3871;
  wire       [35:0]   _zz_3872;
  wire       [26:0]   _zz_3873;
  wire       [35:0]   _zz_3874;
  wire       [17:0]   _zz_3875;
  wire       [17:0]   _zz_3876;
  wire       [35:0]   _zz_3877;
  wire       [35:0]   _zz_3878;
  wire       [17:0]   _zz_3879;
  wire       [35:0]   _zz_3880;
  wire       [35:0]   _zz_3881;
  wire       [35:0]   _zz_3882;
  wire       [17:0]   _zz_3883;
  wire       [35:0]   _zz_3884;
  wire       [35:0]   _zz_3885;
  wire       [35:0]   _zz_3886;
  wire       [35:0]   _zz_3887;
  wire       [35:0]   _zz_3888;
  wire       [35:0]   _zz_3889;
  wire       [26:0]   _zz_3890;
  wire       [35:0]   _zz_3891;
  wire       [17:0]   _zz_3892;
  wire       [35:0]   _zz_3893;
  wire       [35:0]   _zz_3894;
  wire       [35:0]   _zz_3895;
  wire       [35:0]   _zz_3896;
  wire       [35:0]   _zz_3897;
  wire       [26:0]   _zz_3898;
  wire       [35:0]   _zz_3899;
  wire       [17:0]   _zz_3900;
  wire       [35:0]   _zz_3901;
  wire       [35:0]   _zz_3902;
  wire       [35:0]   _zz_3903;
  wire       [35:0]   _zz_3904;
  wire       [35:0]   _zz_3905;
  wire       [26:0]   _zz_3906;
  wire       [35:0]   _zz_3907;
  wire       [17:0]   _zz_3908;
  wire       [35:0]   _zz_3909;
  wire       [35:0]   _zz_3910;
  wire       [35:0]   _zz_3911;
  wire       [35:0]   _zz_3912;
  wire       [35:0]   _zz_3913;
  wire       [26:0]   _zz_3914;
  wire       [35:0]   _zz_3915;
  wire       [17:0]   _zz_3916;
  wire       [17:0]   _zz_3917;
  wire       [35:0]   _zz_3918;
  wire       [35:0]   _zz_3919;
  wire       [17:0]   _zz_3920;
  wire       [35:0]   _zz_3921;
  wire       [35:0]   _zz_3922;
  wire       [35:0]   _zz_3923;
  wire       [17:0]   _zz_3924;
  wire       [35:0]   _zz_3925;
  wire       [35:0]   _zz_3926;
  wire       [35:0]   _zz_3927;
  wire       [35:0]   _zz_3928;
  wire       [35:0]   _zz_3929;
  wire       [35:0]   _zz_3930;
  wire       [26:0]   _zz_3931;
  wire       [35:0]   _zz_3932;
  wire       [17:0]   _zz_3933;
  wire       [35:0]   _zz_3934;
  wire       [35:0]   _zz_3935;
  wire       [35:0]   _zz_3936;
  wire       [35:0]   _zz_3937;
  wire       [35:0]   _zz_3938;
  wire       [26:0]   _zz_3939;
  wire       [35:0]   _zz_3940;
  wire       [17:0]   _zz_3941;
  wire       [35:0]   _zz_3942;
  wire       [35:0]   _zz_3943;
  wire       [35:0]   _zz_3944;
  wire       [35:0]   _zz_3945;
  wire       [35:0]   _zz_3946;
  wire       [26:0]   _zz_3947;
  wire       [35:0]   _zz_3948;
  wire       [17:0]   _zz_3949;
  wire       [35:0]   _zz_3950;
  wire       [35:0]   _zz_3951;
  wire       [35:0]   _zz_3952;
  wire       [35:0]   _zz_3953;
  wire       [35:0]   _zz_3954;
  wire       [26:0]   _zz_3955;
  wire       [35:0]   _zz_3956;
  wire       [17:0]   _zz_3957;
  wire       [17:0]   _zz_3958;
  wire       [35:0]   _zz_3959;
  wire       [35:0]   _zz_3960;
  wire       [17:0]   _zz_3961;
  wire       [35:0]   _zz_3962;
  wire       [35:0]   _zz_3963;
  wire       [35:0]   _zz_3964;
  wire       [17:0]   _zz_3965;
  wire       [35:0]   _zz_3966;
  wire       [35:0]   _zz_3967;
  wire       [35:0]   _zz_3968;
  wire       [35:0]   _zz_3969;
  wire       [35:0]   _zz_3970;
  wire       [35:0]   _zz_3971;
  wire       [26:0]   _zz_3972;
  wire       [35:0]   _zz_3973;
  wire       [17:0]   _zz_3974;
  wire       [35:0]   _zz_3975;
  wire       [35:0]   _zz_3976;
  wire       [35:0]   _zz_3977;
  wire       [35:0]   _zz_3978;
  wire       [35:0]   _zz_3979;
  wire       [26:0]   _zz_3980;
  wire       [35:0]   _zz_3981;
  wire       [17:0]   _zz_3982;
  wire       [35:0]   _zz_3983;
  wire       [35:0]   _zz_3984;
  wire       [35:0]   _zz_3985;
  wire       [35:0]   _zz_3986;
  wire       [35:0]   _zz_3987;
  wire       [26:0]   _zz_3988;
  wire       [35:0]   _zz_3989;
  wire       [17:0]   _zz_3990;
  wire       [35:0]   _zz_3991;
  wire       [35:0]   _zz_3992;
  wire       [35:0]   _zz_3993;
  wire       [35:0]   _zz_3994;
  wire       [35:0]   _zz_3995;
  wire       [26:0]   _zz_3996;
  wire       [35:0]   _zz_3997;
  wire       [17:0]   _zz_3998;
  wire       [17:0]   _zz_3999;
  wire       [35:0]   _zz_4000;
  wire       [35:0]   _zz_4001;
  wire       [17:0]   _zz_4002;
  wire       [35:0]   _zz_4003;
  wire       [35:0]   _zz_4004;
  wire       [35:0]   _zz_4005;
  wire       [17:0]   _zz_4006;
  wire       [35:0]   _zz_4007;
  wire       [35:0]   _zz_4008;
  wire       [35:0]   _zz_4009;
  wire       [35:0]   _zz_4010;
  wire       [35:0]   _zz_4011;
  wire       [35:0]   _zz_4012;
  wire       [26:0]   _zz_4013;
  wire       [35:0]   _zz_4014;
  wire       [17:0]   _zz_4015;
  wire       [35:0]   _zz_4016;
  wire       [35:0]   _zz_4017;
  wire       [35:0]   _zz_4018;
  wire       [35:0]   _zz_4019;
  wire       [35:0]   _zz_4020;
  wire       [26:0]   _zz_4021;
  wire       [35:0]   _zz_4022;
  wire       [17:0]   _zz_4023;
  wire       [35:0]   _zz_4024;
  wire       [35:0]   _zz_4025;
  wire       [35:0]   _zz_4026;
  wire       [35:0]   _zz_4027;
  wire       [35:0]   _zz_4028;
  wire       [26:0]   _zz_4029;
  wire       [35:0]   _zz_4030;
  wire       [17:0]   _zz_4031;
  wire       [35:0]   _zz_4032;
  wire       [35:0]   _zz_4033;
  wire       [35:0]   _zz_4034;
  wire       [35:0]   _zz_4035;
  wire       [35:0]   _zz_4036;
  wire       [26:0]   _zz_4037;
  wire       [35:0]   _zz_4038;
  wire       [17:0]   _zz_4039;
  wire       [17:0]   _zz_4040;
  wire       [35:0]   _zz_4041;
  wire       [35:0]   _zz_4042;
  wire       [17:0]   _zz_4043;
  wire       [35:0]   _zz_4044;
  wire       [35:0]   _zz_4045;
  wire       [35:0]   _zz_4046;
  wire       [17:0]   _zz_4047;
  wire       [35:0]   _zz_4048;
  wire       [35:0]   _zz_4049;
  wire       [35:0]   _zz_4050;
  wire       [35:0]   _zz_4051;
  wire       [35:0]   _zz_4052;
  wire       [35:0]   _zz_4053;
  wire       [26:0]   _zz_4054;
  wire       [35:0]   _zz_4055;
  wire       [17:0]   _zz_4056;
  wire       [35:0]   _zz_4057;
  wire       [35:0]   _zz_4058;
  wire       [35:0]   _zz_4059;
  wire       [35:0]   _zz_4060;
  wire       [35:0]   _zz_4061;
  wire       [26:0]   _zz_4062;
  wire       [35:0]   _zz_4063;
  wire       [17:0]   _zz_4064;
  wire       [35:0]   _zz_4065;
  wire       [35:0]   _zz_4066;
  wire       [35:0]   _zz_4067;
  wire       [35:0]   _zz_4068;
  wire       [35:0]   _zz_4069;
  wire       [26:0]   _zz_4070;
  wire       [35:0]   _zz_4071;
  wire       [17:0]   _zz_4072;
  wire       [35:0]   _zz_4073;
  wire       [35:0]   _zz_4074;
  wire       [35:0]   _zz_4075;
  wire       [35:0]   _zz_4076;
  wire       [35:0]   _zz_4077;
  wire       [26:0]   _zz_4078;
  wire       [35:0]   _zz_4079;
  wire       [17:0]   _zz_4080;
  wire       [17:0]   _zz_4081;
  wire       [35:0]   _zz_4082;
  wire       [35:0]   _zz_4083;
  wire       [17:0]   _zz_4084;
  wire       [35:0]   _zz_4085;
  wire       [35:0]   _zz_4086;
  wire       [35:0]   _zz_4087;
  wire       [17:0]   _zz_4088;
  wire       [35:0]   _zz_4089;
  wire       [35:0]   _zz_4090;
  wire       [35:0]   _zz_4091;
  wire       [35:0]   _zz_4092;
  wire       [35:0]   _zz_4093;
  wire       [35:0]   _zz_4094;
  wire       [26:0]   _zz_4095;
  wire       [35:0]   _zz_4096;
  wire       [17:0]   _zz_4097;
  wire       [35:0]   _zz_4098;
  wire       [35:0]   _zz_4099;
  wire       [35:0]   _zz_4100;
  wire       [35:0]   _zz_4101;
  wire       [35:0]   _zz_4102;
  wire       [26:0]   _zz_4103;
  wire       [35:0]   _zz_4104;
  wire       [17:0]   _zz_4105;
  wire       [35:0]   _zz_4106;
  wire       [35:0]   _zz_4107;
  wire       [35:0]   _zz_4108;
  wire       [35:0]   _zz_4109;
  wire       [35:0]   _zz_4110;
  wire       [26:0]   _zz_4111;
  wire       [35:0]   _zz_4112;
  wire       [17:0]   _zz_4113;
  wire       [35:0]   _zz_4114;
  wire       [35:0]   _zz_4115;
  wire       [35:0]   _zz_4116;
  wire       [35:0]   _zz_4117;
  wire       [35:0]   _zz_4118;
  wire       [26:0]   _zz_4119;
  wire       [35:0]   _zz_4120;
  wire       [17:0]   _zz_4121;
  wire       [17:0]   _zz_4122;
  wire       [35:0]   _zz_4123;
  wire       [35:0]   _zz_4124;
  wire       [17:0]   _zz_4125;
  wire       [35:0]   _zz_4126;
  wire       [35:0]   _zz_4127;
  wire       [35:0]   _zz_4128;
  wire       [17:0]   _zz_4129;
  wire       [35:0]   _zz_4130;
  wire       [35:0]   _zz_4131;
  wire       [35:0]   _zz_4132;
  wire       [35:0]   _zz_4133;
  wire       [35:0]   _zz_4134;
  wire       [35:0]   _zz_4135;
  wire       [26:0]   _zz_4136;
  wire       [35:0]   _zz_4137;
  wire       [17:0]   _zz_4138;
  wire       [35:0]   _zz_4139;
  wire       [35:0]   _zz_4140;
  wire       [35:0]   _zz_4141;
  wire       [35:0]   _zz_4142;
  wire       [35:0]   _zz_4143;
  wire       [26:0]   _zz_4144;
  wire       [35:0]   _zz_4145;
  wire       [17:0]   _zz_4146;
  wire       [35:0]   _zz_4147;
  wire       [35:0]   _zz_4148;
  wire       [35:0]   _zz_4149;
  wire       [35:0]   _zz_4150;
  wire       [35:0]   _zz_4151;
  wire       [26:0]   _zz_4152;
  wire       [35:0]   _zz_4153;
  wire       [17:0]   _zz_4154;
  wire       [35:0]   _zz_4155;
  wire       [35:0]   _zz_4156;
  wire       [35:0]   _zz_4157;
  wire       [35:0]   _zz_4158;
  wire       [35:0]   _zz_4159;
  wire       [26:0]   _zz_4160;
  wire       [35:0]   _zz_4161;
  wire       [17:0]   _zz_4162;
  wire       [17:0]   _zz_4163;
  wire       [35:0]   _zz_4164;
  wire       [35:0]   _zz_4165;
  wire       [17:0]   _zz_4166;
  wire       [35:0]   _zz_4167;
  wire       [35:0]   _zz_4168;
  wire       [35:0]   _zz_4169;
  wire       [17:0]   _zz_4170;
  wire       [35:0]   _zz_4171;
  wire       [35:0]   _zz_4172;
  wire       [35:0]   _zz_4173;
  wire       [35:0]   _zz_4174;
  wire       [35:0]   _zz_4175;
  wire       [35:0]   _zz_4176;
  wire       [26:0]   _zz_4177;
  wire       [35:0]   _zz_4178;
  wire       [17:0]   _zz_4179;
  wire       [35:0]   _zz_4180;
  wire       [35:0]   _zz_4181;
  wire       [35:0]   _zz_4182;
  wire       [35:0]   _zz_4183;
  wire       [35:0]   _zz_4184;
  wire       [26:0]   _zz_4185;
  wire       [35:0]   _zz_4186;
  wire       [17:0]   _zz_4187;
  wire       [35:0]   _zz_4188;
  wire       [35:0]   _zz_4189;
  wire       [35:0]   _zz_4190;
  wire       [35:0]   _zz_4191;
  wire       [35:0]   _zz_4192;
  wire       [26:0]   _zz_4193;
  wire       [35:0]   _zz_4194;
  wire       [17:0]   _zz_4195;
  wire       [35:0]   _zz_4196;
  wire       [35:0]   _zz_4197;
  wire       [35:0]   _zz_4198;
  wire       [35:0]   _zz_4199;
  wire       [35:0]   _zz_4200;
  wire       [26:0]   _zz_4201;
  wire       [35:0]   _zz_4202;
  wire       [17:0]   _zz_4203;
  wire       [17:0]   _zz_4204;
  wire       [35:0]   _zz_4205;
  wire       [35:0]   _zz_4206;
  wire       [17:0]   _zz_4207;
  wire       [35:0]   _zz_4208;
  wire       [35:0]   _zz_4209;
  wire       [35:0]   _zz_4210;
  wire       [17:0]   _zz_4211;
  wire       [35:0]   _zz_4212;
  wire       [35:0]   _zz_4213;
  wire       [35:0]   _zz_4214;
  wire       [35:0]   _zz_4215;
  wire       [35:0]   _zz_4216;
  wire       [35:0]   _zz_4217;
  wire       [26:0]   _zz_4218;
  wire       [35:0]   _zz_4219;
  wire       [17:0]   _zz_4220;
  wire       [35:0]   _zz_4221;
  wire       [35:0]   _zz_4222;
  wire       [35:0]   _zz_4223;
  wire       [35:0]   _zz_4224;
  wire       [35:0]   _zz_4225;
  wire       [26:0]   _zz_4226;
  wire       [35:0]   _zz_4227;
  wire       [17:0]   _zz_4228;
  wire       [35:0]   _zz_4229;
  wire       [35:0]   _zz_4230;
  wire       [35:0]   _zz_4231;
  wire       [35:0]   _zz_4232;
  wire       [35:0]   _zz_4233;
  wire       [26:0]   _zz_4234;
  wire       [35:0]   _zz_4235;
  wire       [17:0]   _zz_4236;
  wire       [35:0]   _zz_4237;
  wire       [35:0]   _zz_4238;
  wire       [35:0]   _zz_4239;
  wire       [35:0]   _zz_4240;
  wire       [35:0]   _zz_4241;
  wire       [26:0]   _zz_4242;
  wire       [35:0]   _zz_4243;
  wire       [17:0]   _zz_4244;
  wire       [17:0]   _zz_4245;
  wire       [35:0]   _zz_4246;
  wire       [35:0]   _zz_4247;
  wire       [17:0]   _zz_4248;
  wire       [35:0]   _zz_4249;
  wire       [35:0]   _zz_4250;
  wire       [35:0]   _zz_4251;
  wire       [17:0]   _zz_4252;
  wire       [35:0]   _zz_4253;
  wire       [35:0]   _zz_4254;
  wire       [35:0]   _zz_4255;
  wire       [35:0]   _zz_4256;
  wire       [35:0]   _zz_4257;
  wire       [35:0]   _zz_4258;
  wire       [26:0]   _zz_4259;
  wire       [35:0]   _zz_4260;
  wire       [17:0]   _zz_4261;
  wire       [35:0]   _zz_4262;
  wire       [35:0]   _zz_4263;
  wire       [35:0]   _zz_4264;
  wire       [35:0]   _zz_4265;
  wire       [35:0]   _zz_4266;
  wire       [26:0]   _zz_4267;
  wire       [35:0]   _zz_4268;
  wire       [17:0]   _zz_4269;
  wire       [35:0]   _zz_4270;
  wire       [35:0]   _zz_4271;
  wire       [35:0]   _zz_4272;
  wire       [35:0]   _zz_4273;
  wire       [35:0]   _zz_4274;
  wire       [26:0]   _zz_4275;
  wire       [35:0]   _zz_4276;
  wire       [17:0]   _zz_4277;
  wire       [35:0]   _zz_4278;
  wire       [35:0]   _zz_4279;
  wire       [35:0]   _zz_4280;
  wire       [35:0]   _zz_4281;
  wire       [35:0]   _zz_4282;
  wire       [26:0]   _zz_4283;
  wire       [35:0]   _zz_4284;
  wire       [17:0]   _zz_4285;
  wire       [17:0]   _zz_4286;
  wire       [35:0]   _zz_4287;
  wire       [35:0]   _zz_4288;
  wire       [17:0]   _zz_4289;
  wire       [35:0]   _zz_4290;
  wire       [35:0]   _zz_4291;
  wire       [35:0]   _zz_4292;
  wire       [17:0]   _zz_4293;
  wire       [35:0]   _zz_4294;
  wire       [35:0]   _zz_4295;
  wire       [35:0]   _zz_4296;
  wire       [35:0]   _zz_4297;
  wire       [35:0]   _zz_4298;
  wire       [35:0]   _zz_4299;
  wire       [26:0]   _zz_4300;
  wire       [35:0]   _zz_4301;
  wire       [17:0]   _zz_4302;
  wire       [35:0]   _zz_4303;
  wire       [35:0]   _zz_4304;
  wire       [35:0]   _zz_4305;
  wire       [35:0]   _zz_4306;
  wire       [35:0]   _zz_4307;
  wire       [26:0]   _zz_4308;
  wire       [35:0]   _zz_4309;
  wire       [17:0]   _zz_4310;
  wire       [35:0]   _zz_4311;
  wire       [35:0]   _zz_4312;
  wire       [35:0]   _zz_4313;
  wire       [35:0]   _zz_4314;
  wire       [35:0]   _zz_4315;
  wire       [26:0]   _zz_4316;
  wire       [35:0]   _zz_4317;
  wire       [17:0]   _zz_4318;
  wire       [35:0]   _zz_4319;
  wire       [35:0]   _zz_4320;
  wire       [35:0]   _zz_4321;
  wire       [35:0]   _zz_4322;
  wire       [35:0]   _zz_4323;
  wire       [26:0]   _zz_4324;
  wire       [35:0]   _zz_4325;
  wire       [17:0]   _zz_4326;
  wire       [17:0]   _zz_4327;
  wire       [35:0]   _zz_4328;
  wire       [35:0]   _zz_4329;
  wire       [17:0]   _zz_4330;
  wire       [35:0]   _zz_4331;
  wire       [35:0]   _zz_4332;
  wire       [35:0]   _zz_4333;
  wire       [17:0]   _zz_4334;
  wire       [35:0]   _zz_4335;
  wire       [35:0]   _zz_4336;
  wire       [35:0]   _zz_4337;
  wire       [35:0]   _zz_4338;
  wire       [35:0]   _zz_4339;
  wire       [35:0]   _zz_4340;
  wire       [26:0]   _zz_4341;
  wire       [35:0]   _zz_4342;
  wire       [17:0]   _zz_4343;
  wire       [35:0]   _zz_4344;
  wire       [35:0]   _zz_4345;
  wire       [35:0]   _zz_4346;
  wire       [35:0]   _zz_4347;
  wire       [35:0]   _zz_4348;
  wire       [26:0]   _zz_4349;
  wire       [35:0]   _zz_4350;
  wire       [17:0]   _zz_4351;
  wire       [35:0]   _zz_4352;
  wire       [35:0]   _zz_4353;
  wire       [35:0]   _zz_4354;
  wire       [35:0]   _zz_4355;
  wire       [35:0]   _zz_4356;
  wire       [26:0]   _zz_4357;
  wire       [35:0]   _zz_4358;
  wire       [17:0]   _zz_4359;
  wire       [35:0]   _zz_4360;
  wire       [35:0]   _zz_4361;
  wire       [35:0]   _zz_4362;
  wire       [35:0]   _zz_4363;
  wire       [35:0]   _zz_4364;
  wire       [26:0]   _zz_4365;
  wire       [35:0]   _zz_4366;
  wire       [17:0]   _zz_4367;
  wire       [17:0]   _zz_4368;
  wire       [35:0]   _zz_4369;
  wire       [35:0]   _zz_4370;
  wire       [17:0]   _zz_4371;
  wire       [35:0]   _zz_4372;
  wire       [35:0]   _zz_4373;
  wire       [35:0]   _zz_4374;
  wire       [17:0]   _zz_4375;
  wire       [35:0]   _zz_4376;
  wire       [35:0]   _zz_4377;
  wire       [35:0]   _zz_4378;
  wire       [35:0]   _zz_4379;
  wire       [35:0]   _zz_4380;
  wire       [35:0]   _zz_4381;
  wire       [26:0]   _zz_4382;
  wire       [35:0]   _zz_4383;
  wire       [17:0]   _zz_4384;
  wire       [35:0]   _zz_4385;
  wire       [35:0]   _zz_4386;
  wire       [35:0]   _zz_4387;
  wire       [35:0]   _zz_4388;
  wire       [35:0]   _zz_4389;
  wire       [26:0]   _zz_4390;
  wire       [35:0]   _zz_4391;
  wire       [17:0]   _zz_4392;
  wire       [35:0]   _zz_4393;
  wire       [35:0]   _zz_4394;
  wire       [35:0]   _zz_4395;
  wire       [35:0]   _zz_4396;
  wire       [35:0]   _zz_4397;
  wire       [26:0]   _zz_4398;
  wire       [35:0]   _zz_4399;
  wire       [17:0]   _zz_4400;
  wire       [35:0]   _zz_4401;
  wire       [35:0]   _zz_4402;
  wire       [35:0]   _zz_4403;
  wire       [35:0]   _zz_4404;
  wire       [35:0]   _zz_4405;
  wire       [26:0]   _zz_4406;
  wire       [35:0]   _zz_4407;
  wire       [17:0]   _zz_4408;
  wire       [17:0]   _zz_4409;
  wire       [35:0]   _zz_4410;
  wire       [35:0]   _zz_4411;
  wire       [17:0]   _zz_4412;
  wire       [35:0]   _zz_4413;
  wire       [35:0]   _zz_4414;
  wire       [35:0]   _zz_4415;
  wire       [17:0]   _zz_4416;
  wire       [35:0]   _zz_4417;
  wire       [35:0]   _zz_4418;
  wire       [35:0]   _zz_4419;
  wire       [35:0]   _zz_4420;
  wire       [35:0]   _zz_4421;
  wire       [35:0]   _zz_4422;
  wire       [26:0]   _zz_4423;
  wire       [35:0]   _zz_4424;
  wire       [17:0]   _zz_4425;
  wire       [35:0]   _zz_4426;
  wire       [35:0]   _zz_4427;
  wire       [35:0]   _zz_4428;
  wire       [35:0]   _zz_4429;
  wire       [35:0]   _zz_4430;
  wire       [26:0]   _zz_4431;
  wire       [35:0]   _zz_4432;
  wire       [17:0]   _zz_4433;
  wire       [35:0]   _zz_4434;
  wire       [35:0]   _zz_4435;
  wire       [35:0]   _zz_4436;
  wire       [35:0]   _zz_4437;
  wire       [35:0]   _zz_4438;
  wire       [26:0]   _zz_4439;
  wire       [35:0]   _zz_4440;
  wire       [17:0]   _zz_4441;
  wire       [35:0]   _zz_4442;
  wire       [35:0]   _zz_4443;
  wire       [35:0]   _zz_4444;
  wire       [35:0]   _zz_4445;
  wire       [35:0]   _zz_4446;
  wire       [26:0]   _zz_4447;
  wire       [35:0]   _zz_4448;
  wire       [17:0]   _zz_4449;
  wire       [17:0]   _zz_4450;
  wire       [35:0]   _zz_4451;
  wire       [35:0]   _zz_4452;
  wire       [17:0]   _zz_4453;
  wire       [35:0]   _zz_4454;
  wire       [35:0]   _zz_4455;
  wire       [35:0]   _zz_4456;
  wire       [17:0]   _zz_4457;
  wire       [35:0]   _zz_4458;
  wire       [35:0]   _zz_4459;
  wire       [35:0]   _zz_4460;
  wire       [35:0]   _zz_4461;
  wire       [35:0]   _zz_4462;
  wire       [35:0]   _zz_4463;
  wire       [26:0]   _zz_4464;
  wire       [35:0]   _zz_4465;
  wire       [17:0]   _zz_4466;
  wire       [35:0]   _zz_4467;
  wire       [35:0]   _zz_4468;
  wire       [35:0]   _zz_4469;
  wire       [35:0]   _zz_4470;
  wire       [35:0]   _zz_4471;
  wire       [26:0]   _zz_4472;
  wire       [35:0]   _zz_4473;
  wire       [17:0]   _zz_4474;
  wire       [35:0]   _zz_4475;
  wire       [35:0]   _zz_4476;
  wire       [35:0]   _zz_4477;
  wire       [35:0]   _zz_4478;
  wire       [35:0]   _zz_4479;
  wire       [26:0]   _zz_4480;
  wire       [35:0]   _zz_4481;
  wire       [17:0]   _zz_4482;
  wire       [35:0]   _zz_4483;
  wire       [35:0]   _zz_4484;
  wire       [35:0]   _zz_4485;
  wire       [35:0]   _zz_4486;
  wire       [35:0]   _zz_4487;
  wire       [26:0]   _zz_4488;
  wire       [35:0]   _zz_4489;
  wire       [17:0]   _zz_4490;
  wire       [17:0]   _zz_4491;
  wire       [35:0]   _zz_4492;
  wire       [35:0]   _zz_4493;
  wire       [17:0]   _zz_4494;
  wire       [35:0]   _zz_4495;
  wire       [35:0]   _zz_4496;
  wire       [35:0]   _zz_4497;
  wire       [17:0]   _zz_4498;
  wire       [35:0]   _zz_4499;
  wire       [35:0]   _zz_4500;
  wire       [35:0]   _zz_4501;
  wire       [35:0]   _zz_4502;
  wire       [35:0]   _zz_4503;
  wire       [35:0]   _zz_4504;
  wire       [26:0]   _zz_4505;
  wire       [35:0]   _zz_4506;
  wire       [17:0]   _zz_4507;
  wire       [35:0]   _zz_4508;
  wire       [35:0]   _zz_4509;
  wire       [35:0]   _zz_4510;
  wire       [35:0]   _zz_4511;
  wire       [35:0]   _zz_4512;
  wire       [26:0]   _zz_4513;
  wire       [35:0]   _zz_4514;
  wire       [17:0]   _zz_4515;
  wire       [35:0]   _zz_4516;
  wire       [35:0]   _zz_4517;
  wire       [35:0]   _zz_4518;
  wire       [35:0]   _zz_4519;
  wire       [35:0]   _zz_4520;
  wire       [26:0]   _zz_4521;
  wire       [35:0]   _zz_4522;
  wire       [17:0]   _zz_4523;
  wire       [35:0]   _zz_4524;
  wire       [35:0]   _zz_4525;
  wire       [35:0]   _zz_4526;
  wire       [35:0]   _zz_4527;
  wire       [35:0]   _zz_4528;
  wire       [26:0]   _zz_4529;
  wire       [35:0]   _zz_4530;
  wire       [17:0]   _zz_4531;
  wire       [17:0]   _zz_4532;
  wire       [35:0]   _zz_4533;
  wire       [35:0]   _zz_4534;
  wire       [17:0]   _zz_4535;
  wire       [35:0]   _zz_4536;
  wire       [35:0]   _zz_4537;
  wire       [35:0]   _zz_4538;
  wire       [17:0]   _zz_4539;
  wire       [35:0]   _zz_4540;
  wire       [35:0]   _zz_4541;
  wire       [35:0]   _zz_4542;
  wire       [35:0]   _zz_4543;
  wire       [35:0]   _zz_4544;
  wire       [35:0]   _zz_4545;
  wire       [26:0]   _zz_4546;
  wire       [35:0]   _zz_4547;
  wire       [17:0]   _zz_4548;
  wire       [35:0]   _zz_4549;
  wire       [35:0]   _zz_4550;
  wire       [35:0]   _zz_4551;
  wire       [35:0]   _zz_4552;
  wire       [35:0]   _zz_4553;
  wire       [26:0]   _zz_4554;
  wire       [35:0]   _zz_4555;
  wire       [17:0]   _zz_4556;
  wire       [35:0]   _zz_4557;
  wire       [35:0]   _zz_4558;
  wire       [35:0]   _zz_4559;
  wire       [35:0]   _zz_4560;
  wire       [35:0]   _zz_4561;
  wire       [26:0]   _zz_4562;
  wire       [35:0]   _zz_4563;
  wire       [17:0]   _zz_4564;
  wire       [35:0]   _zz_4565;
  wire       [35:0]   _zz_4566;
  wire       [35:0]   _zz_4567;
  wire       [35:0]   _zz_4568;
  wire       [35:0]   _zz_4569;
  wire       [26:0]   _zz_4570;
  wire       [35:0]   _zz_4571;
  wire       [17:0]   _zz_4572;
  wire       [17:0]   _zz_4573;
  wire       [35:0]   _zz_4574;
  wire       [35:0]   _zz_4575;
  wire       [17:0]   _zz_4576;
  wire       [35:0]   _zz_4577;
  wire       [35:0]   _zz_4578;
  wire       [35:0]   _zz_4579;
  wire       [17:0]   _zz_4580;
  wire       [35:0]   _zz_4581;
  wire       [35:0]   _zz_4582;
  wire       [35:0]   _zz_4583;
  wire       [35:0]   _zz_4584;
  wire       [35:0]   _zz_4585;
  wire       [35:0]   _zz_4586;
  wire       [26:0]   _zz_4587;
  wire       [35:0]   _zz_4588;
  wire       [17:0]   _zz_4589;
  wire       [35:0]   _zz_4590;
  wire       [35:0]   _zz_4591;
  wire       [35:0]   _zz_4592;
  wire       [35:0]   _zz_4593;
  wire       [35:0]   _zz_4594;
  wire       [26:0]   _zz_4595;
  wire       [35:0]   _zz_4596;
  wire       [17:0]   _zz_4597;
  wire       [35:0]   _zz_4598;
  wire       [35:0]   _zz_4599;
  wire       [35:0]   _zz_4600;
  wire       [35:0]   _zz_4601;
  wire       [35:0]   _zz_4602;
  wire       [26:0]   _zz_4603;
  wire       [35:0]   _zz_4604;
  wire       [17:0]   _zz_4605;
  wire       [35:0]   _zz_4606;
  wire       [35:0]   _zz_4607;
  wire       [35:0]   _zz_4608;
  wire       [35:0]   _zz_4609;
  wire       [35:0]   _zz_4610;
  wire       [26:0]   _zz_4611;
  wire       [35:0]   _zz_4612;
  wire       [17:0]   _zz_4613;
  wire       [17:0]   _zz_4614;
  wire       [35:0]   _zz_4615;
  wire       [35:0]   _zz_4616;
  wire       [17:0]   _zz_4617;
  wire       [35:0]   _zz_4618;
  wire       [35:0]   _zz_4619;
  wire       [35:0]   _zz_4620;
  wire       [17:0]   _zz_4621;
  wire       [35:0]   _zz_4622;
  wire       [35:0]   _zz_4623;
  wire       [35:0]   _zz_4624;
  wire       [35:0]   _zz_4625;
  wire       [35:0]   _zz_4626;
  wire       [35:0]   _zz_4627;
  wire       [26:0]   _zz_4628;
  wire       [35:0]   _zz_4629;
  wire       [17:0]   _zz_4630;
  wire       [35:0]   _zz_4631;
  wire       [35:0]   _zz_4632;
  wire       [35:0]   _zz_4633;
  wire       [35:0]   _zz_4634;
  wire       [35:0]   _zz_4635;
  wire       [26:0]   _zz_4636;
  wire       [35:0]   _zz_4637;
  wire       [17:0]   _zz_4638;
  wire       [35:0]   _zz_4639;
  wire       [35:0]   _zz_4640;
  wire       [35:0]   _zz_4641;
  wire       [35:0]   _zz_4642;
  wire       [35:0]   _zz_4643;
  wire       [26:0]   _zz_4644;
  wire       [35:0]   _zz_4645;
  wire       [17:0]   _zz_4646;
  wire       [35:0]   _zz_4647;
  wire       [35:0]   _zz_4648;
  wire       [35:0]   _zz_4649;
  wire       [35:0]   _zz_4650;
  wire       [35:0]   _zz_4651;
  wire       [26:0]   _zz_4652;
  wire       [35:0]   _zz_4653;
  wire       [17:0]   _zz_4654;
  wire       [17:0]   _zz_4655;
  wire       [35:0]   _zz_4656;
  wire       [35:0]   _zz_4657;
  wire       [17:0]   _zz_4658;
  wire       [35:0]   _zz_4659;
  wire       [35:0]   _zz_4660;
  wire       [35:0]   _zz_4661;
  wire       [17:0]   _zz_4662;
  wire       [35:0]   _zz_4663;
  wire       [35:0]   _zz_4664;
  wire       [35:0]   _zz_4665;
  wire       [35:0]   _zz_4666;
  wire       [35:0]   _zz_4667;
  wire       [35:0]   _zz_4668;
  wire       [26:0]   _zz_4669;
  wire       [35:0]   _zz_4670;
  wire       [17:0]   _zz_4671;
  wire       [35:0]   _zz_4672;
  wire       [35:0]   _zz_4673;
  wire       [35:0]   _zz_4674;
  wire       [35:0]   _zz_4675;
  wire       [35:0]   _zz_4676;
  wire       [26:0]   _zz_4677;
  wire       [35:0]   _zz_4678;
  wire       [17:0]   _zz_4679;
  wire       [35:0]   _zz_4680;
  wire       [35:0]   _zz_4681;
  wire       [35:0]   _zz_4682;
  wire       [35:0]   _zz_4683;
  wire       [35:0]   _zz_4684;
  wire       [26:0]   _zz_4685;
  wire       [35:0]   _zz_4686;
  wire       [17:0]   _zz_4687;
  wire       [35:0]   _zz_4688;
  wire       [35:0]   _zz_4689;
  wire       [35:0]   _zz_4690;
  wire       [35:0]   _zz_4691;
  wire       [35:0]   _zz_4692;
  wire       [26:0]   _zz_4693;
  wire       [35:0]   _zz_4694;
  wire       [17:0]   _zz_4695;
  wire       [17:0]   _zz_4696;
  wire       [35:0]   _zz_4697;
  wire       [35:0]   _zz_4698;
  wire       [17:0]   _zz_4699;
  wire       [35:0]   _zz_4700;
  wire       [35:0]   _zz_4701;
  wire       [35:0]   _zz_4702;
  wire       [17:0]   _zz_4703;
  wire       [35:0]   _zz_4704;
  wire       [35:0]   _zz_4705;
  wire       [35:0]   _zz_4706;
  wire       [35:0]   _zz_4707;
  wire       [35:0]   _zz_4708;
  wire       [35:0]   _zz_4709;
  wire       [26:0]   _zz_4710;
  wire       [35:0]   _zz_4711;
  wire       [17:0]   _zz_4712;
  wire       [35:0]   _zz_4713;
  wire       [35:0]   _zz_4714;
  wire       [35:0]   _zz_4715;
  wire       [35:0]   _zz_4716;
  wire       [35:0]   _zz_4717;
  wire       [26:0]   _zz_4718;
  wire       [35:0]   _zz_4719;
  wire       [17:0]   _zz_4720;
  wire       [35:0]   _zz_4721;
  wire       [35:0]   _zz_4722;
  wire       [35:0]   _zz_4723;
  wire       [35:0]   _zz_4724;
  wire       [35:0]   _zz_4725;
  wire       [26:0]   _zz_4726;
  wire       [35:0]   _zz_4727;
  wire       [17:0]   _zz_4728;
  wire       [35:0]   _zz_4729;
  wire       [35:0]   _zz_4730;
  wire       [35:0]   _zz_4731;
  wire       [35:0]   _zz_4732;
  wire       [35:0]   _zz_4733;
  wire       [26:0]   _zz_4734;
  wire       [35:0]   _zz_4735;
  wire       [17:0]   _zz_4736;
  wire       [17:0]   _zz_4737;
  wire       [35:0]   _zz_4738;
  wire       [35:0]   _zz_4739;
  wire       [17:0]   _zz_4740;
  wire       [35:0]   _zz_4741;
  wire       [35:0]   _zz_4742;
  wire       [35:0]   _zz_4743;
  wire       [17:0]   _zz_4744;
  wire       [35:0]   _zz_4745;
  wire       [35:0]   _zz_4746;
  wire       [35:0]   _zz_4747;
  wire       [35:0]   _zz_4748;
  wire       [35:0]   _zz_4749;
  wire       [35:0]   _zz_4750;
  wire       [26:0]   _zz_4751;
  wire       [35:0]   _zz_4752;
  wire       [17:0]   _zz_4753;
  wire       [35:0]   _zz_4754;
  wire       [35:0]   _zz_4755;
  wire       [35:0]   _zz_4756;
  wire       [35:0]   _zz_4757;
  wire       [35:0]   _zz_4758;
  wire       [26:0]   _zz_4759;
  wire       [35:0]   _zz_4760;
  wire       [17:0]   _zz_4761;
  wire       [35:0]   _zz_4762;
  wire       [35:0]   _zz_4763;
  wire       [35:0]   _zz_4764;
  wire       [35:0]   _zz_4765;
  wire       [35:0]   _zz_4766;
  wire       [26:0]   _zz_4767;
  wire       [35:0]   _zz_4768;
  wire       [17:0]   _zz_4769;
  wire       [35:0]   _zz_4770;
  wire       [35:0]   _zz_4771;
  wire       [35:0]   _zz_4772;
  wire       [35:0]   _zz_4773;
  wire       [35:0]   _zz_4774;
  wire       [26:0]   _zz_4775;
  wire       [35:0]   _zz_4776;
  wire       [17:0]   _zz_4777;
  wire       [17:0]   _zz_4778;
  wire       [35:0]   _zz_4779;
  wire       [35:0]   _zz_4780;
  wire       [17:0]   _zz_4781;
  wire       [35:0]   _zz_4782;
  wire       [35:0]   _zz_4783;
  wire       [35:0]   _zz_4784;
  wire       [17:0]   _zz_4785;
  wire       [35:0]   _zz_4786;
  wire       [35:0]   _zz_4787;
  wire       [35:0]   _zz_4788;
  wire       [35:0]   _zz_4789;
  wire       [35:0]   _zz_4790;
  wire       [35:0]   _zz_4791;
  wire       [26:0]   _zz_4792;
  wire       [35:0]   _zz_4793;
  wire       [17:0]   _zz_4794;
  wire       [35:0]   _zz_4795;
  wire       [35:0]   _zz_4796;
  wire       [35:0]   _zz_4797;
  wire       [35:0]   _zz_4798;
  wire       [35:0]   _zz_4799;
  wire       [26:0]   _zz_4800;
  wire       [35:0]   _zz_4801;
  wire       [17:0]   _zz_4802;
  wire       [35:0]   _zz_4803;
  wire       [35:0]   _zz_4804;
  wire       [35:0]   _zz_4805;
  wire       [35:0]   _zz_4806;
  wire       [35:0]   _zz_4807;
  wire       [26:0]   _zz_4808;
  wire       [35:0]   _zz_4809;
  wire       [17:0]   _zz_4810;
  wire       [35:0]   _zz_4811;
  wire       [35:0]   _zz_4812;
  wire       [35:0]   _zz_4813;
  wire       [35:0]   _zz_4814;
  wire       [35:0]   _zz_4815;
  wire       [26:0]   _zz_4816;
  wire       [35:0]   _zz_4817;
  wire       [17:0]   _zz_4818;
  wire       [17:0]   _zz_4819;
  wire       [35:0]   _zz_4820;
  wire       [35:0]   _zz_4821;
  wire       [17:0]   _zz_4822;
  wire       [35:0]   _zz_4823;
  wire       [35:0]   _zz_4824;
  wire       [35:0]   _zz_4825;
  wire       [17:0]   _zz_4826;
  wire       [35:0]   _zz_4827;
  wire       [35:0]   _zz_4828;
  wire       [35:0]   _zz_4829;
  wire       [35:0]   _zz_4830;
  wire       [35:0]   _zz_4831;
  wire       [35:0]   _zz_4832;
  wire       [26:0]   _zz_4833;
  wire       [35:0]   _zz_4834;
  wire       [17:0]   _zz_4835;
  wire       [35:0]   _zz_4836;
  wire       [35:0]   _zz_4837;
  wire       [35:0]   _zz_4838;
  wire       [35:0]   _zz_4839;
  wire       [35:0]   _zz_4840;
  wire       [26:0]   _zz_4841;
  wire       [35:0]   _zz_4842;
  wire       [17:0]   _zz_4843;
  wire       [35:0]   _zz_4844;
  wire       [35:0]   _zz_4845;
  wire       [35:0]   _zz_4846;
  wire       [35:0]   _zz_4847;
  wire       [35:0]   _zz_4848;
  wire       [26:0]   _zz_4849;
  wire       [35:0]   _zz_4850;
  wire       [17:0]   _zz_4851;
  wire       [35:0]   _zz_4852;
  wire       [35:0]   _zz_4853;
  wire       [35:0]   _zz_4854;
  wire       [35:0]   _zz_4855;
  wire       [35:0]   _zz_4856;
  wire       [26:0]   _zz_4857;
  wire       [35:0]   _zz_4858;
  wire       [17:0]   _zz_4859;
  wire       [17:0]   _zz_4860;
  wire       [35:0]   _zz_4861;
  wire       [35:0]   _zz_4862;
  wire       [17:0]   _zz_4863;
  wire       [35:0]   _zz_4864;
  wire       [35:0]   _zz_4865;
  wire       [35:0]   _zz_4866;
  wire       [17:0]   _zz_4867;
  wire       [35:0]   _zz_4868;
  wire       [35:0]   _zz_4869;
  wire       [35:0]   _zz_4870;
  wire       [35:0]   _zz_4871;
  wire       [35:0]   _zz_4872;
  wire       [35:0]   _zz_4873;
  wire       [26:0]   _zz_4874;
  wire       [35:0]   _zz_4875;
  wire       [17:0]   _zz_4876;
  wire       [35:0]   _zz_4877;
  wire       [35:0]   _zz_4878;
  wire       [35:0]   _zz_4879;
  wire       [35:0]   _zz_4880;
  wire       [35:0]   _zz_4881;
  wire       [26:0]   _zz_4882;
  wire       [35:0]   _zz_4883;
  wire       [17:0]   _zz_4884;
  wire       [35:0]   _zz_4885;
  wire       [35:0]   _zz_4886;
  wire       [35:0]   _zz_4887;
  wire       [35:0]   _zz_4888;
  wire       [35:0]   _zz_4889;
  wire       [26:0]   _zz_4890;
  wire       [35:0]   _zz_4891;
  wire       [17:0]   _zz_4892;
  wire       [35:0]   _zz_4893;
  wire       [35:0]   _zz_4894;
  wire       [35:0]   _zz_4895;
  wire       [35:0]   _zz_4896;
  wire       [35:0]   _zz_4897;
  wire       [26:0]   _zz_4898;
  wire       [35:0]   _zz_4899;
  wire       [17:0]   _zz_4900;
  wire       [17:0]   _zz_4901;
  wire       [35:0]   _zz_4902;
  wire       [35:0]   _zz_4903;
  wire       [17:0]   _zz_4904;
  wire       [35:0]   _zz_4905;
  wire       [35:0]   _zz_4906;
  wire       [35:0]   _zz_4907;
  wire       [17:0]   _zz_4908;
  wire       [35:0]   _zz_4909;
  wire       [35:0]   _zz_4910;
  wire       [35:0]   _zz_4911;
  wire       [35:0]   _zz_4912;
  wire       [35:0]   _zz_4913;
  wire       [35:0]   _zz_4914;
  wire       [26:0]   _zz_4915;
  wire       [35:0]   _zz_4916;
  wire       [17:0]   _zz_4917;
  wire       [35:0]   _zz_4918;
  wire       [35:0]   _zz_4919;
  wire       [35:0]   _zz_4920;
  wire       [35:0]   _zz_4921;
  wire       [35:0]   _zz_4922;
  wire       [26:0]   _zz_4923;
  wire       [35:0]   _zz_4924;
  wire       [17:0]   _zz_4925;
  wire       [35:0]   _zz_4926;
  wire       [35:0]   _zz_4927;
  wire       [35:0]   _zz_4928;
  wire       [35:0]   _zz_4929;
  wire       [35:0]   _zz_4930;
  wire       [26:0]   _zz_4931;
  wire       [35:0]   _zz_4932;
  wire       [17:0]   _zz_4933;
  wire       [35:0]   _zz_4934;
  wire       [35:0]   _zz_4935;
  wire       [35:0]   _zz_4936;
  wire       [35:0]   _zz_4937;
  wire       [35:0]   _zz_4938;
  wire       [26:0]   _zz_4939;
  wire       [35:0]   _zz_4940;
  wire       [17:0]   _zz_4941;
  wire       [17:0]   _zz_4942;
  wire       [35:0]   _zz_4943;
  wire       [35:0]   _zz_4944;
  wire       [17:0]   _zz_4945;
  wire       [35:0]   _zz_4946;
  wire       [35:0]   _zz_4947;
  wire       [35:0]   _zz_4948;
  wire       [17:0]   _zz_4949;
  wire       [35:0]   _zz_4950;
  wire       [35:0]   _zz_4951;
  wire       [35:0]   _zz_4952;
  wire       [35:0]   _zz_4953;
  wire       [35:0]   _zz_4954;
  wire       [35:0]   _zz_4955;
  wire       [26:0]   _zz_4956;
  wire       [35:0]   _zz_4957;
  wire       [17:0]   _zz_4958;
  wire       [35:0]   _zz_4959;
  wire       [35:0]   _zz_4960;
  wire       [35:0]   _zz_4961;
  wire       [35:0]   _zz_4962;
  wire       [35:0]   _zz_4963;
  wire       [26:0]   _zz_4964;
  wire       [35:0]   _zz_4965;
  wire       [17:0]   _zz_4966;
  wire       [35:0]   _zz_4967;
  wire       [35:0]   _zz_4968;
  wire       [35:0]   _zz_4969;
  wire       [35:0]   _zz_4970;
  wire       [35:0]   _zz_4971;
  wire       [26:0]   _zz_4972;
  wire       [35:0]   _zz_4973;
  wire       [17:0]   _zz_4974;
  wire       [35:0]   _zz_4975;
  wire       [35:0]   _zz_4976;
  wire       [35:0]   _zz_4977;
  wire       [35:0]   _zz_4978;
  wire       [35:0]   _zz_4979;
  wire       [26:0]   _zz_4980;
  wire       [35:0]   _zz_4981;
  wire       [17:0]   _zz_4982;
  wire       [17:0]   _zz_4983;
  wire       [35:0]   _zz_4984;
  wire       [35:0]   _zz_4985;
  wire       [17:0]   _zz_4986;
  wire       [35:0]   _zz_4987;
  wire       [35:0]   _zz_4988;
  wire       [35:0]   _zz_4989;
  wire       [17:0]   _zz_4990;
  wire       [35:0]   _zz_4991;
  wire       [35:0]   _zz_4992;
  wire       [35:0]   _zz_4993;
  wire       [35:0]   _zz_4994;
  wire       [35:0]   _zz_4995;
  wire       [35:0]   _zz_4996;
  wire       [26:0]   _zz_4997;
  wire       [35:0]   _zz_4998;
  wire       [17:0]   _zz_4999;
  wire       [35:0]   _zz_5000;
  wire       [35:0]   _zz_5001;
  wire       [35:0]   _zz_5002;
  wire       [35:0]   _zz_5003;
  wire       [35:0]   _zz_5004;
  wire       [26:0]   _zz_5005;
  wire       [35:0]   _zz_5006;
  wire       [17:0]   _zz_5007;
  wire       [35:0]   _zz_5008;
  wire       [35:0]   _zz_5009;
  wire       [35:0]   _zz_5010;
  wire       [35:0]   _zz_5011;
  wire       [35:0]   _zz_5012;
  wire       [26:0]   _zz_5013;
  wire       [35:0]   _zz_5014;
  wire       [17:0]   _zz_5015;
  wire       [35:0]   _zz_5016;
  wire       [35:0]   _zz_5017;
  wire       [35:0]   _zz_5018;
  wire       [35:0]   _zz_5019;
  wire       [35:0]   _zz_5020;
  wire       [26:0]   _zz_5021;
  wire       [35:0]   _zz_5022;
  wire       [17:0]   _zz_5023;
  wire       [17:0]   _zz_5024;
  wire       [35:0]   _zz_5025;
  wire       [35:0]   _zz_5026;
  wire       [17:0]   _zz_5027;
  wire       [35:0]   _zz_5028;
  wire       [35:0]   _zz_5029;
  wire       [35:0]   _zz_5030;
  wire       [17:0]   _zz_5031;
  wire       [35:0]   _zz_5032;
  wire       [35:0]   _zz_5033;
  wire       [35:0]   _zz_5034;
  wire       [35:0]   _zz_5035;
  wire       [35:0]   _zz_5036;
  wire       [35:0]   _zz_5037;
  wire       [26:0]   _zz_5038;
  wire       [35:0]   _zz_5039;
  wire       [17:0]   _zz_5040;
  wire       [35:0]   _zz_5041;
  wire       [35:0]   _zz_5042;
  wire       [35:0]   _zz_5043;
  wire       [35:0]   _zz_5044;
  wire       [35:0]   _zz_5045;
  wire       [26:0]   _zz_5046;
  wire       [35:0]   _zz_5047;
  wire       [17:0]   _zz_5048;
  wire       [35:0]   _zz_5049;
  wire       [35:0]   _zz_5050;
  wire       [35:0]   _zz_5051;
  wire       [35:0]   _zz_5052;
  wire       [35:0]   _zz_5053;
  wire       [26:0]   _zz_5054;
  wire       [35:0]   _zz_5055;
  wire       [17:0]   _zz_5056;
  wire       [35:0]   _zz_5057;
  wire       [35:0]   _zz_5058;
  wire       [35:0]   _zz_5059;
  wire       [35:0]   _zz_5060;
  wire       [35:0]   _zz_5061;
  wire       [26:0]   _zz_5062;
  wire       [35:0]   _zz_5063;
  wire       [17:0]   _zz_5064;
  wire       [17:0]   _zz_5065;
  wire       [35:0]   _zz_5066;
  wire       [35:0]   _zz_5067;
  wire       [17:0]   _zz_5068;
  wire       [35:0]   _zz_5069;
  wire       [35:0]   _zz_5070;
  wire       [35:0]   _zz_5071;
  wire       [17:0]   _zz_5072;
  wire       [35:0]   _zz_5073;
  wire       [35:0]   _zz_5074;
  wire       [35:0]   _zz_5075;
  wire       [35:0]   _zz_5076;
  wire       [35:0]   _zz_5077;
  wire       [35:0]   _zz_5078;
  wire       [26:0]   _zz_5079;
  wire       [35:0]   _zz_5080;
  wire       [17:0]   _zz_5081;
  wire       [35:0]   _zz_5082;
  wire       [35:0]   _zz_5083;
  wire       [35:0]   _zz_5084;
  wire       [35:0]   _zz_5085;
  wire       [35:0]   _zz_5086;
  wire       [26:0]   _zz_5087;
  wire       [35:0]   _zz_5088;
  wire       [17:0]   _zz_5089;
  wire       [35:0]   _zz_5090;
  wire       [35:0]   _zz_5091;
  wire       [35:0]   _zz_5092;
  wire       [35:0]   _zz_5093;
  wire       [35:0]   _zz_5094;
  wire       [26:0]   _zz_5095;
  wire       [35:0]   _zz_5096;
  wire       [17:0]   _zz_5097;
  wire       [35:0]   _zz_5098;
  wire       [35:0]   _zz_5099;
  wire       [35:0]   _zz_5100;
  wire       [35:0]   _zz_5101;
  wire       [35:0]   _zz_5102;
  wire       [26:0]   _zz_5103;
  wire       [35:0]   _zz_5104;
  wire       [17:0]   _zz_5105;
  wire       [17:0]   _zz_5106;
  wire       [35:0]   _zz_5107;
  wire       [35:0]   _zz_5108;
  wire       [17:0]   _zz_5109;
  wire       [35:0]   _zz_5110;
  wire       [35:0]   _zz_5111;
  wire       [35:0]   _zz_5112;
  wire       [17:0]   _zz_5113;
  wire       [35:0]   _zz_5114;
  wire       [35:0]   _zz_5115;
  wire       [35:0]   _zz_5116;
  wire       [35:0]   _zz_5117;
  wire       [35:0]   _zz_5118;
  wire       [35:0]   _zz_5119;
  wire       [26:0]   _zz_5120;
  wire       [35:0]   _zz_5121;
  wire       [17:0]   _zz_5122;
  wire       [35:0]   _zz_5123;
  wire       [35:0]   _zz_5124;
  wire       [35:0]   _zz_5125;
  wire       [35:0]   _zz_5126;
  wire       [35:0]   _zz_5127;
  wire       [26:0]   _zz_5128;
  wire       [35:0]   _zz_5129;
  wire       [17:0]   _zz_5130;
  wire       [35:0]   _zz_5131;
  wire       [35:0]   _zz_5132;
  wire       [35:0]   _zz_5133;
  wire       [35:0]   _zz_5134;
  wire       [35:0]   _zz_5135;
  wire       [26:0]   _zz_5136;
  wire       [35:0]   _zz_5137;
  wire       [17:0]   _zz_5138;
  wire       [35:0]   _zz_5139;
  wire       [35:0]   _zz_5140;
  wire       [35:0]   _zz_5141;
  wire       [35:0]   _zz_5142;
  wire       [35:0]   _zz_5143;
  wire       [26:0]   _zz_5144;
  wire       [35:0]   _zz_5145;
  wire       [17:0]   _zz_5146;
  wire       [17:0]   _zz_5147;
  wire       [35:0]   _zz_5148;
  wire       [35:0]   _zz_5149;
  wire       [17:0]   _zz_5150;
  wire       [35:0]   _zz_5151;
  wire       [35:0]   _zz_5152;
  wire       [35:0]   _zz_5153;
  wire       [17:0]   _zz_5154;
  wire       [35:0]   _zz_5155;
  wire       [35:0]   _zz_5156;
  wire       [35:0]   _zz_5157;
  wire       [35:0]   _zz_5158;
  wire       [35:0]   _zz_5159;
  wire       [35:0]   _zz_5160;
  wire       [26:0]   _zz_5161;
  wire       [35:0]   _zz_5162;
  wire       [17:0]   _zz_5163;
  wire       [35:0]   _zz_5164;
  wire       [35:0]   _zz_5165;
  wire       [35:0]   _zz_5166;
  wire       [35:0]   _zz_5167;
  wire       [35:0]   _zz_5168;
  wire       [26:0]   _zz_5169;
  wire       [35:0]   _zz_5170;
  wire       [17:0]   _zz_5171;
  wire       [35:0]   _zz_5172;
  wire       [35:0]   _zz_5173;
  wire       [35:0]   _zz_5174;
  wire       [35:0]   _zz_5175;
  wire       [35:0]   _zz_5176;
  wire       [26:0]   _zz_5177;
  wire       [35:0]   _zz_5178;
  wire       [17:0]   _zz_5179;
  wire       [35:0]   _zz_5180;
  wire       [35:0]   _zz_5181;
  wire       [35:0]   _zz_5182;
  wire       [35:0]   _zz_5183;
  wire       [35:0]   _zz_5184;
  wire       [26:0]   _zz_5185;
  wire       [35:0]   _zz_5186;
  wire       [17:0]   _zz_5187;
  wire       [17:0]   _zz_5188;
  wire       [35:0]   _zz_5189;
  wire       [35:0]   _zz_5190;
  wire       [17:0]   _zz_5191;
  wire       [35:0]   _zz_5192;
  wire       [35:0]   _zz_5193;
  wire       [35:0]   _zz_5194;
  wire       [17:0]   _zz_5195;
  wire       [35:0]   _zz_5196;
  wire       [35:0]   _zz_5197;
  wire       [35:0]   _zz_5198;
  wire       [35:0]   _zz_5199;
  wire       [35:0]   _zz_5200;
  wire       [35:0]   _zz_5201;
  wire       [26:0]   _zz_5202;
  wire       [35:0]   _zz_5203;
  wire       [17:0]   _zz_5204;
  wire       [35:0]   _zz_5205;
  wire       [35:0]   _zz_5206;
  wire       [35:0]   _zz_5207;
  wire       [35:0]   _zz_5208;
  wire       [35:0]   _zz_5209;
  wire       [26:0]   _zz_5210;
  wire       [35:0]   _zz_5211;
  wire       [17:0]   _zz_5212;
  wire       [35:0]   _zz_5213;
  wire       [35:0]   _zz_5214;
  wire       [35:0]   _zz_5215;
  wire       [35:0]   _zz_5216;
  wire       [35:0]   _zz_5217;
  wire       [26:0]   _zz_5218;
  wire       [35:0]   _zz_5219;
  wire       [17:0]   _zz_5220;
  wire       [35:0]   _zz_5221;
  wire       [35:0]   _zz_5222;
  wire       [35:0]   _zz_5223;
  wire       [35:0]   _zz_5224;
  wire       [35:0]   _zz_5225;
  wire       [26:0]   _zz_5226;
  wire       [35:0]   _zz_5227;
  wire       [17:0]   _zz_5228;
  wire       [17:0]   _zz_5229;
  wire       [35:0]   _zz_5230;
  wire       [35:0]   _zz_5231;
  wire       [17:0]   _zz_5232;
  wire       [35:0]   _zz_5233;
  wire       [35:0]   _zz_5234;
  wire       [35:0]   _zz_5235;
  wire       [17:0]   _zz_5236;
  wire       [35:0]   _zz_5237;
  wire       [35:0]   _zz_5238;
  wire       [35:0]   _zz_5239;
  wire       [35:0]   _zz_5240;
  wire       [35:0]   _zz_5241;
  wire       [35:0]   _zz_5242;
  wire       [26:0]   _zz_5243;
  wire       [35:0]   _zz_5244;
  wire       [17:0]   _zz_5245;
  wire       [35:0]   _zz_5246;
  wire       [35:0]   _zz_5247;
  wire       [35:0]   _zz_5248;
  wire       [35:0]   _zz_5249;
  wire       [35:0]   _zz_5250;
  wire       [26:0]   _zz_5251;
  wire       [35:0]   _zz_5252;
  wire       [17:0]   _zz_5253;
  wire       [35:0]   _zz_5254;
  wire       [35:0]   _zz_5255;
  wire       [35:0]   _zz_5256;
  wire       [35:0]   _zz_5257;
  wire       [35:0]   _zz_5258;
  wire       [26:0]   _zz_5259;
  wire       [35:0]   _zz_5260;
  wire       [17:0]   _zz_5261;
  wire       [35:0]   _zz_5262;
  wire       [35:0]   _zz_5263;
  wire       [35:0]   _zz_5264;
  wire       [35:0]   _zz_5265;
  wire       [35:0]   _zz_5266;
  wire       [26:0]   _zz_5267;
  wire       [35:0]   _zz_5268;
  wire       [17:0]   _zz_5269;
  wire       [17:0]   _zz_5270;
  wire       [35:0]   _zz_5271;
  wire       [35:0]   _zz_5272;
  wire       [17:0]   _zz_5273;
  wire       [35:0]   _zz_5274;
  wire       [35:0]   _zz_5275;
  wire       [35:0]   _zz_5276;
  wire       [17:0]   _zz_5277;
  wire       [35:0]   _zz_5278;
  wire       [35:0]   _zz_5279;
  wire       [35:0]   _zz_5280;
  wire       [35:0]   _zz_5281;
  wire       [35:0]   _zz_5282;
  wire       [35:0]   _zz_5283;
  wire       [26:0]   _zz_5284;
  wire       [35:0]   _zz_5285;
  wire       [17:0]   _zz_5286;
  wire       [35:0]   _zz_5287;
  wire       [35:0]   _zz_5288;
  wire       [35:0]   _zz_5289;
  wire       [35:0]   _zz_5290;
  wire       [35:0]   _zz_5291;
  wire       [26:0]   _zz_5292;
  wire       [35:0]   _zz_5293;
  wire       [17:0]   _zz_5294;
  wire       [35:0]   _zz_5295;
  wire       [35:0]   _zz_5296;
  wire       [35:0]   _zz_5297;
  wire       [35:0]   _zz_5298;
  wire       [35:0]   _zz_5299;
  wire       [26:0]   _zz_5300;
  wire       [35:0]   _zz_5301;
  wire       [17:0]   _zz_5302;
  wire       [35:0]   _zz_5303;
  wire       [35:0]   _zz_5304;
  wire       [35:0]   _zz_5305;
  wire       [35:0]   _zz_5306;
  wire       [35:0]   _zz_5307;
  wire       [26:0]   _zz_5308;
  wire       [35:0]   _zz_5309;
  wire       [17:0]   _zz_5310;
  wire       [17:0]   _zz_5311;
  wire       [35:0]   _zz_5312;
  wire       [35:0]   _zz_5313;
  wire       [17:0]   _zz_5314;
  wire       [35:0]   _zz_5315;
  wire       [35:0]   _zz_5316;
  wire       [35:0]   _zz_5317;
  wire       [17:0]   _zz_5318;
  wire       [35:0]   _zz_5319;
  wire       [35:0]   _zz_5320;
  wire       [35:0]   _zz_5321;
  wire       [35:0]   _zz_5322;
  wire       [35:0]   _zz_5323;
  wire       [35:0]   _zz_5324;
  wire       [26:0]   _zz_5325;
  wire       [35:0]   _zz_5326;
  wire       [17:0]   _zz_5327;
  wire       [35:0]   _zz_5328;
  wire       [35:0]   _zz_5329;
  wire       [35:0]   _zz_5330;
  wire       [35:0]   _zz_5331;
  wire       [35:0]   _zz_5332;
  wire       [26:0]   _zz_5333;
  wire       [35:0]   _zz_5334;
  wire       [17:0]   _zz_5335;
  wire       [35:0]   _zz_5336;
  wire       [35:0]   _zz_5337;
  wire       [35:0]   _zz_5338;
  wire       [35:0]   _zz_5339;
  wire       [35:0]   _zz_5340;
  wire       [26:0]   _zz_5341;
  wire       [35:0]   _zz_5342;
  wire       [17:0]   _zz_5343;
  wire       [35:0]   _zz_5344;
  wire       [35:0]   _zz_5345;
  wire       [35:0]   _zz_5346;
  wire       [35:0]   _zz_5347;
  wire       [35:0]   _zz_5348;
  wire       [26:0]   _zz_5349;
  wire       [35:0]   _zz_5350;
  wire       [17:0]   _zz_5351;
  wire       [17:0]   _zz_5352;
  wire       [35:0]   _zz_5353;
  wire       [35:0]   _zz_5354;
  wire       [17:0]   _zz_5355;
  wire       [35:0]   _zz_5356;
  wire       [35:0]   _zz_5357;
  wire       [35:0]   _zz_5358;
  wire       [17:0]   _zz_5359;
  wire       [35:0]   _zz_5360;
  wire       [35:0]   _zz_5361;
  wire       [35:0]   _zz_5362;
  wire       [35:0]   _zz_5363;
  wire       [35:0]   _zz_5364;
  wire       [35:0]   _zz_5365;
  wire       [26:0]   _zz_5366;
  wire       [35:0]   _zz_5367;
  wire       [17:0]   _zz_5368;
  wire       [35:0]   _zz_5369;
  wire       [35:0]   _zz_5370;
  wire       [35:0]   _zz_5371;
  wire       [35:0]   _zz_5372;
  wire       [35:0]   _zz_5373;
  wire       [26:0]   _zz_5374;
  wire       [35:0]   _zz_5375;
  wire       [17:0]   _zz_5376;
  wire       [35:0]   _zz_5377;
  wire       [35:0]   _zz_5378;
  wire       [35:0]   _zz_5379;
  wire       [35:0]   _zz_5380;
  wire       [35:0]   _zz_5381;
  wire       [26:0]   _zz_5382;
  wire       [35:0]   _zz_5383;
  wire       [17:0]   _zz_5384;
  wire       [35:0]   _zz_5385;
  wire       [35:0]   _zz_5386;
  wire       [35:0]   _zz_5387;
  wire       [35:0]   _zz_5388;
  wire       [35:0]   _zz_5389;
  wire       [26:0]   _zz_5390;
  wire       [35:0]   _zz_5391;
  wire       [17:0]   _zz_5392;
  wire       [17:0]   _zz_5393;
  wire       [35:0]   _zz_5394;
  wire       [35:0]   _zz_5395;
  wire       [17:0]   _zz_5396;
  wire       [35:0]   _zz_5397;
  wire       [35:0]   _zz_5398;
  wire       [35:0]   _zz_5399;
  wire       [17:0]   _zz_5400;
  wire       [35:0]   _zz_5401;
  wire       [35:0]   _zz_5402;
  wire       [35:0]   _zz_5403;
  wire       [35:0]   _zz_5404;
  wire       [35:0]   _zz_5405;
  wire       [35:0]   _zz_5406;
  wire       [26:0]   _zz_5407;
  wire       [35:0]   _zz_5408;
  wire       [17:0]   _zz_5409;
  wire       [35:0]   _zz_5410;
  wire       [35:0]   _zz_5411;
  wire       [35:0]   _zz_5412;
  wire       [35:0]   _zz_5413;
  wire       [35:0]   _zz_5414;
  wire       [26:0]   _zz_5415;
  wire       [35:0]   _zz_5416;
  wire       [17:0]   _zz_5417;
  wire       [35:0]   _zz_5418;
  wire       [35:0]   _zz_5419;
  wire       [35:0]   _zz_5420;
  wire       [35:0]   _zz_5421;
  wire       [35:0]   _zz_5422;
  wire       [26:0]   _zz_5423;
  wire       [35:0]   _zz_5424;
  wire       [17:0]   _zz_5425;
  wire       [35:0]   _zz_5426;
  wire       [35:0]   _zz_5427;
  wire       [35:0]   _zz_5428;
  wire       [35:0]   _zz_5429;
  wire       [35:0]   _zz_5430;
  wire       [26:0]   _zz_5431;
  wire       [35:0]   _zz_5432;
  wire       [17:0]   _zz_5433;
  wire       [17:0]   _zz_5434;
  wire       [35:0]   _zz_5435;
  wire       [35:0]   _zz_5436;
  wire       [17:0]   _zz_5437;
  wire       [35:0]   _zz_5438;
  wire       [35:0]   _zz_5439;
  wire       [35:0]   _zz_5440;
  wire       [17:0]   _zz_5441;
  wire       [35:0]   _zz_5442;
  wire       [35:0]   _zz_5443;
  wire       [35:0]   _zz_5444;
  wire       [35:0]   _zz_5445;
  wire       [35:0]   _zz_5446;
  wire       [35:0]   _zz_5447;
  wire       [26:0]   _zz_5448;
  wire       [35:0]   _zz_5449;
  wire       [17:0]   _zz_5450;
  wire       [35:0]   _zz_5451;
  wire       [35:0]   _zz_5452;
  wire       [35:0]   _zz_5453;
  wire       [35:0]   _zz_5454;
  wire       [35:0]   _zz_5455;
  wire       [26:0]   _zz_5456;
  wire       [35:0]   _zz_5457;
  wire       [17:0]   _zz_5458;
  wire       [35:0]   _zz_5459;
  wire       [35:0]   _zz_5460;
  wire       [35:0]   _zz_5461;
  wire       [35:0]   _zz_5462;
  wire       [35:0]   _zz_5463;
  wire       [26:0]   _zz_5464;
  wire       [35:0]   _zz_5465;
  wire       [17:0]   _zz_5466;
  wire       [35:0]   _zz_5467;
  wire       [35:0]   _zz_5468;
  wire       [35:0]   _zz_5469;
  wire       [35:0]   _zz_5470;
  wire       [35:0]   _zz_5471;
  wire       [26:0]   _zz_5472;
  wire       [35:0]   _zz_5473;
  wire       [17:0]   _zz_5474;
  wire       [17:0]   _zz_5475;
  wire       [35:0]   _zz_5476;
  wire       [35:0]   _zz_5477;
  wire       [17:0]   _zz_5478;
  wire       [35:0]   _zz_5479;
  wire       [35:0]   _zz_5480;
  wire       [35:0]   _zz_5481;
  wire       [17:0]   _zz_5482;
  wire       [35:0]   _zz_5483;
  wire       [35:0]   _zz_5484;
  wire       [35:0]   _zz_5485;
  wire       [35:0]   _zz_5486;
  wire       [35:0]   _zz_5487;
  wire       [35:0]   _zz_5488;
  wire       [26:0]   _zz_5489;
  wire       [35:0]   _zz_5490;
  wire       [17:0]   _zz_5491;
  wire       [35:0]   _zz_5492;
  wire       [35:0]   _zz_5493;
  wire       [35:0]   _zz_5494;
  wire       [35:0]   _zz_5495;
  wire       [35:0]   _zz_5496;
  wire       [26:0]   _zz_5497;
  wire       [35:0]   _zz_5498;
  wire       [17:0]   _zz_5499;
  wire       [35:0]   _zz_5500;
  wire       [35:0]   _zz_5501;
  wire       [35:0]   _zz_5502;
  wire       [35:0]   _zz_5503;
  wire       [35:0]   _zz_5504;
  wire       [26:0]   _zz_5505;
  wire       [35:0]   _zz_5506;
  wire       [17:0]   _zz_5507;
  wire       [35:0]   _zz_5508;
  wire       [35:0]   _zz_5509;
  wire       [35:0]   _zz_5510;
  wire       [35:0]   _zz_5511;
  wire       [35:0]   _zz_5512;
  wire       [26:0]   _zz_5513;
  wire       [35:0]   _zz_5514;
  wire       [17:0]   _zz_5515;
  wire       [17:0]   _zz_5516;
  wire       [35:0]   _zz_5517;
  wire       [35:0]   _zz_5518;
  wire       [17:0]   _zz_5519;
  wire       [35:0]   _zz_5520;
  wire       [35:0]   _zz_5521;
  wire       [35:0]   _zz_5522;
  wire       [17:0]   _zz_5523;
  wire       [35:0]   _zz_5524;
  wire       [35:0]   _zz_5525;
  wire       [35:0]   _zz_5526;
  wire       [35:0]   _zz_5527;
  wire       [35:0]   _zz_5528;
  wire       [35:0]   _zz_5529;
  wire       [26:0]   _zz_5530;
  wire       [35:0]   _zz_5531;
  wire       [17:0]   _zz_5532;
  wire       [35:0]   _zz_5533;
  wire       [35:0]   _zz_5534;
  wire       [35:0]   _zz_5535;
  wire       [35:0]   _zz_5536;
  wire       [35:0]   _zz_5537;
  wire       [26:0]   _zz_5538;
  wire       [35:0]   _zz_5539;
  wire       [17:0]   _zz_5540;
  wire       [35:0]   _zz_5541;
  wire       [35:0]   _zz_5542;
  wire       [35:0]   _zz_5543;
  wire       [35:0]   _zz_5544;
  wire       [35:0]   _zz_5545;
  wire       [26:0]   _zz_5546;
  wire       [35:0]   _zz_5547;
  wire       [17:0]   _zz_5548;
  wire       [35:0]   _zz_5549;
  wire       [35:0]   _zz_5550;
  wire       [35:0]   _zz_5551;
  wire       [35:0]   _zz_5552;
  wire       [35:0]   _zz_5553;
  wire       [26:0]   _zz_5554;
  wire       [35:0]   _zz_5555;
  wire       [17:0]   _zz_5556;
  wire       [17:0]   _zz_5557;
  wire       [35:0]   _zz_5558;
  wire       [35:0]   _zz_5559;
  wire       [17:0]   _zz_5560;
  wire       [35:0]   _zz_5561;
  wire       [35:0]   _zz_5562;
  wire       [35:0]   _zz_5563;
  wire       [17:0]   _zz_5564;
  wire       [35:0]   _zz_5565;
  wire       [35:0]   _zz_5566;
  wire       [35:0]   _zz_5567;
  wire       [35:0]   _zz_5568;
  wire       [35:0]   _zz_5569;
  wire       [35:0]   _zz_5570;
  wire       [26:0]   _zz_5571;
  wire       [35:0]   _zz_5572;
  wire       [17:0]   _zz_5573;
  wire       [35:0]   _zz_5574;
  wire       [35:0]   _zz_5575;
  wire       [35:0]   _zz_5576;
  wire       [35:0]   _zz_5577;
  wire       [35:0]   _zz_5578;
  wire       [26:0]   _zz_5579;
  wire       [35:0]   _zz_5580;
  wire       [17:0]   _zz_5581;
  wire       [35:0]   _zz_5582;
  wire       [35:0]   _zz_5583;
  wire       [35:0]   _zz_5584;
  wire       [35:0]   _zz_5585;
  wire       [35:0]   _zz_5586;
  wire       [26:0]   _zz_5587;
  wire       [35:0]   _zz_5588;
  wire       [17:0]   _zz_5589;
  wire       [35:0]   _zz_5590;
  wire       [35:0]   _zz_5591;
  wire       [35:0]   _zz_5592;
  wire       [35:0]   _zz_5593;
  wire       [35:0]   _zz_5594;
  wire       [26:0]   _zz_5595;
  wire       [35:0]   _zz_5596;
  wire       [17:0]   _zz_5597;
  wire       [17:0]   _zz_5598;
  wire       [35:0]   _zz_5599;
  wire       [35:0]   _zz_5600;
  wire       [17:0]   _zz_5601;
  wire       [35:0]   _zz_5602;
  wire       [35:0]   _zz_5603;
  wire       [35:0]   _zz_5604;
  wire       [17:0]   _zz_5605;
  wire       [35:0]   _zz_5606;
  wire       [35:0]   _zz_5607;
  wire       [35:0]   _zz_5608;
  wire       [35:0]   _zz_5609;
  wire       [35:0]   _zz_5610;
  wire       [35:0]   _zz_5611;
  wire       [26:0]   _zz_5612;
  wire       [35:0]   _zz_5613;
  wire       [17:0]   _zz_5614;
  wire       [35:0]   _zz_5615;
  wire       [35:0]   _zz_5616;
  wire       [35:0]   _zz_5617;
  wire       [35:0]   _zz_5618;
  wire       [35:0]   _zz_5619;
  wire       [26:0]   _zz_5620;
  wire       [35:0]   _zz_5621;
  wire       [17:0]   _zz_5622;
  wire       [35:0]   _zz_5623;
  wire       [35:0]   _zz_5624;
  wire       [35:0]   _zz_5625;
  wire       [35:0]   _zz_5626;
  wire       [35:0]   _zz_5627;
  wire       [26:0]   _zz_5628;
  wire       [35:0]   _zz_5629;
  wire       [17:0]   _zz_5630;
  wire       [35:0]   _zz_5631;
  wire       [35:0]   _zz_5632;
  wire       [35:0]   _zz_5633;
  wire       [35:0]   _zz_5634;
  wire       [35:0]   _zz_5635;
  wire       [26:0]   _zz_5636;
  wire       [35:0]   _zz_5637;
  wire       [17:0]   _zz_5638;
  wire       [17:0]   _zz_5639;
  wire       [35:0]   _zz_5640;
  wire       [35:0]   _zz_5641;
  wire       [17:0]   _zz_5642;
  wire       [35:0]   _zz_5643;
  wire       [35:0]   _zz_5644;
  wire       [35:0]   _zz_5645;
  wire       [17:0]   _zz_5646;
  wire       [35:0]   _zz_5647;
  wire       [35:0]   _zz_5648;
  wire       [35:0]   _zz_5649;
  wire       [35:0]   _zz_5650;
  wire       [35:0]   _zz_5651;
  wire       [35:0]   _zz_5652;
  wire       [26:0]   _zz_5653;
  wire       [35:0]   _zz_5654;
  wire       [17:0]   _zz_5655;
  wire       [35:0]   _zz_5656;
  wire       [35:0]   _zz_5657;
  wire       [35:0]   _zz_5658;
  wire       [35:0]   _zz_5659;
  wire       [35:0]   _zz_5660;
  wire       [26:0]   _zz_5661;
  wire       [35:0]   _zz_5662;
  wire       [17:0]   _zz_5663;
  wire       [35:0]   _zz_5664;
  wire       [35:0]   _zz_5665;
  wire       [35:0]   _zz_5666;
  wire       [35:0]   _zz_5667;
  wire       [35:0]   _zz_5668;
  wire       [26:0]   _zz_5669;
  wire       [35:0]   _zz_5670;
  wire       [17:0]   _zz_5671;
  wire       [35:0]   _zz_5672;
  wire       [35:0]   _zz_5673;
  wire       [35:0]   _zz_5674;
  wire       [35:0]   _zz_5675;
  wire       [35:0]   _zz_5676;
  wire       [26:0]   _zz_5677;
  wire       [35:0]   _zz_5678;
  wire       [17:0]   _zz_5679;
  wire       [17:0]   _zz_5680;
  wire       [35:0]   _zz_5681;
  wire       [35:0]   _zz_5682;
  wire       [17:0]   _zz_5683;
  wire       [35:0]   _zz_5684;
  wire       [35:0]   _zz_5685;
  wire       [35:0]   _zz_5686;
  wire       [17:0]   _zz_5687;
  wire       [35:0]   _zz_5688;
  wire       [35:0]   _zz_5689;
  wire       [35:0]   _zz_5690;
  wire       [35:0]   _zz_5691;
  wire       [35:0]   _zz_5692;
  wire       [35:0]   _zz_5693;
  wire       [26:0]   _zz_5694;
  wire       [35:0]   _zz_5695;
  wire       [17:0]   _zz_5696;
  wire       [35:0]   _zz_5697;
  wire       [35:0]   _zz_5698;
  wire       [35:0]   _zz_5699;
  wire       [35:0]   _zz_5700;
  wire       [35:0]   _zz_5701;
  wire       [26:0]   _zz_5702;
  wire       [35:0]   _zz_5703;
  wire       [17:0]   _zz_5704;
  wire       [35:0]   _zz_5705;
  wire       [35:0]   _zz_5706;
  wire       [35:0]   _zz_5707;
  wire       [35:0]   _zz_5708;
  wire       [35:0]   _zz_5709;
  wire       [26:0]   _zz_5710;
  wire       [35:0]   _zz_5711;
  wire       [17:0]   _zz_5712;
  wire       [35:0]   _zz_5713;
  wire       [35:0]   _zz_5714;
  wire       [35:0]   _zz_5715;
  wire       [35:0]   _zz_5716;
  wire       [35:0]   _zz_5717;
  wire       [26:0]   _zz_5718;
  wire       [35:0]   _zz_5719;
  wire       [17:0]   _zz_5720;
  wire       [17:0]   _zz_5721;
  wire       [35:0]   _zz_5722;
  wire       [35:0]   _zz_5723;
  wire       [17:0]   _zz_5724;
  wire       [35:0]   _zz_5725;
  wire       [35:0]   _zz_5726;
  wire       [35:0]   _zz_5727;
  wire       [17:0]   _zz_5728;
  wire       [35:0]   _zz_5729;
  wire       [35:0]   _zz_5730;
  wire       [35:0]   _zz_5731;
  wire       [35:0]   _zz_5732;
  wire       [35:0]   _zz_5733;
  wire       [35:0]   _zz_5734;
  wire       [26:0]   _zz_5735;
  wire       [35:0]   _zz_5736;
  wire       [17:0]   _zz_5737;
  wire       [35:0]   _zz_5738;
  wire       [35:0]   _zz_5739;
  wire       [35:0]   _zz_5740;
  wire       [35:0]   _zz_5741;
  wire       [35:0]   _zz_5742;
  wire       [26:0]   _zz_5743;
  wire       [35:0]   _zz_5744;
  wire       [17:0]   _zz_5745;
  wire       [35:0]   _zz_5746;
  wire       [35:0]   _zz_5747;
  wire       [35:0]   _zz_5748;
  wire       [35:0]   _zz_5749;
  wire       [35:0]   _zz_5750;
  wire       [26:0]   _zz_5751;
  wire       [35:0]   _zz_5752;
  wire       [17:0]   _zz_5753;
  wire       [35:0]   _zz_5754;
  wire       [35:0]   _zz_5755;
  wire       [35:0]   _zz_5756;
  wire       [35:0]   _zz_5757;
  wire       [35:0]   _zz_5758;
  wire       [26:0]   _zz_5759;
  wire       [35:0]   _zz_5760;
  wire       [17:0]   _zz_5761;
  wire       [17:0]   _zz_5762;
  wire       [35:0]   _zz_5763;
  wire       [35:0]   _zz_5764;
  wire       [17:0]   _zz_5765;
  wire       [35:0]   _zz_5766;
  wire       [35:0]   _zz_5767;
  wire       [35:0]   _zz_5768;
  wire       [17:0]   _zz_5769;
  wire       [35:0]   _zz_5770;
  wire       [35:0]   _zz_5771;
  wire       [35:0]   _zz_5772;
  wire       [35:0]   _zz_5773;
  wire       [35:0]   _zz_5774;
  wire       [35:0]   _zz_5775;
  wire       [26:0]   _zz_5776;
  wire       [35:0]   _zz_5777;
  wire       [17:0]   _zz_5778;
  wire       [35:0]   _zz_5779;
  wire       [35:0]   _zz_5780;
  wire       [35:0]   _zz_5781;
  wire       [35:0]   _zz_5782;
  wire       [35:0]   _zz_5783;
  wire       [26:0]   _zz_5784;
  wire       [35:0]   _zz_5785;
  wire       [17:0]   _zz_5786;
  wire       [35:0]   _zz_5787;
  wire       [35:0]   _zz_5788;
  wire       [35:0]   _zz_5789;
  wire       [35:0]   _zz_5790;
  wire       [35:0]   _zz_5791;
  wire       [26:0]   _zz_5792;
  wire       [35:0]   _zz_5793;
  wire       [17:0]   _zz_5794;
  wire       [35:0]   _zz_5795;
  wire       [35:0]   _zz_5796;
  wire       [35:0]   _zz_5797;
  wire       [35:0]   _zz_5798;
  wire       [35:0]   _zz_5799;
  wire       [26:0]   _zz_5800;
  wire       [35:0]   _zz_5801;
  wire       [17:0]   _zz_5802;
  wire       [17:0]   _zz_5803;
  wire       [35:0]   _zz_5804;
  wire       [35:0]   _zz_5805;
  wire       [17:0]   _zz_5806;
  wire       [35:0]   _zz_5807;
  wire       [35:0]   _zz_5808;
  wire       [35:0]   _zz_5809;
  wire       [17:0]   _zz_5810;
  wire       [35:0]   _zz_5811;
  wire       [35:0]   _zz_5812;
  wire       [35:0]   _zz_5813;
  wire       [35:0]   _zz_5814;
  wire       [35:0]   _zz_5815;
  wire       [35:0]   _zz_5816;
  wire       [26:0]   _zz_5817;
  wire       [35:0]   _zz_5818;
  wire       [17:0]   _zz_5819;
  wire       [35:0]   _zz_5820;
  wire       [35:0]   _zz_5821;
  wire       [35:0]   _zz_5822;
  wire       [35:0]   _zz_5823;
  wire       [35:0]   _zz_5824;
  wire       [26:0]   _zz_5825;
  wire       [35:0]   _zz_5826;
  wire       [17:0]   _zz_5827;
  wire       [35:0]   _zz_5828;
  wire       [35:0]   _zz_5829;
  wire       [35:0]   _zz_5830;
  wire       [35:0]   _zz_5831;
  wire       [35:0]   _zz_5832;
  wire       [26:0]   _zz_5833;
  wire       [35:0]   _zz_5834;
  wire       [17:0]   _zz_5835;
  wire       [35:0]   _zz_5836;
  wire       [35:0]   _zz_5837;
  wire       [35:0]   _zz_5838;
  wire       [35:0]   _zz_5839;
  wire       [35:0]   _zz_5840;
  wire       [26:0]   _zz_5841;
  wire       [35:0]   _zz_5842;
  wire       [17:0]   _zz_5843;
  wire       [17:0]   _zz_5844;
  wire       [35:0]   _zz_5845;
  wire       [35:0]   _zz_5846;
  wire       [17:0]   _zz_5847;
  wire       [35:0]   _zz_5848;
  wire       [35:0]   _zz_5849;
  wire       [35:0]   _zz_5850;
  wire       [17:0]   _zz_5851;
  wire       [35:0]   _zz_5852;
  wire       [35:0]   _zz_5853;
  wire       [35:0]   _zz_5854;
  wire       [35:0]   _zz_5855;
  wire       [35:0]   _zz_5856;
  wire       [35:0]   _zz_5857;
  wire       [26:0]   _zz_5858;
  wire       [35:0]   _zz_5859;
  wire       [17:0]   _zz_5860;
  wire       [35:0]   _zz_5861;
  wire       [35:0]   _zz_5862;
  wire       [35:0]   _zz_5863;
  wire       [35:0]   _zz_5864;
  wire       [35:0]   _zz_5865;
  wire       [26:0]   _zz_5866;
  wire       [35:0]   _zz_5867;
  wire       [17:0]   _zz_5868;
  wire       [35:0]   _zz_5869;
  wire       [35:0]   _zz_5870;
  wire       [35:0]   _zz_5871;
  wire       [35:0]   _zz_5872;
  wire       [35:0]   _zz_5873;
  wire       [26:0]   _zz_5874;
  wire       [35:0]   _zz_5875;
  wire       [17:0]   _zz_5876;
  wire       [35:0]   _zz_5877;
  wire       [35:0]   _zz_5878;
  wire       [35:0]   _zz_5879;
  wire       [35:0]   _zz_5880;
  wire       [35:0]   _zz_5881;
  wire       [26:0]   _zz_5882;
  wire       [35:0]   _zz_5883;
  wire       [17:0]   _zz_5884;
  wire       [17:0]   _zz_5885;
  wire       [35:0]   _zz_5886;
  wire       [35:0]   _zz_5887;
  wire       [17:0]   _zz_5888;
  wire       [35:0]   _zz_5889;
  wire       [35:0]   _zz_5890;
  wire       [35:0]   _zz_5891;
  wire       [17:0]   _zz_5892;
  wire       [35:0]   _zz_5893;
  wire       [35:0]   _zz_5894;
  wire       [35:0]   _zz_5895;
  wire       [35:0]   _zz_5896;
  wire       [35:0]   _zz_5897;
  wire       [35:0]   _zz_5898;
  wire       [26:0]   _zz_5899;
  wire       [35:0]   _zz_5900;
  wire       [17:0]   _zz_5901;
  wire       [35:0]   _zz_5902;
  wire       [35:0]   _zz_5903;
  wire       [35:0]   _zz_5904;
  wire       [35:0]   _zz_5905;
  wire       [35:0]   _zz_5906;
  wire       [26:0]   _zz_5907;
  wire       [35:0]   _zz_5908;
  wire       [17:0]   _zz_5909;
  wire       [35:0]   _zz_5910;
  wire       [35:0]   _zz_5911;
  wire       [35:0]   _zz_5912;
  wire       [35:0]   _zz_5913;
  wire       [35:0]   _zz_5914;
  wire       [26:0]   _zz_5915;
  wire       [35:0]   _zz_5916;
  wire       [17:0]   _zz_5917;
  wire       [35:0]   _zz_5918;
  wire       [35:0]   _zz_5919;
  wire       [35:0]   _zz_5920;
  wire       [35:0]   _zz_5921;
  wire       [35:0]   _zz_5922;
  wire       [26:0]   _zz_5923;
  wire       [35:0]   _zz_5924;
  wire       [17:0]   _zz_5925;
  wire       [17:0]   _zz_5926;
  wire       [35:0]   _zz_5927;
  wire       [35:0]   _zz_5928;
  wire       [17:0]   _zz_5929;
  wire       [35:0]   _zz_5930;
  wire       [35:0]   _zz_5931;
  wire       [35:0]   _zz_5932;
  wire       [17:0]   _zz_5933;
  wire       [35:0]   _zz_5934;
  wire       [35:0]   _zz_5935;
  wire       [35:0]   _zz_5936;
  wire       [35:0]   _zz_5937;
  wire       [35:0]   _zz_5938;
  wire       [35:0]   _zz_5939;
  wire       [26:0]   _zz_5940;
  wire       [35:0]   _zz_5941;
  wire       [17:0]   _zz_5942;
  wire       [35:0]   _zz_5943;
  wire       [35:0]   _zz_5944;
  wire       [35:0]   _zz_5945;
  wire       [35:0]   _zz_5946;
  wire       [35:0]   _zz_5947;
  wire       [26:0]   _zz_5948;
  wire       [35:0]   _zz_5949;
  wire       [17:0]   _zz_5950;
  wire       [35:0]   _zz_5951;
  wire       [35:0]   _zz_5952;
  wire       [35:0]   _zz_5953;
  wire       [35:0]   _zz_5954;
  wire       [35:0]   _zz_5955;
  wire       [26:0]   _zz_5956;
  wire       [35:0]   _zz_5957;
  wire       [17:0]   _zz_5958;
  wire       [35:0]   _zz_5959;
  wire       [35:0]   _zz_5960;
  wire       [35:0]   _zz_5961;
  wire       [35:0]   _zz_5962;
  wire       [35:0]   _zz_5963;
  wire       [26:0]   _zz_5964;
  wire       [35:0]   _zz_5965;
  wire       [17:0]   _zz_5966;
  wire       [17:0]   _zz_5967;
  wire       [35:0]   _zz_5968;
  wire       [35:0]   _zz_5969;
  wire       [17:0]   _zz_5970;
  wire       [35:0]   _zz_5971;
  wire       [35:0]   _zz_5972;
  wire       [35:0]   _zz_5973;
  wire       [17:0]   _zz_5974;
  wire       [35:0]   _zz_5975;
  wire       [35:0]   _zz_5976;
  wire       [35:0]   _zz_5977;
  wire       [35:0]   _zz_5978;
  wire       [35:0]   _zz_5979;
  wire       [35:0]   _zz_5980;
  wire       [26:0]   _zz_5981;
  wire       [35:0]   _zz_5982;
  wire       [17:0]   _zz_5983;
  wire       [35:0]   _zz_5984;
  wire       [35:0]   _zz_5985;
  wire       [35:0]   _zz_5986;
  wire       [35:0]   _zz_5987;
  wire       [35:0]   _zz_5988;
  wire       [26:0]   _zz_5989;
  wire       [35:0]   _zz_5990;
  wire       [17:0]   _zz_5991;
  wire       [35:0]   _zz_5992;
  wire       [35:0]   _zz_5993;
  wire       [35:0]   _zz_5994;
  wire       [35:0]   _zz_5995;
  wire       [35:0]   _zz_5996;
  wire       [26:0]   _zz_5997;
  wire       [35:0]   _zz_5998;
  wire       [17:0]   _zz_5999;
  wire       [35:0]   _zz_6000;
  wire       [35:0]   _zz_6001;
  wire       [35:0]   _zz_6002;
  wire       [35:0]   _zz_6003;
  wire       [35:0]   _zz_6004;
  wire       [26:0]   _zz_6005;
  wire       [35:0]   _zz_6006;
  wire       [17:0]   _zz_6007;
  wire       [17:0]   _zz_6008;
  wire       [35:0]   _zz_6009;
  wire       [35:0]   _zz_6010;
  wire       [17:0]   _zz_6011;
  wire       [35:0]   _zz_6012;
  wire       [35:0]   _zz_6013;
  wire       [35:0]   _zz_6014;
  wire       [17:0]   _zz_6015;
  wire       [35:0]   _zz_6016;
  wire       [35:0]   _zz_6017;
  wire       [35:0]   _zz_6018;
  wire       [35:0]   _zz_6019;
  wire       [35:0]   _zz_6020;
  wire       [35:0]   _zz_6021;
  wire       [26:0]   _zz_6022;
  wire       [35:0]   _zz_6023;
  wire       [17:0]   _zz_6024;
  wire       [35:0]   _zz_6025;
  wire       [35:0]   _zz_6026;
  wire       [35:0]   _zz_6027;
  wire       [35:0]   _zz_6028;
  wire       [35:0]   _zz_6029;
  wire       [26:0]   _zz_6030;
  wire       [35:0]   _zz_6031;
  wire       [17:0]   _zz_6032;
  wire       [35:0]   _zz_6033;
  wire       [35:0]   _zz_6034;
  wire       [35:0]   _zz_6035;
  wire       [35:0]   _zz_6036;
  wire       [35:0]   _zz_6037;
  wire       [26:0]   _zz_6038;
  wire       [35:0]   _zz_6039;
  wire       [17:0]   _zz_6040;
  wire       [35:0]   _zz_6041;
  wire       [35:0]   _zz_6042;
  wire       [35:0]   _zz_6043;
  wire       [35:0]   _zz_6044;
  wire       [35:0]   _zz_6045;
  wire       [26:0]   _zz_6046;
  wire       [35:0]   _zz_6047;
  wire       [17:0]   _zz_6048;
  wire       [17:0]   _zz_6049;
  wire       [35:0]   _zz_6050;
  wire       [35:0]   _zz_6051;
  wire       [17:0]   _zz_6052;
  wire       [35:0]   _zz_6053;
  wire       [35:0]   _zz_6054;
  wire       [35:0]   _zz_6055;
  wire       [17:0]   _zz_6056;
  wire       [35:0]   _zz_6057;
  wire       [35:0]   _zz_6058;
  wire       [35:0]   _zz_6059;
  wire       [35:0]   _zz_6060;
  wire       [35:0]   _zz_6061;
  wire       [35:0]   _zz_6062;
  wire       [26:0]   _zz_6063;
  wire       [35:0]   _zz_6064;
  wire       [17:0]   _zz_6065;
  wire       [35:0]   _zz_6066;
  wire       [35:0]   _zz_6067;
  wire       [35:0]   _zz_6068;
  wire       [35:0]   _zz_6069;
  wire       [35:0]   _zz_6070;
  wire       [26:0]   _zz_6071;
  wire       [35:0]   _zz_6072;
  wire       [17:0]   _zz_6073;
  wire       [35:0]   _zz_6074;
  wire       [35:0]   _zz_6075;
  wire       [35:0]   _zz_6076;
  wire       [35:0]   _zz_6077;
  wire       [35:0]   _zz_6078;
  wire       [26:0]   _zz_6079;
  wire       [35:0]   _zz_6080;
  wire       [17:0]   _zz_6081;
  wire       [35:0]   _zz_6082;
  wire       [35:0]   _zz_6083;
  wire       [35:0]   _zz_6084;
  wire       [35:0]   _zz_6085;
  wire       [35:0]   _zz_6086;
  wire       [26:0]   _zz_6087;
  wire       [35:0]   _zz_6088;
  wire       [17:0]   _zz_6089;
  wire       [17:0]   _zz_6090;
  wire       [35:0]   _zz_6091;
  wire       [35:0]   _zz_6092;
  wire       [17:0]   _zz_6093;
  wire       [35:0]   _zz_6094;
  wire       [35:0]   _zz_6095;
  wire       [35:0]   _zz_6096;
  wire       [17:0]   _zz_6097;
  wire       [35:0]   _zz_6098;
  wire       [35:0]   _zz_6099;
  wire       [35:0]   _zz_6100;
  wire       [35:0]   _zz_6101;
  wire       [35:0]   _zz_6102;
  wire       [35:0]   _zz_6103;
  wire       [26:0]   _zz_6104;
  wire       [35:0]   _zz_6105;
  wire       [17:0]   _zz_6106;
  wire       [35:0]   _zz_6107;
  wire       [35:0]   _zz_6108;
  wire       [35:0]   _zz_6109;
  wire       [35:0]   _zz_6110;
  wire       [35:0]   _zz_6111;
  wire       [26:0]   _zz_6112;
  wire       [35:0]   _zz_6113;
  wire       [17:0]   _zz_6114;
  wire       [35:0]   _zz_6115;
  wire       [35:0]   _zz_6116;
  wire       [35:0]   _zz_6117;
  wire       [35:0]   _zz_6118;
  wire       [35:0]   _zz_6119;
  wire       [26:0]   _zz_6120;
  wire       [35:0]   _zz_6121;
  wire       [17:0]   _zz_6122;
  wire       [35:0]   _zz_6123;
  wire       [35:0]   _zz_6124;
  wire       [35:0]   _zz_6125;
  wire       [35:0]   _zz_6126;
  wire       [35:0]   _zz_6127;
  wire       [26:0]   _zz_6128;
  wire       [35:0]   _zz_6129;
  wire       [17:0]   _zz_6130;
  wire       [17:0]   _zz_6131;
  wire       [35:0]   _zz_6132;
  wire       [35:0]   _zz_6133;
  wire       [17:0]   _zz_6134;
  wire       [35:0]   _zz_6135;
  wire       [35:0]   _zz_6136;
  wire       [35:0]   _zz_6137;
  wire       [17:0]   _zz_6138;
  wire       [35:0]   _zz_6139;
  wire       [35:0]   _zz_6140;
  wire       [35:0]   _zz_6141;
  wire       [35:0]   _zz_6142;
  wire       [35:0]   _zz_6143;
  wire       [35:0]   _zz_6144;
  wire       [26:0]   _zz_6145;
  wire       [35:0]   _zz_6146;
  wire       [17:0]   _zz_6147;
  wire       [35:0]   _zz_6148;
  wire       [35:0]   _zz_6149;
  wire       [35:0]   _zz_6150;
  wire       [35:0]   _zz_6151;
  wire       [35:0]   _zz_6152;
  wire       [26:0]   _zz_6153;
  wire       [35:0]   _zz_6154;
  wire       [17:0]   _zz_6155;
  wire       [35:0]   _zz_6156;
  wire       [35:0]   _zz_6157;
  wire       [35:0]   _zz_6158;
  wire       [35:0]   _zz_6159;
  wire       [35:0]   _zz_6160;
  wire       [26:0]   _zz_6161;
  wire       [35:0]   _zz_6162;
  wire       [17:0]   _zz_6163;
  wire       [35:0]   _zz_6164;
  wire       [35:0]   _zz_6165;
  wire       [35:0]   _zz_6166;
  wire       [35:0]   _zz_6167;
  wire       [35:0]   _zz_6168;
  wire       [26:0]   _zz_6169;
  wire       [35:0]   _zz_6170;
  wire       [17:0]   _zz_6171;
  wire       [17:0]   _zz_6172;
  wire       [35:0]   _zz_6173;
  wire       [35:0]   _zz_6174;
  wire       [17:0]   _zz_6175;
  wire       [35:0]   _zz_6176;
  wire       [35:0]   _zz_6177;
  wire       [35:0]   _zz_6178;
  wire       [17:0]   _zz_6179;
  wire       [35:0]   _zz_6180;
  wire       [35:0]   _zz_6181;
  wire       [35:0]   _zz_6182;
  wire       [35:0]   _zz_6183;
  wire       [35:0]   _zz_6184;
  wire       [35:0]   _zz_6185;
  wire       [26:0]   _zz_6186;
  wire       [35:0]   _zz_6187;
  wire       [17:0]   _zz_6188;
  wire       [35:0]   _zz_6189;
  wire       [35:0]   _zz_6190;
  wire       [35:0]   _zz_6191;
  wire       [35:0]   _zz_6192;
  wire       [35:0]   _zz_6193;
  wire       [26:0]   _zz_6194;
  wire       [35:0]   _zz_6195;
  wire       [17:0]   _zz_6196;
  wire       [35:0]   _zz_6197;
  wire       [35:0]   _zz_6198;
  wire       [35:0]   _zz_6199;
  wire       [35:0]   _zz_6200;
  wire       [35:0]   _zz_6201;
  wire       [26:0]   _zz_6202;
  wire       [35:0]   _zz_6203;
  wire       [17:0]   _zz_6204;
  wire       [35:0]   _zz_6205;
  wire       [35:0]   _zz_6206;
  wire       [35:0]   _zz_6207;
  wire       [35:0]   _zz_6208;
  wire       [35:0]   _zz_6209;
  wire       [26:0]   _zz_6210;
  wire       [35:0]   _zz_6211;
  wire       [17:0]   _zz_6212;
  wire       [17:0]   _zz_6213;
  wire       [35:0]   _zz_6214;
  wire       [35:0]   _zz_6215;
  wire       [17:0]   _zz_6216;
  wire       [35:0]   _zz_6217;
  wire       [35:0]   _zz_6218;
  wire       [35:0]   _zz_6219;
  wire       [17:0]   _zz_6220;
  wire       [35:0]   _zz_6221;
  wire       [35:0]   _zz_6222;
  wire       [35:0]   _zz_6223;
  wire       [35:0]   _zz_6224;
  wire       [35:0]   _zz_6225;
  wire       [35:0]   _zz_6226;
  wire       [26:0]   _zz_6227;
  wire       [35:0]   _zz_6228;
  wire       [17:0]   _zz_6229;
  wire       [35:0]   _zz_6230;
  wire       [35:0]   _zz_6231;
  wire       [35:0]   _zz_6232;
  wire       [35:0]   _zz_6233;
  wire       [35:0]   _zz_6234;
  wire       [26:0]   _zz_6235;
  wire       [35:0]   _zz_6236;
  wire       [17:0]   _zz_6237;
  wire       [35:0]   _zz_6238;
  wire       [35:0]   _zz_6239;
  wire       [35:0]   _zz_6240;
  wire       [35:0]   _zz_6241;
  wire       [35:0]   _zz_6242;
  wire       [26:0]   _zz_6243;
  wire       [35:0]   _zz_6244;
  wire       [17:0]   _zz_6245;
  wire       [35:0]   _zz_6246;
  wire       [35:0]   _zz_6247;
  wire       [35:0]   _zz_6248;
  wire       [35:0]   _zz_6249;
  wire       [35:0]   _zz_6250;
  wire       [26:0]   _zz_6251;
  wire       [35:0]   _zz_6252;
  wire       [17:0]   _zz_6253;
  wire       [17:0]   _zz_6254;
  wire       [35:0]   _zz_6255;
  wire       [35:0]   _zz_6256;
  wire       [17:0]   _zz_6257;
  wire       [35:0]   _zz_6258;
  wire       [35:0]   _zz_6259;
  wire       [35:0]   _zz_6260;
  wire       [17:0]   _zz_6261;
  wire       [35:0]   _zz_6262;
  wire       [35:0]   _zz_6263;
  wire       [35:0]   _zz_6264;
  wire       [35:0]   _zz_6265;
  wire       [35:0]   _zz_6266;
  wire       [35:0]   _zz_6267;
  wire       [26:0]   _zz_6268;
  wire       [35:0]   _zz_6269;
  wire       [17:0]   _zz_6270;
  wire       [35:0]   _zz_6271;
  wire       [35:0]   _zz_6272;
  wire       [35:0]   _zz_6273;
  wire       [35:0]   _zz_6274;
  wire       [35:0]   _zz_6275;
  wire       [26:0]   _zz_6276;
  wire       [35:0]   _zz_6277;
  wire       [17:0]   _zz_6278;
  wire       [35:0]   _zz_6279;
  wire       [35:0]   _zz_6280;
  wire       [35:0]   _zz_6281;
  wire       [35:0]   _zz_6282;
  wire       [35:0]   _zz_6283;
  wire       [26:0]   _zz_6284;
  wire       [35:0]   _zz_6285;
  wire       [17:0]   _zz_6286;
  wire       [35:0]   _zz_6287;
  wire       [35:0]   _zz_6288;
  wire       [35:0]   _zz_6289;
  wire       [35:0]   _zz_6290;
  wire       [35:0]   _zz_6291;
  wire       [26:0]   _zz_6292;
  wire       [35:0]   _zz_6293;
  wire       [17:0]   _zz_6294;
  wire       [17:0]   _zz_6295;
  wire       [35:0]   _zz_6296;
  wire       [35:0]   _zz_6297;
  wire       [17:0]   _zz_6298;
  wire       [35:0]   _zz_6299;
  wire       [35:0]   _zz_6300;
  wire       [35:0]   _zz_6301;
  wire       [17:0]   _zz_6302;
  wire       [35:0]   _zz_6303;
  wire       [35:0]   _zz_6304;
  wire       [35:0]   _zz_6305;
  wire       [35:0]   _zz_6306;
  wire       [35:0]   _zz_6307;
  wire       [35:0]   _zz_6308;
  wire       [26:0]   _zz_6309;
  wire       [35:0]   _zz_6310;
  wire       [17:0]   _zz_6311;
  wire       [35:0]   _zz_6312;
  wire       [35:0]   _zz_6313;
  wire       [35:0]   _zz_6314;
  wire       [35:0]   _zz_6315;
  wire       [35:0]   _zz_6316;
  wire       [26:0]   _zz_6317;
  wire       [35:0]   _zz_6318;
  wire       [17:0]   _zz_6319;
  wire       [35:0]   _zz_6320;
  wire       [35:0]   _zz_6321;
  wire       [35:0]   _zz_6322;
  wire       [35:0]   _zz_6323;
  wire       [35:0]   _zz_6324;
  wire       [26:0]   _zz_6325;
  wire       [35:0]   _zz_6326;
  wire       [17:0]   _zz_6327;
  wire       [35:0]   _zz_6328;
  wire       [35:0]   _zz_6329;
  wire       [35:0]   _zz_6330;
  wire       [35:0]   _zz_6331;
  wire       [35:0]   _zz_6332;
  wire       [26:0]   _zz_6333;
  wire       [35:0]   _zz_6334;
  wire       [17:0]   _zz_6335;
  wire       [17:0]   _zz_6336;
  wire       [35:0]   _zz_6337;
  wire       [35:0]   _zz_6338;
  wire       [17:0]   _zz_6339;
  wire       [35:0]   _zz_6340;
  wire       [35:0]   _zz_6341;
  wire       [35:0]   _zz_6342;
  wire       [17:0]   _zz_6343;
  wire       [35:0]   _zz_6344;
  wire       [35:0]   _zz_6345;
  wire       [35:0]   _zz_6346;
  wire       [35:0]   _zz_6347;
  wire       [35:0]   _zz_6348;
  wire       [35:0]   _zz_6349;
  wire       [26:0]   _zz_6350;
  wire       [35:0]   _zz_6351;
  wire       [17:0]   _zz_6352;
  wire       [35:0]   _zz_6353;
  wire       [35:0]   _zz_6354;
  wire       [35:0]   _zz_6355;
  wire       [35:0]   _zz_6356;
  wire       [35:0]   _zz_6357;
  wire       [26:0]   _zz_6358;
  wire       [35:0]   _zz_6359;
  wire       [17:0]   _zz_6360;
  wire       [35:0]   _zz_6361;
  wire       [35:0]   _zz_6362;
  wire       [35:0]   _zz_6363;
  wire       [35:0]   _zz_6364;
  wire       [35:0]   _zz_6365;
  wire       [26:0]   _zz_6366;
  wire       [35:0]   _zz_6367;
  wire       [17:0]   _zz_6368;
  wire       [35:0]   _zz_6369;
  wire       [35:0]   _zz_6370;
  wire       [35:0]   _zz_6371;
  wire       [35:0]   _zz_6372;
  wire       [35:0]   _zz_6373;
  wire       [26:0]   _zz_6374;
  wire       [35:0]   _zz_6375;
  wire       [17:0]   _zz_6376;
  wire       [17:0]   _zz_6377;
  wire       [35:0]   _zz_6378;
  wire       [35:0]   _zz_6379;
  wire       [17:0]   _zz_6380;
  wire       [35:0]   _zz_6381;
  wire       [35:0]   _zz_6382;
  wire       [35:0]   _zz_6383;
  wire       [17:0]   _zz_6384;
  wire       [35:0]   _zz_6385;
  wire       [35:0]   _zz_6386;
  wire       [35:0]   _zz_6387;
  wire       [35:0]   _zz_6388;
  wire       [35:0]   _zz_6389;
  wire       [35:0]   _zz_6390;
  wire       [26:0]   _zz_6391;
  wire       [35:0]   _zz_6392;
  wire       [17:0]   _zz_6393;
  wire       [35:0]   _zz_6394;
  wire       [35:0]   _zz_6395;
  wire       [35:0]   _zz_6396;
  wire       [35:0]   _zz_6397;
  wire       [35:0]   _zz_6398;
  wire       [26:0]   _zz_6399;
  wire       [35:0]   _zz_6400;
  wire       [17:0]   _zz_6401;
  wire       [35:0]   _zz_6402;
  wire       [35:0]   _zz_6403;
  wire       [35:0]   _zz_6404;
  wire       [35:0]   _zz_6405;
  wire       [35:0]   _zz_6406;
  wire       [26:0]   _zz_6407;
  wire       [35:0]   _zz_6408;
  wire       [17:0]   _zz_6409;
  wire       [35:0]   _zz_6410;
  wire       [35:0]   _zz_6411;
  wire       [35:0]   _zz_6412;
  wire       [35:0]   _zz_6413;
  wire       [35:0]   _zz_6414;
  wire       [26:0]   _zz_6415;
  wire       [35:0]   _zz_6416;
  wire       [17:0]   _zz_6417;
  wire       [17:0]   _zz_6418;
  wire       [35:0]   _zz_6419;
  wire       [35:0]   _zz_6420;
  wire       [17:0]   _zz_6421;
  wire       [35:0]   _zz_6422;
  wire       [35:0]   _zz_6423;
  wire       [35:0]   _zz_6424;
  wire       [17:0]   _zz_6425;
  wire       [35:0]   _zz_6426;
  wire       [35:0]   _zz_6427;
  wire       [35:0]   _zz_6428;
  wire       [35:0]   _zz_6429;
  wire       [35:0]   _zz_6430;
  wire       [35:0]   _zz_6431;
  wire       [26:0]   _zz_6432;
  wire       [35:0]   _zz_6433;
  wire       [17:0]   _zz_6434;
  wire       [35:0]   _zz_6435;
  wire       [35:0]   _zz_6436;
  wire       [35:0]   _zz_6437;
  wire       [35:0]   _zz_6438;
  wire       [35:0]   _zz_6439;
  wire       [26:0]   _zz_6440;
  wire       [35:0]   _zz_6441;
  wire       [17:0]   _zz_6442;
  wire       [35:0]   _zz_6443;
  wire       [35:0]   _zz_6444;
  wire       [35:0]   _zz_6445;
  wire       [35:0]   _zz_6446;
  wire       [35:0]   _zz_6447;
  wire       [26:0]   _zz_6448;
  wire       [35:0]   _zz_6449;
  wire       [17:0]   _zz_6450;
  wire       [35:0]   _zz_6451;
  wire       [35:0]   _zz_6452;
  wire       [35:0]   _zz_6453;
  wire       [35:0]   _zz_6454;
  wire       [35:0]   _zz_6455;
  wire       [26:0]   _zz_6456;
  wire       [35:0]   _zz_6457;
  wire       [17:0]   _zz_6458;
  wire       [17:0]   _zz_6459;
  wire       [35:0]   _zz_6460;
  wire       [35:0]   _zz_6461;
  wire       [17:0]   _zz_6462;
  wire       [35:0]   _zz_6463;
  wire       [35:0]   _zz_6464;
  wire       [35:0]   _zz_6465;
  wire       [17:0]   _zz_6466;
  wire       [35:0]   _zz_6467;
  wire       [35:0]   _zz_6468;
  wire       [35:0]   _zz_6469;
  wire       [35:0]   _zz_6470;
  wire       [35:0]   _zz_6471;
  wire       [35:0]   _zz_6472;
  wire       [26:0]   _zz_6473;
  wire       [35:0]   _zz_6474;
  wire       [17:0]   _zz_6475;
  wire       [35:0]   _zz_6476;
  wire       [35:0]   _zz_6477;
  wire       [35:0]   _zz_6478;
  wire       [35:0]   _zz_6479;
  wire       [35:0]   _zz_6480;
  wire       [26:0]   _zz_6481;
  wire       [35:0]   _zz_6482;
  wire       [17:0]   _zz_6483;
  wire       [35:0]   _zz_6484;
  wire       [35:0]   _zz_6485;
  wire       [35:0]   _zz_6486;
  wire       [35:0]   _zz_6487;
  wire       [35:0]   _zz_6488;
  wire       [26:0]   _zz_6489;
  wire       [35:0]   _zz_6490;
  wire       [17:0]   _zz_6491;
  wire       [35:0]   _zz_6492;
  wire       [35:0]   _zz_6493;
  wire       [35:0]   _zz_6494;
  wire       [35:0]   _zz_6495;
  wire       [35:0]   _zz_6496;
  wire       [26:0]   _zz_6497;
  wire       [35:0]   _zz_6498;
  wire       [17:0]   _zz_6499;
  wire       [17:0]   _zz_6500;
  wire       [35:0]   _zz_6501;
  wire       [35:0]   _zz_6502;
  wire       [17:0]   _zz_6503;
  wire       [35:0]   _zz_6504;
  wire       [35:0]   _zz_6505;
  wire       [35:0]   _zz_6506;
  wire       [17:0]   _zz_6507;
  wire       [35:0]   _zz_6508;
  wire       [35:0]   _zz_6509;
  wire       [35:0]   _zz_6510;
  wire       [35:0]   _zz_6511;
  wire       [35:0]   _zz_6512;
  wire       [35:0]   _zz_6513;
  wire       [26:0]   _zz_6514;
  wire       [35:0]   _zz_6515;
  wire       [17:0]   _zz_6516;
  wire       [35:0]   _zz_6517;
  wire       [35:0]   _zz_6518;
  wire       [35:0]   _zz_6519;
  wire       [35:0]   _zz_6520;
  wire       [35:0]   _zz_6521;
  wire       [26:0]   _zz_6522;
  wire       [35:0]   _zz_6523;
  wire       [17:0]   _zz_6524;
  wire       [35:0]   _zz_6525;
  wire       [35:0]   _zz_6526;
  wire       [35:0]   _zz_6527;
  wire       [35:0]   _zz_6528;
  wire       [35:0]   _zz_6529;
  wire       [26:0]   _zz_6530;
  wire       [35:0]   _zz_6531;
  wire       [17:0]   _zz_6532;
  wire       [35:0]   _zz_6533;
  wire       [35:0]   _zz_6534;
  wire       [35:0]   _zz_6535;
  wire       [35:0]   _zz_6536;
  wire       [35:0]   _zz_6537;
  wire       [26:0]   _zz_6538;
  wire       [35:0]   _zz_6539;
  wire       [17:0]   _zz_6540;
  wire       [17:0]   _zz_6541;
  wire       [35:0]   _zz_6542;
  wire       [35:0]   _zz_6543;
  wire       [17:0]   _zz_6544;
  wire       [35:0]   _zz_6545;
  wire       [35:0]   _zz_6546;
  wire       [35:0]   _zz_6547;
  wire       [17:0]   _zz_6548;
  wire       [35:0]   _zz_6549;
  wire       [35:0]   _zz_6550;
  wire       [35:0]   _zz_6551;
  wire       [35:0]   _zz_6552;
  wire       [35:0]   _zz_6553;
  wire       [35:0]   _zz_6554;
  wire       [26:0]   _zz_6555;
  wire       [35:0]   _zz_6556;
  wire       [17:0]   _zz_6557;
  wire       [35:0]   _zz_6558;
  wire       [35:0]   _zz_6559;
  wire       [35:0]   _zz_6560;
  wire       [35:0]   _zz_6561;
  wire       [35:0]   _zz_6562;
  wire       [26:0]   _zz_6563;
  wire       [35:0]   _zz_6564;
  wire       [17:0]   _zz_6565;
  wire       [35:0]   _zz_6566;
  wire       [35:0]   _zz_6567;
  wire       [35:0]   _zz_6568;
  wire       [35:0]   _zz_6569;
  wire       [35:0]   _zz_6570;
  wire       [26:0]   _zz_6571;
  wire       [35:0]   _zz_6572;
  wire       [17:0]   _zz_6573;
  wire       [35:0]   _zz_6574;
  wire       [35:0]   _zz_6575;
  wire       [35:0]   _zz_6576;
  wire       [35:0]   _zz_6577;
  wire       [35:0]   _zz_6578;
  wire       [26:0]   _zz_6579;
  wire       [35:0]   _zz_6580;
  wire       [17:0]   _zz_6581;
  wire       [17:0]   _zz_6582;
  wire       [35:0]   _zz_6583;
  wire       [35:0]   _zz_6584;
  wire       [17:0]   _zz_6585;
  wire       [35:0]   _zz_6586;
  wire       [35:0]   _zz_6587;
  wire       [35:0]   _zz_6588;
  wire       [17:0]   _zz_6589;
  wire       [35:0]   _zz_6590;
  wire       [35:0]   _zz_6591;
  wire       [35:0]   _zz_6592;
  wire       [35:0]   _zz_6593;
  wire       [35:0]   _zz_6594;
  wire       [35:0]   _zz_6595;
  wire       [26:0]   _zz_6596;
  wire       [35:0]   _zz_6597;
  wire       [17:0]   _zz_6598;
  wire       [35:0]   _zz_6599;
  wire       [35:0]   _zz_6600;
  wire       [35:0]   _zz_6601;
  wire       [35:0]   _zz_6602;
  wire       [35:0]   _zz_6603;
  wire       [26:0]   _zz_6604;
  wire       [35:0]   _zz_6605;
  wire       [17:0]   _zz_6606;
  wire       [35:0]   _zz_6607;
  wire       [35:0]   _zz_6608;
  wire       [35:0]   _zz_6609;
  wire       [35:0]   _zz_6610;
  wire       [35:0]   _zz_6611;
  wire       [26:0]   _zz_6612;
  wire       [35:0]   _zz_6613;
  wire       [17:0]   _zz_6614;
  wire       [35:0]   _zz_6615;
  wire       [35:0]   _zz_6616;
  wire       [35:0]   _zz_6617;
  wire       [35:0]   _zz_6618;
  wire       [35:0]   _zz_6619;
  wire       [26:0]   _zz_6620;
  wire       [35:0]   _zz_6621;
  wire       [17:0]   _zz_6622;
  wire       [17:0]   _zz_6623;
  wire       [35:0]   _zz_6624;
  wire       [35:0]   _zz_6625;
  wire       [17:0]   _zz_6626;
  wire       [35:0]   _zz_6627;
  wire       [35:0]   _zz_6628;
  wire       [35:0]   _zz_6629;
  wire       [17:0]   _zz_6630;
  wire       [35:0]   _zz_6631;
  wire       [35:0]   _zz_6632;
  wire       [35:0]   _zz_6633;
  wire       [35:0]   _zz_6634;
  wire       [35:0]   _zz_6635;
  wire       [35:0]   _zz_6636;
  wire       [26:0]   _zz_6637;
  wire       [35:0]   _zz_6638;
  wire       [17:0]   _zz_6639;
  wire       [35:0]   _zz_6640;
  wire       [35:0]   _zz_6641;
  wire       [35:0]   _zz_6642;
  wire       [35:0]   _zz_6643;
  wire       [35:0]   _zz_6644;
  wire       [26:0]   _zz_6645;
  wire       [35:0]   _zz_6646;
  wire       [17:0]   _zz_6647;
  wire       [35:0]   _zz_6648;
  wire       [35:0]   _zz_6649;
  wire       [35:0]   _zz_6650;
  wire       [35:0]   _zz_6651;
  wire       [35:0]   _zz_6652;
  wire       [26:0]   _zz_6653;
  wire       [35:0]   _zz_6654;
  wire       [17:0]   _zz_6655;
  wire       [35:0]   _zz_6656;
  wire       [35:0]   _zz_6657;
  wire       [35:0]   _zz_6658;
  wire       [35:0]   _zz_6659;
  wire       [35:0]   _zz_6660;
  wire       [26:0]   _zz_6661;
  wire       [35:0]   _zz_6662;
  wire       [17:0]   _zz_6663;
  wire       [17:0]   _zz_6664;
  wire       [35:0]   _zz_6665;
  wire       [35:0]   _zz_6666;
  wire       [17:0]   _zz_6667;
  wire       [35:0]   _zz_6668;
  wire       [35:0]   _zz_6669;
  wire       [35:0]   _zz_6670;
  wire       [17:0]   _zz_6671;
  wire       [35:0]   _zz_6672;
  wire       [35:0]   _zz_6673;
  wire       [35:0]   _zz_6674;
  wire       [35:0]   _zz_6675;
  wire       [35:0]   _zz_6676;
  wire       [35:0]   _zz_6677;
  wire       [26:0]   _zz_6678;
  wire       [35:0]   _zz_6679;
  wire       [17:0]   _zz_6680;
  wire       [35:0]   _zz_6681;
  wire       [35:0]   _zz_6682;
  wire       [35:0]   _zz_6683;
  wire       [35:0]   _zz_6684;
  wire       [35:0]   _zz_6685;
  wire       [26:0]   _zz_6686;
  wire       [35:0]   _zz_6687;
  wire       [17:0]   _zz_6688;
  wire       [35:0]   _zz_6689;
  wire       [35:0]   _zz_6690;
  wire       [35:0]   _zz_6691;
  wire       [35:0]   _zz_6692;
  wire       [35:0]   _zz_6693;
  wire       [26:0]   _zz_6694;
  wire       [35:0]   _zz_6695;
  wire       [17:0]   _zz_6696;
  wire       [35:0]   _zz_6697;
  wire       [35:0]   _zz_6698;
  wire       [35:0]   _zz_6699;
  wire       [35:0]   _zz_6700;
  wire       [35:0]   _zz_6701;
  wire       [26:0]   _zz_6702;
  wire       [35:0]   _zz_6703;
  wire       [17:0]   _zz_6704;
  wire       [17:0]   _zz_6705;
  wire       [35:0]   _zz_6706;
  wire       [35:0]   _zz_6707;
  wire       [17:0]   _zz_6708;
  wire       [35:0]   _zz_6709;
  wire       [35:0]   _zz_6710;
  wire       [35:0]   _zz_6711;
  wire       [17:0]   _zz_6712;
  wire       [35:0]   _zz_6713;
  wire       [35:0]   _zz_6714;
  wire       [35:0]   _zz_6715;
  wire       [35:0]   _zz_6716;
  wire       [35:0]   _zz_6717;
  wire       [35:0]   _zz_6718;
  wire       [26:0]   _zz_6719;
  wire       [35:0]   _zz_6720;
  wire       [17:0]   _zz_6721;
  wire       [35:0]   _zz_6722;
  wire       [35:0]   _zz_6723;
  wire       [35:0]   _zz_6724;
  wire       [35:0]   _zz_6725;
  wire       [35:0]   _zz_6726;
  wire       [26:0]   _zz_6727;
  wire       [35:0]   _zz_6728;
  wire       [17:0]   _zz_6729;
  wire       [35:0]   _zz_6730;
  wire       [35:0]   _zz_6731;
  wire       [35:0]   _zz_6732;
  wire       [35:0]   _zz_6733;
  wire       [35:0]   _zz_6734;
  wire       [26:0]   _zz_6735;
  wire       [35:0]   _zz_6736;
  wire       [17:0]   _zz_6737;
  wire       [35:0]   _zz_6738;
  wire       [35:0]   _zz_6739;
  wire       [35:0]   _zz_6740;
  wire       [35:0]   _zz_6741;
  wire       [35:0]   _zz_6742;
  wire       [26:0]   _zz_6743;
  wire       [35:0]   _zz_6744;
  wire       [17:0]   _zz_6745;
  wire       [17:0]   _zz_6746;
  wire       [35:0]   _zz_6747;
  wire       [35:0]   _zz_6748;
  wire       [17:0]   _zz_6749;
  wire       [35:0]   _zz_6750;
  wire       [35:0]   _zz_6751;
  wire       [35:0]   _zz_6752;
  wire       [17:0]   _zz_6753;
  wire       [35:0]   _zz_6754;
  wire       [35:0]   _zz_6755;
  wire       [35:0]   _zz_6756;
  wire       [35:0]   _zz_6757;
  wire       [35:0]   _zz_6758;
  wire       [35:0]   _zz_6759;
  wire       [26:0]   _zz_6760;
  wire       [35:0]   _zz_6761;
  wire       [17:0]   _zz_6762;
  wire       [35:0]   _zz_6763;
  wire       [35:0]   _zz_6764;
  wire       [35:0]   _zz_6765;
  wire       [35:0]   _zz_6766;
  wire       [35:0]   _zz_6767;
  wire       [26:0]   _zz_6768;
  wire       [35:0]   _zz_6769;
  wire       [17:0]   _zz_6770;
  wire       [35:0]   _zz_6771;
  wire       [35:0]   _zz_6772;
  wire       [35:0]   _zz_6773;
  wire       [35:0]   _zz_6774;
  wire       [35:0]   _zz_6775;
  wire       [26:0]   _zz_6776;
  wire       [35:0]   _zz_6777;
  wire       [17:0]   _zz_6778;
  wire       [35:0]   _zz_6779;
  wire       [35:0]   _zz_6780;
  wire       [35:0]   _zz_6781;
  wire       [35:0]   _zz_6782;
  wire       [35:0]   _zz_6783;
  wire       [26:0]   _zz_6784;
  wire       [35:0]   _zz_6785;
  wire       [17:0]   _zz_6786;
  wire       [17:0]   _zz_6787;
  wire       [35:0]   _zz_6788;
  wire       [35:0]   _zz_6789;
  wire       [17:0]   _zz_6790;
  wire       [35:0]   _zz_6791;
  wire       [35:0]   _zz_6792;
  wire       [35:0]   _zz_6793;
  wire       [17:0]   _zz_6794;
  wire       [35:0]   _zz_6795;
  wire       [35:0]   _zz_6796;
  wire       [35:0]   _zz_6797;
  wire       [35:0]   _zz_6798;
  wire       [35:0]   _zz_6799;
  wire       [35:0]   _zz_6800;
  wire       [26:0]   _zz_6801;
  wire       [35:0]   _zz_6802;
  wire       [17:0]   _zz_6803;
  wire       [35:0]   _zz_6804;
  wire       [35:0]   _zz_6805;
  wire       [35:0]   _zz_6806;
  wire       [35:0]   _zz_6807;
  wire       [35:0]   _zz_6808;
  wire       [26:0]   _zz_6809;
  wire       [35:0]   _zz_6810;
  wire       [17:0]   _zz_6811;
  wire       [35:0]   _zz_6812;
  wire       [35:0]   _zz_6813;
  wire       [35:0]   _zz_6814;
  wire       [35:0]   _zz_6815;
  wire       [35:0]   _zz_6816;
  wire       [26:0]   _zz_6817;
  wire       [35:0]   _zz_6818;
  wire       [17:0]   _zz_6819;
  wire       [35:0]   _zz_6820;
  wire       [35:0]   _zz_6821;
  wire       [35:0]   _zz_6822;
  wire       [35:0]   _zz_6823;
  wire       [35:0]   _zz_6824;
  wire       [26:0]   _zz_6825;
  wire       [35:0]   _zz_6826;
  wire       [17:0]   _zz_6827;
  wire       [17:0]   _zz_6828;
  wire       [35:0]   _zz_6829;
  wire       [35:0]   _zz_6830;
  wire       [17:0]   _zz_6831;
  wire       [35:0]   _zz_6832;
  wire       [35:0]   _zz_6833;
  wire       [35:0]   _zz_6834;
  wire       [17:0]   _zz_6835;
  wire       [35:0]   _zz_6836;
  wire       [35:0]   _zz_6837;
  wire       [35:0]   _zz_6838;
  wire       [35:0]   _zz_6839;
  wire       [35:0]   _zz_6840;
  wire       [35:0]   _zz_6841;
  wire       [26:0]   _zz_6842;
  wire       [35:0]   _zz_6843;
  wire       [17:0]   _zz_6844;
  wire       [35:0]   _zz_6845;
  wire       [35:0]   _zz_6846;
  wire       [35:0]   _zz_6847;
  wire       [35:0]   _zz_6848;
  wire       [35:0]   _zz_6849;
  wire       [26:0]   _zz_6850;
  wire       [35:0]   _zz_6851;
  wire       [17:0]   _zz_6852;
  wire       [35:0]   _zz_6853;
  wire       [35:0]   _zz_6854;
  wire       [35:0]   _zz_6855;
  wire       [35:0]   _zz_6856;
  wire       [35:0]   _zz_6857;
  wire       [26:0]   _zz_6858;
  wire       [35:0]   _zz_6859;
  wire       [17:0]   _zz_6860;
  wire       [35:0]   _zz_6861;
  wire       [35:0]   _zz_6862;
  wire       [35:0]   _zz_6863;
  wire       [35:0]   _zz_6864;
  wire       [35:0]   _zz_6865;
  wire       [26:0]   _zz_6866;
  wire       [35:0]   _zz_6867;
  wire       [17:0]   _zz_6868;
  wire       [17:0]   _zz_6869;
  wire       [35:0]   _zz_6870;
  wire       [35:0]   _zz_6871;
  wire       [17:0]   _zz_6872;
  wire       [35:0]   _zz_6873;
  wire       [35:0]   _zz_6874;
  wire       [35:0]   _zz_6875;
  wire       [17:0]   _zz_6876;
  wire       [35:0]   _zz_6877;
  wire       [35:0]   _zz_6878;
  wire       [35:0]   _zz_6879;
  wire       [35:0]   _zz_6880;
  wire       [35:0]   _zz_6881;
  wire       [35:0]   _zz_6882;
  wire       [26:0]   _zz_6883;
  wire       [35:0]   _zz_6884;
  wire       [17:0]   _zz_6885;
  wire       [35:0]   _zz_6886;
  wire       [35:0]   _zz_6887;
  wire       [35:0]   _zz_6888;
  wire       [35:0]   _zz_6889;
  wire       [35:0]   _zz_6890;
  wire       [26:0]   _zz_6891;
  wire       [35:0]   _zz_6892;
  wire       [17:0]   _zz_6893;
  wire       [35:0]   _zz_6894;
  wire       [35:0]   _zz_6895;
  wire       [35:0]   _zz_6896;
  wire       [35:0]   _zz_6897;
  wire       [35:0]   _zz_6898;
  wire       [26:0]   _zz_6899;
  wire       [35:0]   _zz_6900;
  wire       [17:0]   _zz_6901;
  wire       [35:0]   _zz_6902;
  wire       [35:0]   _zz_6903;
  wire       [35:0]   _zz_6904;
  wire       [35:0]   _zz_6905;
  wire       [35:0]   _zz_6906;
  wire       [26:0]   _zz_6907;
  wire       [35:0]   _zz_6908;
  wire       [17:0]   _zz_6909;
  wire       [17:0]   _zz_6910;
  wire       [35:0]   _zz_6911;
  wire       [35:0]   _zz_6912;
  wire       [17:0]   _zz_6913;
  wire       [35:0]   _zz_6914;
  wire       [35:0]   _zz_6915;
  wire       [35:0]   _zz_6916;
  wire       [17:0]   _zz_6917;
  wire       [35:0]   _zz_6918;
  wire       [35:0]   _zz_6919;
  wire       [35:0]   _zz_6920;
  wire       [35:0]   _zz_6921;
  wire       [35:0]   _zz_6922;
  wire       [35:0]   _zz_6923;
  wire       [26:0]   _zz_6924;
  wire       [35:0]   _zz_6925;
  wire       [17:0]   _zz_6926;
  wire       [35:0]   _zz_6927;
  wire       [35:0]   _zz_6928;
  wire       [35:0]   _zz_6929;
  wire       [35:0]   _zz_6930;
  wire       [35:0]   _zz_6931;
  wire       [26:0]   _zz_6932;
  wire       [35:0]   _zz_6933;
  wire       [17:0]   _zz_6934;
  wire       [35:0]   _zz_6935;
  wire       [35:0]   _zz_6936;
  wire       [35:0]   _zz_6937;
  wire       [35:0]   _zz_6938;
  wire       [35:0]   _zz_6939;
  wire       [26:0]   _zz_6940;
  wire       [35:0]   _zz_6941;
  wire       [17:0]   _zz_6942;
  wire       [35:0]   _zz_6943;
  wire       [35:0]   _zz_6944;
  wire       [35:0]   _zz_6945;
  wire       [35:0]   _zz_6946;
  wire       [35:0]   _zz_6947;
  wire       [26:0]   _zz_6948;
  wire       [35:0]   _zz_6949;
  wire       [17:0]   _zz_6950;
  wire       [17:0]   _zz_6951;
  wire       [35:0]   _zz_6952;
  wire       [35:0]   _zz_6953;
  wire       [17:0]   _zz_6954;
  wire       [35:0]   _zz_6955;
  wire       [35:0]   _zz_6956;
  wire       [35:0]   _zz_6957;
  wire       [17:0]   _zz_6958;
  wire       [35:0]   _zz_6959;
  wire       [35:0]   _zz_6960;
  wire       [35:0]   _zz_6961;
  wire       [35:0]   _zz_6962;
  wire       [35:0]   _zz_6963;
  wire       [35:0]   _zz_6964;
  wire       [26:0]   _zz_6965;
  wire       [35:0]   _zz_6966;
  wire       [17:0]   _zz_6967;
  wire       [35:0]   _zz_6968;
  wire       [35:0]   _zz_6969;
  wire       [35:0]   _zz_6970;
  wire       [35:0]   _zz_6971;
  wire       [35:0]   _zz_6972;
  wire       [26:0]   _zz_6973;
  wire       [35:0]   _zz_6974;
  wire       [17:0]   _zz_6975;
  wire       [35:0]   _zz_6976;
  wire       [35:0]   _zz_6977;
  wire       [35:0]   _zz_6978;
  wire       [35:0]   _zz_6979;
  wire       [35:0]   _zz_6980;
  wire       [26:0]   _zz_6981;
  wire       [35:0]   _zz_6982;
  wire       [17:0]   _zz_6983;
  wire       [35:0]   _zz_6984;
  wire       [35:0]   _zz_6985;
  wire       [35:0]   _zz_6986;
  wire       [35:0]   _zz_6987;
  wire       [35:0]   _zz_6988;
  wire       [26:0]   _zz_6989;
  wire       [35:0]   _zz_6990;
  wire       [17:0]   _zz_6991;
  wire       [17:0]   _zz_6992;
  wire       [35:0]   _zz_6993;
  wire       [35:0]   _zz_6994;
  wire       [17:0]   _zz_6995;
  wire       [35:0]   _zz_6996;
  wire       [35:0]   _zz_6997;
  wire       [35:0]   _zz_6998;
  wire       [17:0]   _zz_6999;
  wire       [35:0]   _zz_7000;
  wire       [35:0]   _zz_7001;
  wire       [35:0]   _zz_7002;
  wire       [35:0]   _zz_7003;
  wire       [35:0]   _zz_7004;
  wire       [35:0]   _zz_7005;
  wire       [26:0]   _zz_7006;
  wire       [35:0]   _zz_7007;
  wire       [17:0]   _zz_7008;
  wire       [35:0]   _zz_7009;
  wire       [35:0]   _zz_7010;
  wire       [35:0]   _zz_7011;
  wire       [35:0]   _zz_7012;
  wire       [35:0]   _zz_7013;
  wire       [26:0]   _zz_7014;
  wire       [35:0]   _zz_7015;
  wire       [17:0]   _zz_7016;
  wire       [35:0]   _zz_7017;
  wire       [35:0]   _zz_7018;
  wire       [35:0]   _zz_7019;
  wire       [35:0]   _zz_7020;
  wire       [35:0]   _zz_7021;
  wire       [26:0]   _zz_7022;
  wire       [35:0]   _zz_7023;
  wire       [17:0]   _zz_7024;
  wire       [35:0]   _zz_7025;
  wire       [35:0]   _zz_7026;
  wire       [35:0]   _zz_7027;
  wire       [35:0]   _zz_7028;
  wire       [35:0]   _zz_7029;
  wire       [26:0]   _zz_7030;
  wire       [35:0]   _zz_7031;
  wire       [17:0]   _zz_7032;
  wire       [17:0]   _zz_7033;
  wire       [35:0]   _zz_7034;
  wire       [35:0]   _zz_7035;
  wire       [17:0]   _zz_7036;
  wire       [35:0]   _zz_7037;
  wire       [35:0]   _zz_7038;
  wire       [35:0]   _zz_7039;
  wire       [17:0]   _zz_7040;
  wire       [35:0]   _zz_7041;
  wire       [35:0]   _zz_7042;
  wire       [35:0]   _zz_7043;
  wire       [35:0]   _zz_7044;
  wire       [35:0]   _zz_7045;
  wire       [35:0]   _zz_7046;
  wire       [26:0]   _zz_7047;
  wire       [35:0]   _zz_7048;
  wire       [17:0]   _zz_7049;
  wire       [35:0]   _zz_7050;
  wire       [35:0]   _zz_7051;
  wire       [35:0]   _zz_7052;
  wire       [35:0]   _zz_7053;
  wire       [35:0]   _zz_7054;
  wire       [26:0]   _zz_7055;
  wire       [35:0]   _zz_7056;
  wire       [17:0]   _zz_7057;
  wire       [35:0]   _zz_7058;
  wire       [35:0]   _zz_7059;
  wire       [35:0]   _zz_7060;
  wire       [35:0]   _zz_7061;
  wire       [35:0]   _zz_7062;
  wire       [26:0]   _zz_7063;
  wire       [35:0]   _zz_7064;
  wire       [17:0]   _zz_7065;
  wire       [35:0]   _zz_7066;
  wire       [35:0]   _zz_7067;
  wire       [35:0]   _zz_7068;
  wire       [35:0]   _zz_7069;
  wire       [35:0]   _zz_7070;
  wire       [26:0]   _zz_7071;
  wire       [35:0]   _zz_7072;
  wire       [17:0]   _zz_7073;
  wire       [17:0]   _zz_7074;
  wire       [35:0]   _zz_7075;
  wire       [35:0]   _zz_7076;
  wire       [17:0]   _zz_7077;
  wire       [35:0]   _zz_7078;
  wire       [35:0]   _zz_7079;
  wire       [35:0]   _zz_7080;
  wire       [17:0]   _zz_7081;
  wire       [35:0]   _zz_7082;
  wire       [35:0]   _zz_7083;
  wire       [35:0]   _zz_7084;
  wire       [35:0]   _zz_7085;
  wire       [35:0]   _zz_7086;
  wire       [35:0]   _zz_7087;
  wire       [26:0]   _zz_7088;
  wire       [35:0]   _zz_7089;
  wire       [17:0]   _zz_7090;
  wire       [35:0]   _zz_7091;
  wire       [35:0]   _zz_7092;
  wire       [35:0]   _zz_7093;
  wire       [35:0]   _zz_7094;
  wire       [35:0]   _zz_7095;
  wire       [26:0]   _zz_7096;
  wire       [35:0]   _zz_7097;
  wire       [17:0]   _zz_7098;
  wire       [35:0]   _zz_7099;
  wire       [35:0]   _zz_7100;
  wire       [35:0]   _zz_7101;
  wire       [35:0]   _zz_7102;
  wire       [35:0]   _zz_7103;
  wire       [26:0]   _zz_7104;
  wire       [35:0]   _zz_7105;
  wire       [17:0]   _zz_7106;
  wire       [35:0]   _zz_7107;
  wire       [35:0]   _zz_7108;
  wire       [35:0]   _zz_7109;
  wire       [35:0]   _zz_7110;
  wire       [35:0]   _zz_7111;
  wire       [26:0]   _zz_7112;
  wire       [35:0]   _zz_7113;
  wire       [17:0]   _zz_7114;
  wire       [17:0]   _zz_7115;
  wire       [35:0]   _zz_7116;
  wire       [35:0]   _zz_7117;
  wire       [17:0]   _zz_7118;
  wire       [35:0]   _zz_7119;
  wire       [35:0]   _zz_7120;
  wire       [35:0]   _zz_7121;
  wire       [17:0]   _zz_7122;
  wire       [35:0]   _zz_7123;
  wire       [35:0]   _zz_7124;
  wire       [35:0]   _zz_7125;
  wire       [35:0]   _zz_7126;
  wire       [35:0]   _zz_7127;
  wire       [35:0]   _zz_7128;
  wire       [26:0]   _zz_7129;
  wire       [35:0]   _zz_7130;
  wire       [17:0]   _zz_7131;
  wire       [35:0]   _zz_7132;
  wire       [35:0]   _zz_7133;
  wire       [35:0]   _zz_7134;
  wire       [35:0]   _zz_7135;
  wire       [35:0]   _zz_7136;
  wire       [26:0]   _zz_7137;
  wire       [35:0]   _zz_7138;
  wire       [17:0]   _zz_7139;
  wire       [35:0]   _zz_7140;
  wire       [35:0]   _zz_7141;
  wire       [35:0]   _zz_7142;
  wire       [35:0]   _zz_7143;
  wire       [35:0]   _zz_7144;
  wire       [26:0]   _zz_7145;
  wire       [35:0]   _zz_7146;
  wire       [17:0]   _zz_7147;
  wire       [35:0]   _zz_7148;
  wire       [35:0]   _zz_7149;
  wire       [35:0]   _zz_7150;
  wire       [35:0]   _zz_7151;
  wire       [35:0]   _zz_7152;
  wire       [26:0]   _zz_7153;
  wire       [35:0]   _zz_7154;
  wire       [17:0]   _zz_7155;
  wire       [17:0]   _zz_7156;
  wire       [35:0]   _zz_7157;
  wire       [35:0]   _zz_7158;
  wire       [17:0]   _zz_7159;
  wire       [35:0]   _zz_7160;
  wire       [35:0]   _zz_7161;
  wire       [35:0]   _zz_7162;
  wire       [17:0]   _zz_7163;
  wire       [35:0]   _zz_7164;
  wire       [35:0]   _zz_7165;
  wire       [35:0]   _zz_7166;
  wire       [35:0]   _zz_7167;
  wire       [35:0]   _zz_7168;
  wire       [35:0]   _zz_7169;
  wire       [26:0]   _zz_7170;
  wire       [35:0]   _zz_7171;
  wire       [17:0]   _zz_7172;
  wire       [35:0]   _zz_7173;
  wire       [35:0]   _zz_7174;
  wire       [35:0]   _zz_7175;
  wire       [35:0]   _zz_7176;
  wire       [35:0]   _zz_7177;
  wire       [26:0]   _zz_7178;
  wire       [35:0]   _zz_7179;
  wire       [17:0]   _zz_7180;
  wire       [35:0]   _zz_7181;
  wire       [35:0]   _zz_7182;
  wire       [35:0]   _zz_7183;
  wire       [35:0]   _zz_7184;
  wire       [35:0]   _zz_7185;
  wire       [26:0]   _zz_7186;
  wire       [35:0]   _zz_7187;
  wire       [17:0]   _zz_7188;
  wire       [35:0]   _zz_7189;
  wire       [35:0]   _zz_7190;
  wire       [35:0]   _zz_7191;
  wire       [35:0]   _zz_7192;
  wire       [35:0]   _zz_7193;
  wire       [26:0]   _zz_7194;
  wire       [35:0]   _zz_7195;
  wire       [17:0]   _zz_7196;
  wire       [17:0]   _zz_7197;
  wire       [35:0]   _zz_7198;
  wire       [35:0]   _zz_7199;
  wire       [17:0]   _zz_7200;
  wire       [35:0]   _zz_7201;
  wire       [35:0]   _zz_7202;
  wire       [35:0]   _zz_7203;
  wire       [17:0]   _zz_7204;
  wire       [35:0]   _zz_7205;
  wire       [35:0]   _zz_7206;
  wire       [35:0]   _zz_7207;
  wire       [35:0]   _zz_7208;
  wire       [35:0]   _zz_7209;
  wire       [35:0]   _zz_7210;
  wire       [26:0]   _zz_7211;
  wire       [35:0]   _zz_7212;
  wire       [17:0]   _zz_7213;
  wire       [35:0]   _zz_7214;
  wire       [35:0]   _zz_7215;
  wire       [35:0]   _zz_7216;
  wire       [35:0]   _zz_7217;
  wire       [35:0]   _zz_7218;
  wire       [26:0]   _zz_7219;
  wire       [35:0]   _zz_7220;
  wire       [17:0]   _zz_7221;
  wire       [35:0]   _zz_7222;
  wire       [35:0]   _zz_7223;
  wire       [35:0]   _zz_7224;
  wire       [35:0]   _zz_7225;
  wire       [35:0]   _zz_7226;
  wire       [26:0]   _zz_7227;
  wire       [35:0]   _zz_7228;
  wire       [17:0]   _zz_7229;
  wire       [35:0]   _zz_7230;
  wire       [35:0]   _zz_7231;
  wire       [35:0]   _zz_7232;
  wire       [35:0]   _zz_7233;
  wire       [35:0]   _zz_7234;
  wire       [26:0]   _zz_7235;
  wire       [35:0]   _zz_7236;
  wire       [17:0]   _zz_7237;
  wire       [17:0]   _zz_7238;
  wire       [35:0]   _zz_7239;
  wire       [35:0]   _zz_7240;
  wire       [17:0]   _zz_7241;
  wire       [35:0]   _zz_7242;
  wire       [35:0]   _zz_7243;
  wire       [35:0]   _zz_7244;
  wire       [17:0]   _zz_7245;
  wire       [35:0]   _zz_7246;
  wire       [35:0]   _zz_7247;
  wire       [35:0]   _zz_7248;
  wire       [35:0]   _zz_7249;
  wire       [35:0]   _zz_7250;
  wire       [35:0]   _zz_7251;
  wire       [26:0]   _zz_7252;
  wire       [35:0]   _zz_7253;
  wire       [17:0]   _zz_7254;
  wire       [35:0]   _zz_7255;
  wire       [35:0]   _zz_7256;
  wire       [35:0]   _zz_7257;
  wire       [35:0]   _zz_7258;
  wire       [35:0]   _zz_7259;
  wire       [26:0]   _zz_7260;
  wire       [35:0]   _zz_7261;
  wire       [17:0]   _zz_7262;
  wire       [35:0]   _zz_7263;
  wire       [35:0]   _zz_7264;
  wire       [35:0]   _zz_7265;
  wire       [35:0]   _zz_7266;
  wire       [35:0]   _zz_7267;
  wire       [26:0]   _zz_7268;
  wire       [35:0]   _zz_7269;
  wire       [17:0]   _zz_7270;
  wire       [35:0]   _zz_7271;
  wire       [35:0]   _zz_7272;
  wire       [35:0]   _zz_7273;
  wire       [35:0]   _zz_7274;
  wire       [35:0]   _zz_7275;
  wire       [26:0]   _zz_7276;
  wire       [35:0]   _zz_7277;
  wire       [17:0]   _zz_7278;
  wire       [17:0]   _zz_7279;
  wire       [35:0]   _zz_7280;
  wire       [35:0]   _zz_7281;
  wire       [17:0]   _zz_7282;
  wire       [35:0]   _zz_7283;
  wire       [35:0]   _zz_7284;
  wire       [35:0]   _zz_7285;
  wire       [17:0]   _zz_7286;
  wire       [35:0]   _zz_7287;
  wire       [35:0]   _zz_7288;
  wire       [35:0]   _zz_7289;
  wire       [35:0]   _zz_7290;
  wire       [35:0]   _zz_7291;
  wire       [35:0]   _zz_7292;
  wire       [26:0]   _zz_7293;
  wire       [35:0]   _zz_7294;
  wire       [17:0]   _zz_7295;
  wire       [35:0]   _zz_7296;
  wire       [35:0]   _zz_7297;
  wire       [35:0]   _zz_7298;
  wire       [35:0]   _zz_7299;
  wire       [35:0]   _zz_7300;
  wire       [26:0]   _zz_7301;
  wire       [35:0]   _zz_7302;
  wire       [17:0]   _zz_7303;
  wire       [35:0]   _zz_7304;
  wire       [35:0]   _zz_7305;
  wire       [35:0]   _zz_7306;
  wire       [35:0]   _zz_7307;
  wire       [35:0]   _zz_7308;
  wire       [26:0]   _zz_7309;
  wire       [35:0]   _zz_7310;
  wire       [17:0]   _zz_7311;
  wire       [35:0]   _zz_7312;
  wire       [35:0]   _zz_7313;
  wire       [35:0]   _zz_7314;
  wire       [35:0]   _zz_7315;
  wire       [35:0]   _zz_7316;
  wire       [26:0]   _zz_7317;
  wire       [35:0]   _zz_7318;
  wire       [17:0]   _zz_7319;
  wire       [17:0]   _zz_7320;
  wire       [35:0]   _zz_7321;
  wire       [35:0]   _zz_7322;
  wire       [17:0]   _zz_7323;
  wire       [35:0]   _zz_7324;
  wire       [35:0]   _zz_7325;
  wire       [35:0]   _zz_7326;
  wire       [17:0]   _zz_7327;
  wire       [35:0]   _zz_7328;
  wire       [35:0]   _zz_7329;
  wire       [35:0]   _zz_7330;
  wire       [35:0]   _zz_7331;
  wire       [35:0]   _zz_7332;
  wire       [35:0]   _zz_7333;
  wire       [26:0]   _zz_7334;
  wire       [35:0]   _zz_7335;
  wire       [17:0]   _zz_7336;
  wire       [35:0]   _zz_7337;
  wire       [35:0]   _zz_7338;
  wire       [35:0]   _zz_7339;
  wire       [35:0]   _zz_7340;
  wire       [35:0]   _zz_7341;
  wire       [26:0]   _zz_7342;
  wire       [35:0]   _zz_7343;
  wire       [17:0]   _zz_7344;
  wire       [35:0]   _zz_7345;
  wire       [35:0]   _zz_7346;
  wire       [35:0]   _zz_7347;
  wire       [35:0]   _zz_7348;
  wire       [35:0]   _zz_7349;
  wire       [26:0]   _zz_7350;
  wire       [35:0]   _zz_7351;
  wire       [17:0]   _zz_7352;
  wire       [35:0]   _zz_7353;
  wire       [35:0]   _zz_7354;
  wire       [35:0]   _zz_7355;
  wire       [35:0]   _zz_7356;
  wire       [35:0]   _zz_7357;
  wire       [26:0]   _zz_7358;
  wire       [35:0]   _zz_7359;
  wire       [17:0]   _zz_7360;
  wire       [17:0]   _zz_7361;
  wire       [35:0]   _zz_7362;
  wire       [35:0]   _zz_7363;
  wire       [17:0]   _zz_7364;
  wire       [35:0]   _zz_7365;
  wire       [35:0]   _zz_7366;
  wire       [35:0]   _zz_7367;
  wire       [17:0]   _zz_7368;
  wire       [35:0]   _zz_7369;
  wire       [35:0]   _zz_7370;
  wire       [35:0]   _zz_7371;
  wire       [35:0]   _zz_7372;
  wire       [35:0]   _zz_7373;
  wire       [35:0]   _zz_7374;
  wire       [26:0]   _zz_7375;
  wire       [35:0]   _zz_7376;
  wire       [17:0]   _zz_7377;
  wire       [35:0]   _zz_7378;
  wire       [35:0]   _zz_7379;
  wire       [35:0]   _zz_7380;
  wire       [35:0]   _zz_7381;
  wire       [35:0]   _zz_7382;
  wire       [26:0]   _zz_7383;
  wire       [35:0]   _zz_7384;
  wire       [17:0]   _zz_7385;
  wire       [35:0]   _zz_7386;
  wire       [35:0]   _zz_7387;
  wire       [35:0]   _zz_7388;
  wire       [35:0]   _zz_7389;
  wire       [35:0]   _zz_7390;
  wire       [26:0]   _zz_7391;
  wire       [35:0]   _zz_7392;
  wire       [17:0]   _zz_7393;
  wire       [35:0]   _zz_7394;
  wire       [35:0]   _zz_7395;
  wire       [35:0]   _zz_7396;
  wire       [35:0]   _zz_7397;
  wire       [35:0]   _zz_7398;
  wire       [26:0]   _zz_7399;
  wire       [35:0]   _zz_7400;
  wire       [17:0]   _zz_7401;
  wire       [17:0]   _zz_7402;
  wire       [35:0]   _zz_7403;
  wire       [35:0]   _zz_7404;
  wire       [17:0]   _zz_7405;
  wire       [35:0]   _zz_7406;
  wire       [35:0]   _zz_7407;
  wire       [35:0]   _zz_7408;
  wire       [17:0]   _zz_7409;
  wire       [35:0]   _zz_7410;
  wire       [35:0]   _zz_7411;
  wire       [35:0]   _zz_7412;
  wire       [35:0]   _zz_7413;
  wire       [35:0]   _zz_7414;
  wire       [35:0]   _zz_7415;
  wire       [26:0]   _zz_7416;
  wire       [35:0]   _zz_7417;
  wire       [17:0]   _zz_7418;
  wire       [35:0]   _zz_7419;
  wire       [35:0]   _zz_7420;
  wire       [35:0]   _zz_7421;
  wire       [35:0]   _zz_7422;
  wire       [35:0]   _zz_7423;
  wire       [26:0]   _zz_7424;
  wire       [35:0]   _zz_7425;
  wire       [17:0]   _zz_7426;
  wire       [35:0]   _zz_7427;
  wire       [35:0]   _zz_7428;
  wire       [35:0]   _zz_7429;
  wire       [35:0]   _zz_7430;
  wire       [35:0]   _zz_7431;
  wire       [26:0]   _zz_7432;
  wire       [35:0]   _zz_7433;
  wire       [17:0]   _zz_7434;
  wire       [35:0]   _zz_7435;
  wire       [35:0]   _zz_7436;
  wire       [35:0]   _zz_7437;
  wire       [35:0]   _zz_7438;
  wire       [35:0]   _zz_7439;
  wire       [26:0]   _zz_7440;
  wire       [35:0]   _zz_7441;
  wire       [17:0]   _zz_7442;
  wire       [17:0]   _zz_7443;
  wire       [35:0]   _zz_7444;
  wire       [35:0]   _zz_7445;
  wire       [17:0]   _zz_7446;
  wire       [35:0]   _zz_7447;
  wire       [35:0]   _zz_7448;
  wire       [35:0]   _zz_7449;
  wire       [17:0]   _zz_7450;
  wire       [35:0]   _zz_7451;
  wire       [35:0]   _zz_7452;
  wire       [35:0]   _zz_7453;
  wire       [35:0]   _zz_7454;
  wire       [35:0]   _zz_7455;
  wire       [35:0]   _zz_7456;
  wire       [26:0]   _zz_7457;
  wire       [35:0]   _zz_7458;
  wire       [17:0]   _zz_7459;
  wire       [35:0]   _zz_7460;
  wire       [35:0]   _zz_7461;
  wire       [35:0]   _zz_7462;
  wire       [35:0]   _zz_7463;
  wire       [35:0]   _zz_7464;
  wire       [26:0]   _zz_7465;
  wire       [35:0]   _zz_7466;
  wire       [17:0]   _zz_7467;
  wire       [35:0]   _zz_7468;
  wire       [35:0]   _zz_7469;
  wire       [35:0]   _zz_7470;
  wire       [35:0]   _zz_7471;
  wire       [35:0]   _zz_7472;
  wire       [26:0]   _zz_7473;
  wire       [35:0]   _zz_7474;
  wire       [17:0]   _zz_7475;
  wire       [35:0]   _zz_7476;
  wire       [35:0]   _zz_7477;
  wire       [35:0]   _zz_7478;
  wire       [35:0]   _zz_7479;
  wire       [35:0]   _zz_7480;
  wire       [26:0]   _zz_7481;
  wire       [35:0]   _zz_7482;
  wire       [17:0]   _zz_7483;
  wire       [17:0]   _zz_7484;
  wire       [35:0]   _zz_7485;
  wire       [35:0]   _zz_7486;
  wire       [17:0]   _zz_7487;
  wire       [35:0]   _zz_7488;
  wire       [35:0]   _zz_7489;
  wire       [35:0]   _zz_7490;
  wire       [17:0]   _zz_7491;
  wire       [35:0]   _zz_7492;
  wire       [35:0]   _zz_7493;
  wire       [35:0]   _zz_7494;
  wire       [35:0]   _zz_7495;
  wire       [35:0]   _zz_7496;
  wire       [35:0]   _zz_7497;
  wire       [26:0]   _zz_7498;
  wire       [35:0]   _zz_7499;
  wire       [17:0]   _zz_7500;
  wire       [35:0]   _zz_7501;
  wire       [35:0]   _zz_7502;
  wire       [35:0]   _zz_7503;
  wire       [35:0]   _zz_7504;
  wire       [35:0]   _zz_7505;
  wire       [26:0]   _zz_7506;
  wire       [35:0]   _zz_7507;
  wire       [17:0]   _zz_7508;
  wire       [35:0]   _zz_7509;
  wire       [35:0]   _zz_7510;
  wire       [35:0]   _zz_7511;
  wire       [35:0]   _zz_7512;
  wire       [35:0]   _zz_7513;
  wire       [26:0]   _zz_7514;
  wire       [35:0]   _zz_7515;
  wire       [17:0]   _zz_7516;
  wire       [35:0]   _zz_7517;
  wire       [35:0]   _zz_7518;
  wire       [35:0]   _zz_7519;
  wire       [35:0]   _zz_7520;
  wire       [35:0]   _zz_7521;
  wire       [26:0]   _zz_7522;
  wire       [35:0]   _zz_7523;
  wire       [17:0]   _zz_7524;
  wire       [17:0]   _zz_7525;
  wire       [35:0]   _zz_7526;
  wire       [35:0]   _zz_7527;
  wire       [17:0]   _zz_7528;
  wire       [35:0]   _zz_7529;
  wire       [35:0]   _zz_7530;
  wire       [35:0]   _zz_7531;
  wire       [17:0]   _zz_7532;
  wire       [35:0]   _zz_7533;
  wire       [35:0]   _zz_7534;
  wire       [35:0]   _zz_7535;
  wire       [35:0]   _zz_7536;
  wire       [35:0]   _zz_7537;
  wire       [35:0]   _zz_7538;
  wire       [26:0]   _zz_7539;
  wire       [35:0]   _zz_7540;
  wire       [17:0]   _zz_7541;
  wire       [35:0]   _zz_7542;
  wire       [35:0]   _zz_7543;
  wire       [35:0]   _zz_7544;
  wire       [35:0]   _zz_7545;
  wire       [35:0]   _zz_7546;
  wire       [26:0]   _zz_7547;
  wire       [35:0]   _zz_7548;
  wire       [17:0]   _zz_7549;
  wire       [35:0]   _zz_7550;
  wire       [35:0]   _zz_7551;
  wire       [35:0]   _zz_7552;
  wire       [35:0]   _zz_7553;
  wire       [35:0]   _zz_7554;
  wire       [26:0]   _zz_7555;
  wire       [35:0]   _zz_7556;
  wire       [17:0]   _zz_7557;
  wire       [35:0]   _zz_7558;
  wire       [35:0]   _zz_7559;
  wire       [35:0]   _zz_7560;
  wire       [35:0]   _zz_7561;
  wire       [35:0]   _zz_7562;
  wire       [26:0]   _zz_7563;
  wire       [35:0]   _zz_7564;
  wire       [17:0]   _zz_7565;
  wire       [17:0]   _zz_7566;
  wire       [35:0]   _zz_7567;
  wire       [35:0]   _zz_7568;
  wire       [17:0]   _zz_7569;
  wire       [35:0]   _zz_7570;
  wire       [35:0]   _zz_7571;
  wire       [35:0]   _zz_7572;
  wire       [17:0]   _zz_7573;
  wire       [35:0]   _zz_7574;
  wire       [35:0]   _zz_7575;
  wire       [35:0]   _zz_7576;
  wire       [35:0]   _zz_7577;
  wire       [35:0]   _zz_7578;
  wire       [35:0]   _zz_7579;
  wire       [26:0]   _zz_7580;
  wire       [35:0]   _zz_7581;
  wire       [17:0]   _zz_7582;
  wire       [35:0]   _zz_7583;
  wire       [35:0]   _zz_7584;
  wire       [35:0]   _zz_7585;
  wire       [35:0]   _zz_7586;
  wire       [35:0]   _zz_7587;
  wire       [26:0]   _zz_7588;
  wire       [35:0]   _zz_7589;
  wire       [17:0]   _zz_7590;
  wire       [35:0]   _zz_7591;
  wire       [35:0]   _zz_7592;
  wire       [35:0]   _zz_7593;
  wire       [35:0]   _zz_7594;
  wire       [35:0]   _zz_7595;
  wire       [26:0]   _zz_7596;
  wire       [35:0]   _zz_7597;
  wire       [17:0]   _zz_7598;
  wire       [35:0]   _zz_7599;
  wire       [35:0]   _zz_7600;
  wire       [35:0]   _zz_7601;
  wire       [35:0]   _zz_7602;
  wire       [35:0]   _zz_7603;
  wire       [26:0]   _zz_7604;
  wire       [35:0]   _zz_7605;
  wire       [17:0]   _zz_7606;
  wire       [17:0]   _zz_7607;
  wire       [35:0]   _zz_7608;
  wire       [35:0]   _zz_7609;
  wire       [17:0]   _zz_7610;
  wire       [35:0]   _zz_7611;
  wire       [35:0]   _zz_7612;
  wire       [35:0]   _zz_7613;
  wire       [17:0]   _zz_7614;
  wire       [35:0]   _zz_7615;
  wire       [35:0]   _zz_7616;
  wire       [35:0]   _zz_7617;
  wire       [35:0]   _zz_7618;
  wire       [35:0]   _zz_7619;
  wire       [35:0]   _zz_7620;
  wire       [26:0]   _zz_7621;
  wire       [35:0]   _zz_7622;
  wire       [17:0]   _zz_7623;
  wire       [35:0]   _zz_7624;
  wire       [35:0]   _zz_7625;
  wire       [35:0]   _zz_7626;
  wire       [35:0]   _zz_7627;
  wire       [35:0]   _zz_7628;
  wire       [26:0]   _zz_7629;
  wire       [35:0]   _zz_7630;
  wire       [17:0]   _zz_7631;
  wire       [35:0]   _zz_7632;
  wire       [35:0]   _zz_7633;
  wire       [35:0]   _zz_7634;
  wire       [35:0]   _zz_7635;
  wire       [35:0]   _zz_7636;
  wire       [26:0]   _zz_7637;
  wire       [35:0]   _zz_7638;
  wire       [17:0]   _zz_7639;
  wire       [35:0]   _zz_7640;
  wire       [35:0]   _zz_7641;
  wire       [35:0]   _zz_7642;
  wire       [35:0]   _zz_7643;
  wire       [35:0]   _zz_7644;
  wire       [26:0]   _zz_7645;
  wire       [35:0]   _zz_7646;
  wire       [17:0]   _zz_7647;
  wire       [17:0]   _zz_7648;
  wire       [35:0]   _zz_7649;
  wire       [35:0]   _zz_7650;
  wire       [17:0]   _zz_7651;
  wire       [35:0]   _zz_7652;
  wire       [35:0]   _zz_7653;
  wire       [35:0]   _zz_7654;
  wire       [17:0]   _zz_7655;
  wire       [35:0]   _zz_7656;
  wire       [35:0]   _zz_7657;
  wire       [35:0]   _zz_7658;
  wire       [35:0]   _zz_7659;
  wire       [35:0]   _zz_7660;
  wire       [35:0]   _zz_7661;
  wire       [26:0]   _zz_7662;
  wire       [35:0]   _zz_7663;
  wire       [17:0]   _zz_7664;
  wire       [35:0]   _zz_7665;
  wire       [35:0]   _zz_7666;
  wire       [35:0]   _zz_7667;
  wire       [35:0]   _zz_7668;
  wire       [35:0]   _zz_7669;
  wire       [26:0]   _zz_7670;
  wire       [35:0]   _zz_7671;
  wire       [17:0]   _zz_7672;
  wire       [35:0]   _zz_7673;
  wire       [35:0]   _zz_7674;
  wire       [35:0]   _zz_7675;
  wire       [35:0]   _zz_7676;
  wire       [35:0]   _zz_7677;
  wire       [26:0]   _zz_7678;
  wire       [35:0]   _zz_7679;
  wire       [17:0]   _zz_7680;
  wire       [35:0]   _zz_7681;
  wire       [35:0]   _zz_7682;
  wire       [35:0]   _zz_7683;
  wire       [35:0]   _zz_7684;
  wire       [35:0]   _zz_7685;
  wire       [26:0]   _zz_7686;
  wire       [35:0]   _zz_7687;
  wire       [17:0]   _zz_7688;
  wire       [17:0]   _zz_7689;
  wire       [35:0]   _zz_7690;
  wire       [35:0]   _zz_7691;
  wire       [17:0]   _zz_7692;
  wire       [35:0]   _zz_7693;
  wire       [35:0]   _zz_7694;
  wire       [35:0]   _zz_7695;
  wire       [17:0]   _zz_7696;
  wire       [35:0]   _zz_7697;
  wire       [35:0]   _zz_7698;
  wire       [35:0]   _zz_7699;
  wire       [35:0]   _zz_7700;
  wire       [35:0]   _zz_7701;
  wire       [35:0]   _zz_7702;
  wire       [26:0]   _zz_7703;
  wire       [35:0]   _zz_7704;
  wire       [17:0]   _zz_7705;
  wire       [35:0]   _zz_7706;
  wire       [35:0]   _zz_7707;
  wire       [35:0]   _zz_7708;
  wire       [35:0]   _zz_7709;
  wire       [35:0]   _zz_7710;
  wire       [26:0]   _zz_7711;
  wire       [35:0]   _zz_7712;
  wire       [17:0]   _zz_7713;
  wire       [35:0]   _zz_7714;
  wire       [35:0]   _zz_7715;
  wire       [35:0]   _zz_7716;
  wire       [35:0]   _zz_7717;
  wire       [35:0]   _zz_7718;
  wire       [26:0]   _zz_7719;
  wire       [35:0]   _zz_7720;
  wire       [17:0]   _zz_7721;
  wire       [35:0]   _zz_7722;
  wire       [35:0]   _zz_7723;
  wire       [35:0]   _zz_7724;
  wire       [35:0]   _zz_7725;
  wire       [35:0]   _zz_7726;
  wire       [26:0]   _zz_7727;
  wire       [35:0]   _zz_7728;
  wire       [17:0]   _zz_7729;
  wire       [17:0]   _zz_7730;
  wire       [35:0]   _zz_7731;
  wire       [35:0]   _zz_7732;
  wire       [17:0]   _zz_7733;
  wire       [35:0]   _zz_7734;
  wire       [35:0]   _zz_7735;
  wire       [35:0]   _zz_7736;
  wire       [17:0]   _zz_7737;
  wire       [35:0]   _zz_7738;
  wire       [35:0]   _zz_7739;
  wire       [35:0]   _zz_7740;
  wire       [35:0]   _zz_7741;
  wire       [35:0]   _zz_7742;
  wire       [35:0]   _zz_7743;
  wire       [26:0]   _zz_7744;
  wire       [35:0]   _zz_7745;
  wire       [17:0]   _zz_7746;
  wire       [35:0]   _zz_7747;
  wire       [35:0]   _zz_7748;
  wire       [35:0]   _zz_7749;
  wire       [35:0]   _zz_7750;
  wire       [35:0]   _zz_7751;
  wire       [26:0]   _zz_7752;
  wire       [35:0]   _zz_7753;
  wire       [17:0]   _zz_7754;
  wire       [35:0]   _zz_7755;
  wire       [35:0]   _zz_7756;
  wire       [35:0]   _zz_7757;
  wire       [35:0]   _zz_7758;
  wire       [35:0]   _zz_7759;
  wire       [26:0]   _zz_7760;
  wire       [35:0]   _zz_7761;
  wire       [17:0]   _zz_7762;
  wire       [35:0]   _zz_7763;
  wire       [35:0]   _zz_7764;
  wire       [35:0]   _zz_7765;
  wire       [35:0]   _zz_7766;
  wire       [35:0]   _zz_7767;
  wire       [26:0]   _zz_7768;
  wire       [35:0]   _zz_7769;
  wire       [17:0]   _zz_7770;
  wire       [17:0]   _zz_7771;
  wire       [35:0]   _zz_7772;
  wire       [35:0]   _zz_7773;
  wire       [17:0]   _zz_7774;
  wire       [35:0]   _zz_7775;
  wire       [35:0]   _zz_7776;
  wire       [35:0]   _zz_7777;
  wire       [17:0]   _zz_7778;
  wire       [35:0]   _zz_7779;
  wire       [35:0]   _zz_7780;
  wire       [35:0]   _zz_7781;
  wire       [35:0]   _zz_7782;
  wire       [35:0]   _zz_7783;
  wire       [35:0]   _zz_7784;
  wire       [26:0]   _zz_7785;
  wire       [35:0]   _zz_7786;
  wire       [17:0]   _zz_7787;
  wire       [35:0]   _zz_7788;
  wire       [35:0]   _zz_7789;
  wire       [35:0]   _zz_7790;
  wire       [35:0]   _zz_7791;
  wire       [35:0]   _zz_7792;
  wire       [26:0]   _zz_7793;
  wire       [35:0]   _zz_7794;
  wire       [17:0]   _zz_7795;
  wire       [35:0]   _zz_7796;
  wire       [35:0]   _zz_7797;
  wire       [35:0]   _zz_7798;
  wire       [35:0]   _zz_7799;
  wire       [35:0]   _zz_7800;
  wire       [26:0]   _zz_7801;
  wire       [35:0]   _zz_7802;
  wire       [17:0]   _zz_7803;
  wire       [35:0]   _zz_7804;
  wire       [35:0]   _zz_7805;
  wire       [35:0]   _zz_7806;
  wire       [35:0]   _zz_7807;
  wire       [35:0]   _zz_7808;
  wire       [26:0]   _zz_7809;
  wire       [35:0]   _zz_7810;
  wire       [17:0]   _zz_7811;
  wire       [17:0]   _zz_7812;
  wire       [35:0]   _zz_7813;
  wire       [35:0]   _zz_7814;
  wire       [17:0]   _zz_7815;
  wire       [35:0]   _zz_7816;
  wire       [35:0]   _zz_7817;
  wire       [35:0]   _zz_7818;
  wire       [17:0]   _zz_7819;
  wire       [35:0]   _zz_7820;
  wire       [35:0]   _zz_7821;
  wire       [35:0]   _zz_7822;
  wire       [35:0]   _zz_7823;
  wire       [35:0]   _zz_7824;
  wire       [35:0]   _zz_7825;
  wire       [26:0]   _zz_7826;
  wire       [35:0]   _zz_7827;
  wire       [17:0]   _zz_7828;
  wire       [35:0]   _zz_7829;
  wire       [35:0]   _zz_7830;
  wire       [35:0]   _zz_7831;
  wire       [35:0]   _zz_7832;
  wire       [35:0]   _zz_7833;
  wire       [26:0]   _zz_7834;
  wire       [35:0]   _zz_7835;
  wire       [17:0]   _zz_7836;
  wire       [35:0]   _zz_7837;
  wire       [35:0]   _zz_7838;
  wire       [35:0]   _zz_7839;
  wire       [35:0]   _zz_7840;
  wire       [35:0]   _zz_7841;
  wire       [26:0]   _zz_7842;
  wire       [35:0]   _zz_7843;
  wire       [17:0]   _zz_7844;
  wire       [35:0]   _zz_7845;
  wire       [35:0]   _zz_7846;
  wire       [35:0]   _zz_7847;
  wire       [35:0]   _zz_7848;
  wire       [35:0]   _zz_7849;
  wire       [26:0]   _zz_7850;
  wire       [35:0]   _zz_7851;
  wire       [17:0]   _zz_7852;
  wire       [17:0]   _zz_7853;
  wire       [35:0]   _zz_7854;
  wire       [35:0]   _zz_7855;
  wire       [17:0]   _zz_7856;
  wire       [35:0]   _zz_7857;
  wire       [35:0]   _zz_7858;
  wire       [35:0]   _zz_7859;
  wire       [17:0]   _zz_7860;
  wire       [35:0]   _zz_7861;
  wire       [35:0]   _zz_7862;
  wire       [35:0]   _zz_7863;
  wire       [35:0]   _zz_7864;
  wire       [35:0]   _zz_7865;
  wire       [35:0]   _zz_7866;
  wire       [26:0]   _zz_7867;
  wire       [35:0]   _zz_7868;
  wire       [17:0]   _zz_7869;
  wire       [35:0]   _zz_7870;
  wire       [35:0]   _zz_7871;
  wire       [35:0]   _zz_7872;
  wire       [35:0]   _zz_7873;
  wire       [35:0]   _zz_7874;
  wire       [26:0]   _zz_7875;
  wire       [35:0]   _zz_7876;
  wire       [17:0]   _zz_7877;
  wire       [35:0]   _zz_7878;
  wire       [35:0]   _zz_7879;
  wire       [35:0]   _zz_7880;
  wire       [35:0]   _zz_7881;
  wire       [35:0]   _zz_7882;
  wire       [26:0]   _zz_7883;
  wire       [35:0]   _zz_7884;
  wire       [17:0]   _zz_7885;
  wire       [35:0]   _zz_7886;
  wire       [35:0]   _zz_7887;
  wire       [35:0]   _zz_7888;
  wire       [35:0]   _zz_7889;
  wire       [35:0]   _zz_7890;
  wire       [26:0]   _zz_7891;
  wire       [35:0]   _zz_7892;
  wire       [17:0]   _zz_7893;
  wire       [17:0]   _zz_7894;
  wire       [35:0]   _zz_7895;
  wire       [35:0]   _zz_7896;
  wire       [17:0]   _zz_7897;
  wire       [35:0]   _zz_7898;
  wire       [35:0]   _zz_7899;
  wire       [35:0]   _zz_7900;
  wire       [17:0]   _zz_7901;
  wire       [35:0]   _zz_7902;
  wire       [35:0]   _zz_7903;
  wire       [35:0]   _zz_7904;
  wire       [35:0]   _zz_7905;
  wire       [35:0]   _zz_7906;
  wire       [35:0]   _zz_7907;
  wire       [26:0]   _zz_7908;
  wire       [35:0]   _zz_7909;
  wire       [17:0]   _zz_7910;
  wire       [35:0]   _zz_7911;
  wire       [35:0]   _zz_7912;
  wire       [35:0]   _zz_7913;
  wire       [35:0]   _zz_7914;
  wire       [35:0]   _zz_7915;
  wire       [26:0]   _zz_7916;
  wire       [35:0]   _zz_7917;
  wire       [17:0]   _zz_7918;
  wire       [35:0]   _zz_7919;
  wire       [35:0]   _zz_7920;
  wire       [35:0]   _zz_7921;
  wire       [35:0]   _zz_7922;
  wire       [35:0]   _zz_7923;
  wire       [26:0]   _zz_7924;
  wire       [35:0]   _zz_7925;
  wire       [17:0]   _zz_7926;
  wire       [35:0]   _zz_7927;
  wire       [35:0]   _zz_7928;
  wire       [35:0]   _zz_7929;
  wire       [35:0]   _zz_7930;
  wire       [35:0]   _zz_7931;
  wire       [26:0]   _zz_7932;
  wire       [35:0]   _zz_7933;
  wire       [17:0]   _zz_7934;
  wire       [17:0]   _zz_7935;
  wire       [35:0]   _zz_7936;
  wire       [35:0]   _zz_7937;
  wire       [17:0]   _zz_7938;
  wire       [35:0]   _zz_7939;
  wire       [35:0]   _zz_7940;
  wire       [35:0]   _zz_7941;
  wire       [17:0]   _zz_7942;
  wire       [35:0]   _zz_7943;
  wire       [35:0]   _zz_7944;
  wire       [35:0]   _zz_7945;
  wire       [35:0]   _zz_7946;
  wire       [35:0]   _zz_7947;
  wire       [35:0]   _zz_7948;
  wire       [26:0]   _zz_7949;
  wire       [35:0]   _zz_7950;
  wire       [17:0]   _zz_7951;
  wire       [35:0]   _zz_7952;
  wire       [35:0]   _zz_7953;
  wire       [35:0]   _zz_7954;
  wire       [35:0]   _zz_7955;
  wire       [35:0]   _zz_7956;
  wire       [26:0]   _zz_7957;
  wire       [35:0]   _zz_7958;
  wire       [17:0]   _zz_7959;
  wire       [35:0]   _zz_7960;
  wire       [35:0]   _zz_7961;
  wire       [35:0]   _zz_7962;
  wire       [35:0]   _zz_7963;
  wire       [35:0]   _zz_7964;
  wire       [26:0]   _zz_7965;
  wire       [35:0]   _zz_7966;
  wire       [17:0]   _zz_7967;
  wire       [35:0]   _zz_7968;
  wire       [35:0]   _zz_7969;
  wire       [35:0]   _zz_7970;
  wire       [35:0]   _zz_7971;
  wire       [35:0]   _zz_7972;
  wire       [26:0]   _zz_7973;
  wire       [35:0]   _zz_7974;
  wire       [17:0]   _zz_7975;
  wire       [17:0]   _zz_7976;
  wire       [35:0]   _zz_7977;
  wire       [35:0]   _zz_7978;
  wire       [17:0]   _zz_7979;
  wire       [35:0]   _zz_7980;
  wire       [35:0]   _zz_7981;
  wire       [35:0]   _zz_7982;
  wire       [17:0]   _zz_7983;
  wire       [35:0]   _zz_7984;
  wire       [35:0]   _zz_7985;
  wire       [35:0]   _zz_7986;
  wire       [35:0]   _zz_7987;
  wire       [35:0]   _zz_7988;
  wire       [35:0]   _zz_7989;
  wire       [26:0]   _zz_7990;
  wire       [35:0]   _zz_7991;
  wire       [17:0]   _zz_7992;
  wire       [35:0]   _zz_7993;
  wire       [35:0]   _zz_7994;
  wire       [35:0]   _zz_7995;
  wire       [35:0]   _zz_7996;
  wire       [35:0]   _zz_7997;
  wire       [26:0]   _zz_7998;
  wire       [35:0]   _zz_7999;
  wire       [17:0]   _zz_8000;
  wire       [35:0]   _zz_8001;
  wire       [35:0]   _zz_8002;
  wire       [35:0]   _zz_8003;
  wire       [35:0]   _zz_8004;
  wire       [35:0]   _zz_8005;
  wire       [26:0]   _zz_8006;
  wire       [35:0]   _zz_8007;
  wire       [17:0]   _zz_8008;
  wire       [35:0]   _zz_8009;
  wire       [35:0]   _zz_8010;
  wire       [35:0]   _zz_8011;
  wire       [35:0]   _zz_8012;
  wire       [35:0]   _zz_8013;
  wire       [26:0]   _zz_8014;
  wire       [35:0]   _zz_8015;
  wire       [17:0]   _zz_8016;
  wire       [17:0]   _zz_8017;
  wire       [35:0]   _zz_8018;
  wire       [35:0]   _zz_8019;
  wire       [17:0]   _zz_8020;
  wire       [35:0]   _zz_8021;
  wire       [35:0]   _zz_8022;
  wire       [35:0]   _zz_8023;
  wire       [17:0]   _zz_8024;
  wire       [35:0]   _zz_8025;
  wire       [35:0]   _zz_8026;
  wire       [35:0]   _zz_8027;
  wire       [35:0]   _zz_8028;
  wire       [35:0]   _zz_8029;
  wire       [35:0]   _zz_8030;
  wire       [26:0]   _zz_8031;
  wire       [35:0]   _zz_8032;
  wire       [17:0]   _zz_8033;
  wire       [35:0]   _zz_8034;
  wire       [35:0]   _zz_8035;
  wire       [35:0]   _zz_8036;
  wire       [35:0]   _zz_8037;
  wire       [35:0]   _zz_8038;
  wire       [26:0]   _zz_8039;
  wire       [35:0]   _zz_8040;
  wire       [17:0]   _zz_8041;
  wire       [35:0]   _zz_8042;
  wire       [35:0]   _zz_8043;
  wire       [35:0]   _zz_8044;
  wire       [35:0]   _zz_8045;
  wire       [35:0]   _zz_8046;
  wire       [26:0]   _zz_8047;
  wire       [35:0]   _zz_8048;
  wire       [17:0]   _zz_8049;
  wire       [35:0]   _zz_8050;
  wire       [35:0]   _zz_8051;
  wire       [35:0]   _zz_8052;
  wire       [35:0]   _zz_8053;
  wire       [35:0]   _zz_8054;
  wire       [26:0]   _zz_8055;
  wire       [35:0]   _zz_8056;
  wire       [17:0]   _zz_8057;
  wire       [17:0]   _zz_8058;
  wire       [35:0]   _zz_8059;
  wire       [35:0]   _zz_8060;
  wire       [17:0]   _zz_8061;
  wire       [35:0]   _zz_8062;
  wire       [35:0]   _zz_8063;
  wire       [35:0]   _zz_8064;
  wire       [17:0]   _zz_8065;
  wire       [35:0]   _zz_8066;
  wire       [35:0]   _zz_8067;
  wire       [35:0]   _zz_8068;
  wire       [35:0]   _zz_8069;
  wire       [35:0]   _zz_8070;
  wire       [35:0]   _zz_8071;
  wire       [26:0]   _zz_8072;
  wire       [35:0]   _zz_8073;
  wire       [17:0]   _zz_8074;
  wire       [35:0]   _zz_8075;
  wire       [35:0]   _zz_8076;
  wire       [35:0]   _zz_8077;
  wire       [35:0]   _zz_8078;
  wire       [35:0]   _zz_8079;
  wire       [26:0]   _zz_8080;
  wire       [35:0]   _zz_8081;
  wire       [17:0]   _zz_8082;
  wire       [35:0]   _zz_8083;
  wire       [35:0]   _zz_8084;
  wire       [35:0]   _zz_8085;
  wire       [35:0]   _zz_8086;
  wire       [35:0]   _zz_8087;
  wire       [26:0]   _zz_8088;
  wire       [35:0]   _zz_8089;
  wire       [17:0]   _zz_8090;
  wire       [35:0]   _zz_8091;
  wire       [35:0]   _zz_8092;
  wire       [35:0]   _zz_8093;
  wire       [35:0]   _zz_8094;
  wire       [35:0]   _zz_8095;
  wire       [26:0]   _zz_8096;
  wire       [35:0]   _zz_8097;
  wire       [17:0]   _zz_8098;
  wire       [17:0]   _zz_8099;
  wire       [35:0]   _zz_8100;
  wire       [35:0]   _zz_8101;
  wire       [17:0]   _zz_8102;
  wire       [35:0]   _zz_8103;
  wire       [35:0]   _zz_8104;
  wire       [35:0]   _zz_8105;
  wire       [17:0]   _zz_8106;
  wire       [35:0]   _zz_8107;
  wire       [35:0]   _zz_8108;
  wire       [35:0]   _zz_8109;
  wire       [35:0]   _zz_8110;
  wire       [35:0]   _zz_8111;
  wire       [35:0]   _zz_8112;
  wire       [26:0]   _zz_8113;
  wire       [35:0]   _zz_8114;
  wire       [17:0]   _zz_8115;
  wire       [35:0]   _zz_8116;
  wire       [35:0]   _zz_8117;
  wire       [35:0]   _zz_8118;
  wire       [35:0]   _zz_8119;
  wire       [35:0]   _zz_8120;
  wire       [26:0]   _zz_8121;
  wire       [35:0]   _zz_8122;
  wire       [17:0]   _zz_8123;
  wire       [35:0]   _zz_8124;
  wire       [35:0]   _zz_8125;
  wire       [35:0]   _zz_8126;
  wire       [35:0]   _zz_8127;
  wire       [35:0]   _zz_8128;
  wire       [26:0]   _zz_8129;
  wire       [35:0]   _zz_8130;
  wire       [17:0]   _zz_8131;
  wire       [35:0]   _zz_8132;
  wire       [35:0]   _zz_8133;
  wire       [35:0]   _zz_8134;
  wire       [35:0]   _zz_8135;
  wire       [35:0]   _zz_8136;
  wire       [26:0]   _zz_8137;
  wire       [35:0]   _zz_8138;
  wire       [17:0]   _zz_8139;
  wire       [17:0]   _zz_8140;
  wire       [35:0]   _zz_8141;
  wire       [35:0]   _zz_8142;
  wire       [17:0]   _zz_8143;
  wire       [35:0]   _zz_8144;
  wire       [35:0]   _zz_8145;
  wire       [35:0]   _zz_8146;
  wire       [17:0]   _zz_8147;
  wire       [35:0]   _zz_8148;
  wire       [35:0]   _zz_8149;
  wire       [35:0]   _zz_8150;
  wire       [35:0]   _zz_8151;
  wire       [35:0]   _zz_8152;
  wire       [35:0]   _zz_8153;
  wire       [26:0]   _zz_8154;
  wire       [35:0]   _zz_8155;
  wire       [17:0]   _zz_8156;
  wire       [35:0]   _zz_8157;
  wire       [35:0]   _zz_8158;
  wire       [35:0]   _zz_8159;
  wire       [35:0]   _zz_8160;
  wire       [35:0]   _zz_8161;
  wire       [26:0]   _zz_8162;
  wire       [35:0]   _zz_8163;
  wire       [17:0]   _zz_8164;
  wire       [35:0]   _zz_8165;
  wire       [35:0]   _zz_8166;
  wire       [35:0]   _zz_8167;
  wire       [35:0]   _zz_8168;
  wire       [35:0]   _zz_8169;
  wire       [26:0]   _zz_8170;
  wire       [35:0]   _zz_8171;
  wire       [17:0]   _zz_8172;
  wire       [35:0]   _zz_8173;
  wire       [35:0]   _zz_8174;
  wire       [35:0]   _zz_8175;
  wire       [35:0]   _zz_8176;
  wire       [35:0]   _zz_8177;
  wire       [26:0]   _zz_8178;
  wire       [35:0]   _zz_8179;
  wire       [17:0]   _zz_8180;
  wire       [17:0]   _zz_8181;
  wire       [35:0]   _zz_8182;
  wire       [35:0]   _zz_8183;
  wire       [17:0]   _zz_8184;
  wire       [35:0]   _zz_8185;
  wire       [35:0]   _zz_8186;
  wire       [35:0]   _zz_8187;
  wire       [17:0]   _zz_8188;
  wire       [35:0]   _zz_8189;
  wire       [35:0]   _zz_8190;
  wire       [35:0]   _zz_8191;
  wire       [35:0]   _zz_8192;
  wire       [35:0]   _zz_8193;
  wire       [35:0]   _zz_8194;
  wire       [26:0]   _zz_8195;
  wire       [35:0]   _zz_8196;
  wire       [17:0]   _zz_8197;
  wire       [35:0]   _zz_8198;
  wire       [35:0]   _zz_8199;
  wire       [35:0]   _zz_8200;
  wire       [35:0]   _zz_8201;
  wire       [35:0]   _zz_8202;
  wire       [26:0]   _zz_8203;
  wire       [35:0]   _zz_8204;
  wire       [17:0]   _zz_8205;
  wire       [35:0]   _zz_8206;
  wire       [35:0]   _zz_8207;
  wire       [35:0]   _zz_8208;
  wire       [35:0]   _zz_8209;
  wire       [35:0]   _zz_8210;
  wire       [26:0]   _zz_8211;
  wire       [35:0]   _zz_8212;
  wire       [17:0]   _zz_8213;
  wire       [35:0]   _zz_8214;
  wire       [35:0]   _zz_8215;
  wire       [35:0]   _zz_8216;
  wire       [35:0]   _zz_8217;
  wire       [35:0]   _zz_8218;
  wire       [26:0]   _zz_8219;
  wire       [35:0]   _zz_8220;
  wire       [17:0]   _zz_8221;
  wire       [17:0]   _zz_8222;
  wire       [35:0]   _zz_8223;
  wire       [35:0]   _zz_8224;
  wire       [17:0]   _zz_8225;
  wire       [35:0]   _zz_8226;
  wire       [35:0]   _zz_8227;
  wire       [35:0]   _zz_8228;
  wire       [17:0]   _zz_8229;
  wire       [35:0]   _zz_8230;
  wire       [35:0]   _zz_8231;
  wire       [35:0]   _zz_8232;
  wire       [35:0]   _zz_8233;
  wire       [35:0]   _zz_8234;
  wire       [35:0]   _zz_8235;
  wire       [26:0]   _zz_8236;
  wire       [35:0]   _zz_8237;
  wire       [17:0]   _zz_8238;
  wire       [35:0]   _zz_8239;
  wire       [35:0]   _zz_8240;
  wire       [35:0]   _zz_8241;
  wire       [35:0]   _zz_8242;
  wire       [35:0]   _zz_8243;
  wire       [26:0]   _zz_8244;
  wire       [35:0]   _zz_8245;
  wire       [17:0]   _zz_8246;
  wire       [35:0]   _zz_8247;
  wire       [35:0]   _zz_8248;
  wire       [35:0]   _zz_8249;
  wire       [35:0]   _zz_8250;
  wire       [35:0]   _zz_8251;
  wire       [26:0]   _zz_8252;
  wire       [35:0]   _zz_8253;
  wire       [17:0]   _zz_8254;
  wire       [35:0]   _zz_8255;
  wire       [35:0]   _zz_8256;
  wire       [35:0]   _zz_8257;
  wire       [35:0]   _zz_8258;
  wire       [35:0]   _zz_8259;
  wire       [26:0]   _zz_8260;
  wire       [35:0]   _zz_8261;
  wire       [17:0]   _zz_8262;
  wire       [17:0]   _zz_8263;
  wire       [35:0]   _zz_8264;
  wire       [35:0]   _zz_8265;
  wire       [17:0]   _zz_8266;
  wire       [35:0]   _zz_8267;
  wire       [35:0]   _zz_8268;
  wire       [35:0]   _zz_8269;
  wire       [17:0]   _zz_8270;
  wire       [35:0]   _zz_8271;
  wire       [35:0]   _zz_8272;
  wire       [35:0]   _zz_8273;
  wire       [35:0]   _zz_8274;
  wire       [35:0]   _zz_8275;
  wire       [35:0]   _zz_8276;
  wire       [26:0]   _zz_8277;
  wire       [35:0]   _zz_8278;
  wire       [17:0]   _zz_8279;
  wire       [35:0]   _zz_8280;
  wire       [35:0]   _zz_8281;
  wire       [35:0]   _zz_8282;
  wire       [35:0]   _zz_8283;
  wire       [35:0]   _zz_8284;
  wire       [26:0]   _zz_8285;
  wire       [35:0]   _zz_8286;
  wire       [17:0]   _zz_8287;
  wire       [35:0]   _zz_8288;
  wire       [35:0]   _zz_8289;
  wire       [35:0]   _zz_8290;
  wire       [35:0]   _zz_8291;
  wire       [35:0]   _zz_8292;
  wire       [26:0]   _zz_8293;
  wire       [35:0]   _zz_8294;
  wire       [17:0]   _zz_8295;
  wire       [35:0]   _zz_8296;
  wire       [35:0]   _zz_8297;
  wire       [35:0]   _zz_8298;
  wire       [35:0]   _zz_8299;
  wire       [35:0]   _zz_8300;
  wire       [26:0]   _zz_8301;
  wire       [35:0]   _zz_8302;
  wire       [17:0]   _zz_8303;
  wire       [17:0]   _zz_8304;
  wire       [35:0]   _zz_8305;
  wire       [35:0]   _zz_8306;
  wire       [17:0]   _zz_8307;
  wire       [35:0]   _zz_8308;
  wire       [35:0]   _zz_8309;
  wire       [35:0]   _zz_8310;
  wire       [17:0]   _zz_8311;
  wire       [35:0]   _zz_8312;
  wire       [35:0]   _zz_8313;
  wire       [35:0]   _zz_8314;
  wire       [35:0]   _zz_8315;
  wire       [35:0]   _zz_8316;
  wire       [35:0]   _zz_8317;
  wire       [26:0]   _zz_8318;
  wire       [35:0]   _zz_8319;
  wire       [17:0]   _zz_8320;
  wire       [35:0]   _zz_8321;
  wire       [35:0]   _zz_8322;
  wire       [35:0]   _zz_8323;
  wire       [35:0]   _zz_8324;
  wire       [35:0]   _zz_8325;
  wire       [26:0]   _zz_8326;
  wire       [35:0]   _zz_8327;
  wire       [17:0]   _zz_8328;
  wire       [35:0]   _zz_8329;
  wire       [35:0]   _zz_8330;
  wire       [35:0]   _zz_8331;
  wire       [35:0]   _zz_8332;
  wire       [35:0]   _zz_8333;
  wire       [26:0]   _zz_8334;
  wire       [35:0]   _zz_8335;
  wire       [17:0]   _zz_8336;
  wire       [35:0]   _zz_8337;
  wire       [35:0]   _zz_8338;
  wire       [35:0]   _zz_8339;
  wire       [35:0]   _zz_8340;
  wire       [35:0]   _zz_8341;
  wire       [26:0]   _zz_8342;
  wire       [35:0]   _zz_8343;
  wire       [17:0]   _zz_8344;
  wire       [17:0]   _zz_8345;
  wire       [35:0]   _zz_8346;
  wire       [35:0]   _zz_8347;
  wire       [17:0]   _zz_8348;
  wire       [35:0]   _zz_8349;
  wire       [35:0]   _zz_8350;
  wire       [35:0]   _zz_8351;
  wire       [17:0]   _zz_8352;
  wire       [35:0]   _zz_8353;
  wire       [35:0]   _zz_8354;
  wire       [35:0]   _zz_8355;
  wire       [35:0]   _zz_8356;
  wire       [35:0]   _zz_8357;
  wire       [35:0]   _zz_8358;
  wire       [26:0]   _zz_8359;
  wire       [35:0]   _zz_8360;
  wire       [17:0]   _zz_8361;
  wire       [35:0]   _zz_8362;
  wire       [35:0]   _zz_8363;
  wire       [35:0]   _zz_8364;
  wire       [35:0]   _zz_8365;
  wire       [35:0]   _zz_8366;
  wire       [26:0]   _zz_8367;
  wire       [35:0]   _zz_8368;
  wire       [17:0]   _zz_8369;
  wire       [35:0]   _zz_8370;
  wire       [35:0]   _zz_8371;
  wire       [35:0]   _zz_8372;
  wire       [35:0]   _zz_8373;
  wire       [35:0]   _zz_8374;
  wire       [26:0]   _zz_8375;
  wire       [35:0]   _zz_8376;
  wire       [17:0]   _zz_8377;
  wire       [35:0]   _zz_8378;
  wire       [35:0]   _zz_8379;
  wire       [35:0]   _zz_8380;
  wire       [35:0]   _zz_8381;
  wire       [35:0]   _zz_8382;
  wire       [26:0]   _zz_8383;
  wire       [35:0]   _zz_8384;
  wire       [17:0]   _zz_8385;
  wire       [17:0]   _zz_8386;
  wire       [35:0]   _zz_8387;
  wire       [35:0]   _zz_8388;
  wire       [17:0]   _zz_8389;
  wire       [35:0]   _zz_8390;
  wire       [35:0]   _zz_8391;
  wire       [35:0]   _zz_8392;
  wire       [17:0]   _zz_8393;
  wire       [35:0]   _zz_8394;
  wire       [35:0]   _zz_8395;
  wire       [35:0]   _zz_8396;
  wire       [35:0]   _zz_8397;
  wire       [35:0]   _zz_8398;
  wire       [35:0]   _zz_8399;
  wire       [26:0]   _zz_8400;
  wire       [35:0]   _zz_8401;
  wire       [17:0]   _zz_8402;
  wire       [35:0]   _zz_8403;
  wire       [35:0]   _zz_8404;
  wire       [35:0]   _zz_8405;
  wire       [35:0]   _zz_8406;
  wire       [35:0]   _zz_8407;
  wire       [26:0]   _zz_8408;
  wire       [35:0]   _zz_8409;
  wire       [17:0]   _zz_8410;
  wire       [35:0]   _zz_8411;
  wire       [35:0]   _zz_8412;
  wire       [35:0]   _zz_8413;
  wire       [35:0]   _zz_8414;
  wire       [35:0]   _zz_8415;
  wire       [26:0]   _zz_8416;
  wire       [35:0]   _zz_8417;
  wire       [17:0]   _zz_8418;
  wire       [35:0]   _zz_8419;
  wire       [35:0]   _zz_8420;
  wire       [35:0]   _zz_8421;
  wire       [35:0]   _zz_8422;
  wire       [35:0]   _zz_8423;
  wire       [26:0]   _zz_8424;
  wire       [35:0]   _zz_8425;
  wire       [17:0]   _zz_8426;
  wire       [17:0]   _zz_8427;
  wire       [35:0]   _zz_8428;
  wire       [35:0]   _zz_8429;
  wire       [17:0]   _zz_8430;
  wire       [35:0]   _zz_8431;
  wire       [35:0]   _zz_8432;
  wire       [35:0]   _zz_8433;
  wire       [17:0]   _zz_8434;
  wire       [35:0]   _zz_8435;
  wire       [35:0]   _zz_8436;
  wire       [35:0]   _zz_8437;
  wire       [35:0]   _zz_8438;
  wire       [35:0]   _zz_8439;
  wire       [35:0]   _zz_8440;
  wire       [26:0]   _zz_8441;
  wire       [35:0]   _zz_8442;
  wire       [17:0]   _zz_8443;
  wire       [35:0]   _zz_8444;
  wire       [35:0]   _zz_8445;
  wire       [35:0]   _zz_8446;
  wire       [35:0]   _zz_8447;
  wire       [35:0]   _zz_8448;
  wire       [26:0]   _zz_8449;
  wire       [35:0]   _zz_8450;
  wire       [17:0]   _zz_8451;
  wire       [35:0]   _zz_8452;
  wire       [35:0]   _zz_8453;
  wire       [35:0]   _zz_8454;
  wire       [35:0]   _zz_8455;
  wire       [35:0]   _zz_8456;
  wire       [26:0]   _zz_8457;
  wire       [35:0]   _zz_8458;
  wire       [17:0]   _zz_8459;
  wire       [35:0]   _zz_8460;
  wire       [35:0]   _zz_8461;
  wire       [35:0]   _zz_8462;
  wire       [35:0]   _zz_8463;
  wire       [35:0]   _zz_8464;
  wire       [26:0]   _zz_8465;
  wire       [35:0]   _zz_8466;
  wire       [17:0]   _zz_8467;
  wire       [17:0]   _zz_8468;
  wire       [35:0]   _zz_8469;
  wire       [35:0]   _zz_8470;
  wire       [17:0]   _zz_8471;
  wire       [35:0]   _zz_8472;
  wire       [35:0]   _zz_8473;
  wire       [35:0]   _zz_8474;
  wire       [17:0]   _zz_8475;
  wire       [35:0]   _zz_8476;
  wire       [35:0]   _zz_8477;
  wire       [35:0]   _zz_8478;
  wire       [35:0]   _zz_8479;
  wire       [35:0]   _zz_8480;
  wire       [35:0]   _zz_8481;
  wire       [26:0]   _zz_8482;
  wire       [35:0]   _zz_8483;
  wire       [17:0]   _zz_8484;
  wire       [35:0]   _zz_8485;
  wire       [35:0]   _zz_8486;
  wire       [35:0]   _zz_8487;
  wire       [35:0]   _zz_8488;
  wire       [35:0]   _zz_8489;
  wire       [26:0]   _zz_8490;
  wire       [35:0]   _zz_8491;
  wire       [17:0]   _zz_8492;
  wire       [35:0]   _zz_8493;
  wire       [35:0]   _zz_8494;
  wire       [35:0]   _zz_8495;
  wire       [35:0]   _zz_8496;
  wire       [35:0]   _zz_8497;
  wire       [26:0]   _zz_8498;
  wire       [35:0]   _zz_8499;
  wire       [17:0]   _zz_8500;
  wire       [35:0]   _zz_8501;
  wire       [35:0]   _zz_8502;
  wire       [35:0]   _zz_8503;
  wire       [35:0]   _zz_8504;
  wire       [35:0]   _zz_8505;
  wire       [26:0]   _zz_8506;
  wire       [35:0]   _zz_8507;
  wire       [17:0]   _zz_8508;
  wire       [17:0]   _zz_8509;
  wire       [35:0]   _zz_8510;
  wire       [35:0]   _zz_8511;
  wire       [17:0]   _zz_8512;
  wire       [35:0]   _zz_8513;
  wire       [35:0]   _zz_8514;
  wire       [35:0]   _zz_8515;
  wire       [17:0]   _zz_8516;
  wire       [35:0]   _zz_8517;
  wire       [35:0]   _zz_8518;
  wire       [35:0]   _zz_8519;
  wire       [35:0]   _zz_8520;
  wire       [35:0]   _zz_8521;
  wire       [35:0]   _zz_8522;
  wire       [26:0]   _zz_8523;
  wire       [35:0]   _zz_8524;
  wire       [17:0]   _zz_8525;
  wire       [35:0]   _zz_8526;
  wire       [35:0]   _zz_8527;
  wire       [35:0]   _zz_8528;
  wire       [35:0]   _zz_8529;
  wire       [35:0]   _zz_8530;
  wire       [26:0]   _zz_8531;
  wire       [35:0]   _zz_8532;
  wire       [17:0]   _zz_8533;
  wire       [35:0]   _zz_8534;
  wire       [35:0]   _zz_8535;
  wire       [35:0]   _zz_8536;
  wire       [35:0]   _zz_8537;
  wire       [35:0]   _zz_8538;
  wire       [26:0]   _zz_8539;
  wire       [35:0]   _zz_8540;
  wire       [17:0]   _zz_8541;
  wire       [35:0]   _zz_8542;
  wire       [35:0]   _zz_8543;
  wire       [35:0]   _zz_8544;
  wire       [35:0]   _zz_8545;
  wire       [35:0]   _zz_8546;
  wire       [26:0]   _zz_8547;
  wire       [35:0]   _zz_8548;
  wire       [17:0]   _zz_8549;
  wire       [17:0]   _zz_8550;
  wire       [35:0]   _zz_8551;
  wire       [35:0]   _zz_8552;
  wire       [17:0]   _zz_8553;
  wire       [35:0]   _zz_8554;
  wire       [35:0]   _zz_8555;
  wire       [35:0]   _zz_8556;
  wire       [17:0]   _zz_8557;
  wire       [35:0]   _zz_8558;
  wire       [35:0]   _zz_8559;
  wire       [35:0]   _zz_8560;
  wire       [35:0]   _zz_8561;
  wire       [35:0]   _zz_8562;
  wire       [35:0]   _zz_8563;
  wire       [26:0]   _zz_8564;
  wire       [35:0]   _zz_8565;
  wire       [17:0]   _zz_8566;
  wire       [35:0]   _zz_8567;
  wire       [35:0]   _zz_8568;
  wire       [35:0]   _zz_8569;
  wire       [35:0]   _zz_8570;
  wire       [35:0]   _zz_8571;
  wire       [26:0]   _zz_8572;
  wire       [35:0]   _zz_8573;
  wire       [17:0]   _zz_8574;
  wire       [35:0]   _zz_8575;
  wire       [35:0]   _zz_8576;
  wire       [35:0]   _zz_8577;
  wire       [35:0]   _zz_8578;
  wire       [35:0]   _zz_8579;
  wire       [26:0]   _zz_8580;
  wire       [35:0]   _zz_8581;
  wire       [17:0]   _zz_8582;
  wire       [35:0]   _zz_8583;
  wire       [35:0]   _zz_8584;
  wire       [35:0]   _zz_8585;
  wire       [35:0]   _zz_8586;
  wire       [35:0]   _zz_8587;
  wire       [26:0]   _zz_8588;
  wire       [35:0]   _zz_8589;
  wire       [17:0]   _zz_8590;
  wire       [17:0]   _zz_8591;
  wire       [35:0]   _zz_8592;
  wire       [35:0]   _zz_8593;
  wire       [17:0]   _zz_8594;
  wire       [35:0]   _zz_8595;
  wire       [35:0]   _zz_8596;
  wire       [35:0]   _zz_8597;
  wire       [17:0]   _zz_8598;
  wire       [35:0]   _zz_8599;
  wire       [35:0]   _zz_8600;
  wire       [35:0]   _zz_8601;
  wire       [35:0]   _zz_8602;
  wire       [35:0]   _zz_8603;
  wire       [35:0]   _zz_8604;
  wire       [26:0]   _zz_8605;
  wire       [35:0]   _zz_8606;
  wire       [17:0]   _zz_8607;
  wire       [35:0]   _zz_8608;
  wire       [35:0]   _zz_8609;
  wire       [35:0]   _zz_8610;
  wire       [35:0]   _zz_8611;
  wire       [35:0]   _zz_8612;
  wire       [26:0]   _zz_8613;
  wire       [35:0]   _zz_8614;
  wire       [17:0]   _zz_8615;
  wire       [35:0]   _zz_8616;
  wire       [35:0]   _zz_8617;
  wire       [35:0]   _zz_8618;
  wire       [35:0]   _zz_8619;
  wire       [35:0]   _zz_8620;
  wire       [26:0]   _zz_8621;
  wire       [35:0]   _zz_8622;
  wire       [17:0]   _zz_8623;
  wire       [35:0]   _zz_8624;
  wire       [35:0]   _zz_8625;
  wire       [35:0]   _zz_8626;
  wire       [35:0]   _zz_8627;
  wire       [35:0]   _zz_8628;
  wire       [26:0]   _zz_8629;
  wire       [35:0]   _zz_8630;
  wire       [17:0]   _zz_8631;
  wire       [17:0]   _zz_8632;
  wire       [35:0]   _zz_8633;
  wire       [35:0]   _zz_8634;
  wire       [17:0]   _zz_8635;
  wire       [35:0]   _zz_8636;
  wire       [35:0]   _zz_8637;
  wire       [35:0]   _zz_8638;
  wire       [17:0]   _zz_8639;
  wire       [35:0]   _zz_8640;
  wire       [35:0]   _zz_8641;
  wire       [35:0]   _zz_8642;
  wire       [35:0]   _zz_8643;
  wire       [35:0]   _zz_8644;
  wire       [35:0]   _zz_8645;
  wire       [26:0]   _zz_8646;
  wire       [35:0]   _zz_8647;
  wire       [17:0]   _zz_8648;
  wire       [35:0]   _zz_8649;
  wire       [35:0]   _zz_8650;
  wire       [35:0]   _zz_8651;
  wire       [35:0]   _zz_8652;
  wire       [35:0]   _zz_8653;
  wire       [26:0]   _zz_8654;
  wire       [35:0]   _zz_8655;
  wire       [17:0]   _zz_8656;
  wire       [35:0]   _zz_8657;
  wire       [35:0]   _zz_8658;
  wire       [35:0]   _zz_8659;
  wire       [35:0]   _zz_8660;
  wire       [35:0]   _zz_8661;
  wire       [26:0]   _zz_8662;
  wire       [35:0]   _zz_8663;
  wire       [17:0]   _zz_8664;
  wire       [35:0]   _zz_8665;
  wire       [35:0]   _zz_8666;
  wire       [35:0]   _zz_8667;
  wire       [35:0]   _zz_8668;
  wire       [35:0]   _zz_8669;
  wire       [26:0]   _zz_8670;
  wire       [35:0]   _zz_8671;
  wire       [17:0]   _zz_8672;
  wire       [17:0]   _zz_8673;
  wire       [35:0]   _zz_8674;
  wire       [35:0]   _zz_8675;
  wire       [17:0]   _zz_8676;
  wire       [35:0]   _zz_8677;
  wire       [35:0]   _zz_8678;
  wire       [35:0]   _zz_8679;
  wire       [17:0]   _zz_8680;
  wire       [35:0]   _zz_8681;
  wire       [35:0]   _zz_8682;
  wire       [35:0]   _zz_8683;
  wire       [35:0]   _zz_8684;
  wire       [35:0]   _zz_8685;
  wire       [35:0]   _zz_8686;
  wire       [26:0]   _zz_8687;
  wire       [35:0]   _zz_8688;
  wire       [17:0]   _zz_8689;
  wire       [35:0]   _zz_8690;
  wire       [35:0]   _zz_8691;
  wire       [35:0]   _zz_8692;
  wire       [35:0]   _zz_8693;
  wire       [35:0]   _zz_8694;
  wire       [26:0]   _zz_8695;
  wire       [35:0]   _zz_8696;
  wire       [17:0]   _zz_8697;
  wire       [35:0]   _zz_8698;
  wire       [35:0]   _zz_8699;
  wire       [35:0]   _zz_8700;
  wire       [35:0]   _zz_8701;
  wire       [35:0]   _zz_8702;
  wire       [26:0]   _zz_8703;
  wire       [35:0]   _zz_8704;
  wire       [17:0]   _zz_8705;
  wire       [35:0]   _zz_8706;
  wire       [35:0]   _zz_8707;
  wire       [35:0]   _zz_8708;
  wire       [35:0]   _zz_8709;
  wire       [35:0]   _zz_8710;
  wire       [26:0]   _zz_8711;
  wire       [35:0]   _zz_8712;
  wire       [17:0]   _zz_8713;
  wire       [17:0]   _zz_8714;
  wire       [35:0]   _zz_8715;
  wire       [35:0]   _zz_8716;
  wire       [17:0]   _zz_8717;
  wire       [35:0]   _zz_8718;
  wire       [35:0]   _zz_8719;
  wire       [35:0]   _zz_8720;
  wire       [17:0]   _zz_8721;
  wire       [35:0]   _zz_8722;
  wire       [35:0]   _zz_8723;
  wire       [35:0]   _zz_8724;
  wire       [35:0]   _zz_8725;
  wire       [35:0]   _zz_8726;
  wire       [35:0]   _zz_8727;
  wire       [26:0]   _zz_8728;
  wire       [35:0]   _zz_8729;
  wire       [17:0]   _zz_8730;
  wire       [35:0]   _zz_8731;
  wire       [35:0]   _zz_8732;
  wire       [35:0]   _zz_8733;
  wire       [35:0]   _zz_8734;
  wire       [35:0]   _zz_8735;
  wire       [26:0]   _zz_8736;
  wire       [35:0]   _zz_8737;
  wire       [17:0]   _zz_8738;
  wire       [35:0]   _zz_8739;
  wire       [35:0]   _zz_8740;
  wire       [35:0]   _zz_8741;
  wire       [35:0]   _zz_8742;
  wire       [35:0]   _zz_8743;
  wire       [26:0]   _zz_8744;
  wire       [35:0]   _zz_8745;
  wire       [17:0]   _zz_8746;
  wire       [35:0]   _zz_8747;
  wire       [35:0]   _zz_8748;
  wire       [35:0]   _zz_8749;
  wire       [35:0]   _zz_8750;
  wire       [35:0]   _zz_8751;
  wire       [26:0]   _zz_8752;
  wire       [35:0]   _zz_8753;
  wire       [17:0]   _zz_8754;
  wire       [17:0]   _zz_8755;
  wire       [35:0]   _zz_8756;
  wire       [35:0]   _zz_8757;
  wire       [17:0]   _zz_8758;
  wire       [35:0]   _zz_8759;
  wire       [35:0]   _zz_8760;
  wire       [35:0]   _zz_8761;
  wire       [17:0]   _zz_8762;
  wire       [35:0]   _zz_8763;
  wire       [35:0]   _zz_8764;
  wire       [35:0]   _zz_8765;
  wire       [35:0]   _zz_8766;
  wire       [35:0]   _zz_8767;
  wire       [35:0]   _zz_8768;
  wire       [26:0]   _zz_8769;
  wire       [35:0]   _zz_8770;
  wire       [17:0]   _zz_8771;
  wire       [35:0]   _zz_8772;
  wire       [35:0]   _zz_8773;
  wire       [35:0]   _zz_8774;
  wire       [35:0]   _zz_8775;
  wire       [35:0]   _zz_8776;
  wire       [26:0]   _zz_8777;
  wire       [35:0]   _zz_8778;
  wire       [17:0]   _zz_8779;
  wire       [35:0]   _zz_8780;
  wire       [35:0]   _zz_8781;
  wire       [35:0]   _zz_8782;
  wire       [35:0]   _zz_8783;
  wire       [35:0]   _zz_8784;
  wire       [26:0]   _zz_8785;
  wire       [35:0]   _zz_8786;
  wire       [17:0]   _zz_8787;
  wire       [35:0]   _zz_8788;
  wire       [35:0]   _zz_8789;
  wire       [35:0]   _zz_8790;
  wire       [35:0]   _zz_8791;
  wire       [35:0]   _zz_8792;
  wire       [26:0]   _zz_8793;
  wire       [35:0]   _zz_8794;
  wire       [17:0]   _zz_8795;
  wire       [17:0]   _zz_8796;
  wire       [35:0]   _zz_8797;
  wire       [35:0]   _zz_8798;
  wire       [17:0]   _zz_8799;
  wire       [35:0]   _zz_8800;
  wire       [35:0]   _zz_8801;
  wire       [35:0]   _zz_8802;
  wire       [17:0]   _zz_8803;
  wire       [35:0]   _zz_8804;
  wire       [35:0]   _zz_8805;
  wire       [35:0]   _zz_8806;
  wire       [35:0]   _zz_8807;
  wire       [35:0]   _zz_8808;
  wire       [35:0]   _zz_8809;
  wire       [26:0]   _zz_8810;
  wire       [35:0]   _zz_8811;
  wire       [17:0]   _zz_8812;
  wire       [35:0]   _zz_8813;
  wire       [35:0]   _zz_8814;
  wire       [35:0]   _zz_8815;
  wire       [35:0]   _zz_8816;
  wire       [35:0]   _zz_8817;
  wire       [26:0]   _zz_8818;
  wire       [35:0]   _zz_8819;
  wire       [17:0]   _zz_8820;
  wire       [35:0]   _zz_8821;
  wire       [35:0]   _zz_8822;
  wire       [35:0]   _zz_8823;
  wire       [35:0]   _zz_8824;
  wire       [35:0]   _zz_8825;
  wire       [26:0]   _zz_8826;
  wire       [35:0]   _zz_8827;
  wire       [17:0]   _zz_8828;
  wire       [35:0]   _zz_8829;
  wire       [35:0]   _zz_8830;
  wire       [35:0]   _zz_8831;
  wire       [35:0]   _zz_8832;
  wire       [35:0]   _zz_8833;
  wire       [26:0]   _zz_8834;
  wire       [35:0]   _zz_8835;
  wire       [17:0]   _zz_8836;
  wire       [17:0]   _zz_8837;
  wire       [35:0]   _zz_8838;
  wire       [35:0]   _zz_8839;
  wire       [17:0]   _zz_8840;
  wire       [35:0]   _zz_8841;
  wire       [35:0]   _zz_8842;
  wire       [35:0]   _zz_8843;
  wire       [17:0]   _zz_8844;
  wire       [35:0]   _zz_8845;
  wire       [35:0]   _zz_8846;
  wire       [35:0]   _zz_8847;
  wire       [35:0]   _zz_8848;
  wire       [35:0]   _zz_8849;
  wire       [35:0]   _zz_8850;
  wire       [26:0]   _zz_8851;
  wire       [35:0]   _zz_8852;
  wire       [17:0]   _zz_8853;
  wire       [35:0]   _zz_8854;
  wire       [35:0]   _zz_8855;
  wire       [35:0]   _zz_8856;
  wire       [35:0]   _zz_8857;
  wire       [35:0]   _zz_8858;
  wire       [26:0]   _zz_8859;
  wire       [35:0]   _zz_8860;
  wire       [17:0]   _zz_8861;
  wire       [35:0]   _zz_8862;
  wire       [35:0]   _zz_8863;
  wire       [35:0]   _zz_8864;
  wire       [35:0]   _zz_8865;
  wire       [35:0]   _zz_8866;
  wire       [26:0]   _zz_8867;
  wire       [35:0]   _zz_8868;
  wire       [17:0]   _zz_8869;
  wire       [35:0]   _zz_8870;
  wire       [35:0]   _zz_8871;
  wire       [35:0]   _zz_8872;
  wire       [35:0]   _zz_8873;
  wire       [35:0]   _zz_8874;
  wire       [26:0]   _zz_8875;
  wire       [35:0]   _zz_8876;
  wire       [17:0]   _zz_8877;
  wire       [17:0]   _zz_8878;
  wire       [35:0]   _zz_8879;
  wire       [35:0]   _zz_8880;
  wire       [17:0]   _zz_8881;
  wire       [35:0]   _zz_8882;
  wire       [35:0]   _zz_8883;
  wire       [35:0]   _zz_8884;
  wire       [17:0]   _zz_8885;
  wire       [35:0]   _zz_8886;
  wire       [35:0]   _zz_8887;
  wire       [35:0]   _zz_8888;
  wire       [35:0]   _zz_8889;
  wire       [35:0]   _zz_8890;
  wire       [35:0]   _zz_8891;
  wire       [26:0]   _zz_8892;
  wire       [35:0]   _zz_8893;
  wire       [17:0]   _zz_8894;
  wire       [35:0]   _zz_8895;
  wire       [35:0]   _zz_8896;
  wire       [35:0]   _zz_8897;
  wire       [35:0]   _zz_8898;
  wire       [35:0]   _zz_8899;
  wire       [26:0]   _zz_8900;
  wire       [35:0]   _zz_8901;
  wire       [17:0]   _zz_8902;
  wire       [35:0]   _zz_8903;
  wire       [35:0]   _zz_8904;
  wire       [35:0]   _zz_8905;
  wire       [35:0]   _zz_8906;
  wire       [35:0]   _zz_8907;
  wire       [26:0]   _zz_8908;
  wire       [35:0]   _zz_8909;
  wire       [17:0]   _zz_8910;
  wire       [35:0]   _zz_8911;
  wire       [35:0]   _zz_8912;
  wire       [35:0]   _zz_8913;
  wire       [35:0]   _zz_8914;
  wire       [35:0]   _zz_8915;
  wire       [26:0]   _zz_8916;
  wire       [35:0]   _zz_8917;
  wire       [17:0]   _zz_8918;
  wire       [17:0]   _zz_8919;
  wire       [35:0]   _zz_8920;
  wire       [35:0]   _zz_8921;
  wire       [17:0]   _zz_8922;
  wire       [35:0]   _zz_8923;
  wire       [35:0]   _zz_8924;
  wire       [35:0]   _zz_8925;
  wire       [17:0]   _zz_8926;
  wire       [35:0]   _zz_8927;
  wire       [35:0]   _zz_8928;
  wire       [35:0]   _zz_8929;
  wire       [35:0]   _zz_8930;
  wire       [35:0]   _zz_8931;
  wire       [35:0]   _zz_8932;
  wire       [26:0]   _zz_8933;
  wire       [35:0]   _zz_8934;
  wire       [17:0]   _zz_8935;
  wire       [35:0]   _zz_8936;
  wire       [35:0]   _zz_8937;
  wire       [35:0]   _zz_8938;
  wire       [35:0]   _zz_8939;
  wire       [35:0]   _zz_8940;
  wire       [26:0]   _zz_8941;
  wire       [35:0]   _zz_8942;
  wire       [17:0]   _zz_8943;
  wire       [35:0]   _zz_8944;
  wire       [35:0]   _zz_8945;
  wire       [35:0]   _zz_8946;
  wire       [35:0]   _zz_8947;
  wire       [35:0]   _zz_8948;
  wire       [26:0]   _zz_8949;
  wire       [35:0]   _zz_8950;
  wire       [17:0]   _zz_8951;
  wire       [35:0]   _zz_8952;
  wire       [35:0]   _zz_8953;
  wire       [35:0]   _zz_8954;
  wire       [35:0]   _zz_8955;
  wire       [35:0]   _zz_8956;
  wire       [26:0]   _zz_8957;
  wire       [35:0]   _zz_8958;
  wire       [17:0]   _zz_8959;
  wire       [17:0]   _zz_8960;
  wire       [35:0]   _zz_8961;
  wire       [35:0]   _zz_8962;
  wire       [17:0]   _zz_8963;
  wire       [35:0]   _zz_8964;
  wire       [35:0]   _zz_8965;
  wire       [35:0]   _zz_8966;
  wire       [17:0]   _zz_8967;
  wire       [35:0]   _zz_8968;
  wire       [35:0]   _zz_8969;
  wire       [35:0]   _zz_8970;
  wire       [35:0]   _zz_8971;
  wire       [35:0]   _zz_8972;
  wire       [35:0]   _zz_8973;
  wire       [26:0]   _zz_8974;
  wire       [35:0]   _zz_8975;
  wire       [17:0]   _zz_8976;
  wire       [35:0]   _zz_8977;
  wire       [35:0]   _zz_8978;
  wire       [35:0]   _zz_8979;
  wire       [35:0]   _zz_8980;
  wire       [35:0]   _zz_8981;
  wire       [26:0]   _zz_8982;
  wire       [35:0]   _zz_8983;
  wire       [17:0]   _zz_8984;
  wire       [35:0]   _zz_8985;
  wire       [35:0]   _zz_8986;
  wire       [35:0]   _zz_8987;
  wire       [35:0]   _zz_8988;
  wire       [35:0]   _zz_8989;
  wire       [26:0]   _zz_8990;
  wire       [35:0]   _zz_8991;
  wire       [17:0]   _zz_8992;
  wire       [35:0]   _zz_8993;
  wire       [35:0]   _zz_8994;
  wire       [35:0]   _zz_8995;
  wire       [35:0]   _zz_8996;
  wire       [35:0]   _zz_8997;
  wire       [26:0]   _zz_8998;
  wire       [35:0]   _zz_8999;
  wire       [17:0]   _zz_9000;
  wire       [17:0]   _zz_9001;
  wire       [35:0]   _zz_9002;
  wire       [35:0]   _zz_9003;
  wire       [17:0]   _zz_9004;
  wire       [35:0]   _zz_9005;
  wire       [35:0]   _zz_9006;
  wire       [35:0]   _zz_9007;
  wire       [17:0]   _zz_9008;
  wire       [35:0]   _zz_9009;
  wire       [35:0]   _zz_9010;
  wire       [35:0]   _zz_9011;
  wire       [35:0]   _zz_9012;
  wire       [35:0]   _zz_9013;
  wire       [35:0]   _zz_9014;
  wire       [26:0]   _zz_9015;
  wire       [35:0]   _zz_9016;
  wire       [17:0]   _zz_9017;
  wire       [35:0]   _zz_9018;
  wire       [35:0]   _zz_9019;
  wire       [35:0]   _zz_9020;
  wire       [35:0]   _zz_9021;
  wire       [35:0]   _zz_9022;
  wire       [26:0]   _zz_9023;
  wire       [35:0]   _zz_9024;
  wire       [17:0]   _zz_9025;
  wire       [35:0]   _zz_9026;
  wire       [35:0]   _zz_9027;
  wire       [35:0]   _zz_9028;
  wire       [35:0]   _zz_9029;
  wire       [35:0]   _zz_9030;
  wire       [26:0]   _zz_9031;
  wire       [35:0]   _zz_9032;
  wire       [17:0]   _zz_9033;
  wire       [35:0]   _zz_9034;
  wire       [35:0]   _zz_9035;
  wire       [35:0]   _zz_9036;
  wire       [35:0]   _zz_9037;
  wire       [35:0]   _zz_9038;
  wire       [26:0]   _zz_9039;
  wire       [35:0]   _zz_9040;
  wire       [17:0]   _zz_9041;
  wire       [17:0]   _zz_9042;
  wire       [35:0]   _zz_9043;
  wire       [35:0]   _zz_9044;
  wire       [17:0]   _zz_9045;
  wire       [35:0]   _zz_9046;
  wire       [35:0]   _zz_9047;
  wire       [35:0]   _zz_9048;
  wire       [17:0]   _zz_9049;
  wire       [35:0]   _zz_9050;
  wire       [35:0]   _zz_9051;
  wire       [35:0]   _zz_9052;
  wire       [35:0]   _zz_9053;
  wire       [35:0]   _zz_9054;
  wire       [35:0]   _zz_9055;
  wire       [26:0]   _zz_9056;
  wire       [35:0]   _zz_9057;
  wire       [17:0]   _zz_9058;
  wire       [35:0]   _zz_9059;
  wire       [35:0]   _zz_9060;
  wire       [35:0]   _zz_9061;
  wire       [35:0]   _zz_9062;
  wire       [35:0]   _zz_9063;
  wire       [26:0]   _zz_9064;
  wire       [35:0]   _zz_9065;
  wire       [17:0]   _zz_9066;
  wire       [35:0]   _zz_9067;
  wire       [35:0]   _zz_9068;
  wire       [35:0]   _zz_9069;
  wire       [35:0]   _zz_9070;
  wire       [35:0]   _zz_9071;
  wire       [26:0]   _zz_9072;
  wire       [35:0]   _zz_9073;
  wire       [17:0]   _zz_9074;
  wire       [35:0]   _zz_9075;
  wire       [35:0]   _zz_9076;
  wire       [35:0]   _zz_9077;
  wire       [35:0]   _zz_9078;
  wire       [35:0]   _zz_9079;
  wire       [26:0]   _zz_9080;
  wire       [35:0]   _zz_9081;
  wire       [17:0]   _zz_9082;
  wire       [17:0]   _zz_9083;
  wire       [35:0]   _zz_9084;
  wire       [35:0]   _zz_9085;
  wire       [17:0]   _zz_9086;
  wire       [35:0]   _zz_9087;
  wire       [35:0]   _zz_9088;
  wire       [35:0]   _zz_9089;
  wire       [17:0]   _zz_9090;
  wire       [35:0]   _zz_9091;
  wire       [35:0]   _zz_9092;
  wire       [35:0]   _zz_9093;
  wire       [35:0]   _zz_9094;
  wire       [35:0]   _zz_9095;
  wire       [35:0]   _zz_9096;
  wire       [26:0]   _zz_9097;
  wire       [35:0]   _zz_9098;
  wire       [17:0]   _zz_9099;
  wire       [35:0]   _zz_9100;
  wire       [35:0]   _zz_9101;
  wire       [35:0]   _zz_9102;
  wire       [35:0]   _zz_9103;
  wire       [35:0]   _zz_9104;
  wire       [26:0]   _zz_9105;
  wire       [35:0]   _zz_9106;
  wire       [17:0]   _zz_9107;
  wire       [35:0]   _zz_9108;
  wire       [35:0]   _zz_9109;
  wire       [35:0]   _zz_9110;
  wire       [35:0]   _zz_9111;
  wire       [35:0]   _zz_9112;
  wire       [26:0]   _zz_9113;
  wire       [35:0]   _zz_9114;
  wire       [17:0]   _zz_9115;
  wire       [35:0]   _zz_9116;
  wire       [35:0]   _zz_9117;
  wire       [35:0]   _zz_9118;
  wire       [35:0]   _zz_9119;
  wire       [35:0]   _zz_9120;
  wire       [26:0]   _zz_9121;
  wire       [35:0]   _zz_9122;
  wire       [17:0]   _zz_9123;
  wire       [17:0]   _zz_9124;
  wire       [35:0]   _zz_9125;
  wire       [35:0]   _zz_9126;
  wire       [17:0]   _zz_9127;
  wire       [35:0]   _zz_9128;
  wire       [35:0]   _zz_9129;
  wire       [35:0]   _zz_9130;
  wire       [17:0]   _zz_9131;
  wire       [35:0]   _zz_9132;
  wire       [35:0]   _zz_9133;
  wire       [35:0]   _zz_9134;
  wire       [35:0]   _zz_9135;
  wire       [35:0]   _zz_9136;
  wire       [35:0]   _zz_9137;
  wire       [26:0]   _zz_9138;
  wire       [35:0]   _zz_9139;
  wire       [17:0]   _zz_9140;
  wire       [35:0]   _zz_9141;
  wire       [35:0]   _zz_9142;
  wire       [35:0]   _zz_9143;
  wire       [35:0]   _zz_9144;
  wire       [35:0]   _zz_9145;
  wire       [26:0]   _zz_9146;
  wire       [35:0]   _zz_9147;
  wire       [17:0]   _zz_9148;
  wire       [35:0]   _zz_9149;
  wire       [35:0]   _zz_9150;
  wire       [35:0]   _zz_9151;
  wire       [35:0]   _zz_9152;
  wire       [35:0]   _zz_9153;
  wire       [26:0]   _zz_9154;
  wire       [35:0]   _zz_9155;
  wire       [17:0]   _zz_9156;
  wire       [35:0]   _zz_9157;
  wire       [35:0]   _zz_9158;
  wire       [35:0]   _zz_9159;
  wire       [35:0]   _zz_9160;
  wire       [35:0]   _zz_9161;
  wire       [26:0]   _zz_9162;
  wire       [35:0]   _zz_9163;
  wire       [17:0]   _zz_9164;
  wire       [17:0]   _zz_9165;
  wire       [35:0]   _zz_9166;
  wire       [35:0]   _zz_9167;
  wire       [17:0]   _zz_9168;
  wire       [35:0]   _zz_9169;
  wire       [35:0]   _zz_9170;
  wire       [35:0]   _zz_9171;
  wire       [17:0]   _zz_9172;
  wire       [35:0]   _zz_9173;
  wire       [35:0]   _zz_9174;
  wire       [35:0]   _zz_9175;
  wire       [35:0]   _zz_9176;
  wire       [35:0]   _zz_9177;
  wire       [35:0]   _zz_9178;
  wire       [26:0]   _zz_9179;
  wire       [35:0]   _zz_9180;
  wire       [17:0]   _zz_9181;
  wire       [35:0]   _zz_9182;
  wire       [35:0]   _zz_9183;
  wire       [35:0]   _zz_9184;
  wire       [35:0]   _zz_9185;
  wire       [35:0]   _zz_9186;
  wire       [26:0]   _zz_9187;
  wire       [35:0]   _zz_9188;
  wire       [17:0]   _zz_9189;
  wire       [35:0]   _zz_9190;
  wire       [35:0]   _zz_9191;
  wire       [35:0]   _zz_9192;
  wire       [35:0]   _zz_9193;
  wire       [35:0]   _zz_9194;
  wire       [26:0]   _zz_9195;
  wire       [35:0]   _zz_9196;
  wire       [17:0]   _zz_9197;
  wire       [35:0]   _zz_9198;
  wire       [35:0]   _zz_9199;
  wire       [35:0]   _zz_9200;
  wire       [35:0]   _zz_9201;
  wire       [35:0]   _zz_9202;
  wire       [26:0]   _zz_9203;
  wire       [35:0]   _zz_9204;
  wire       [17:0]   _zz_9205;
  wire       [17:0]   _zz_9206;
  wire       [35:0]   _zz_9207;
  wire       [35:0]   _zz_9208;
  wire       [17:0]   _zz_9209;
  wire       [35:0]   _zz_9210;
  wire       [35:0]   _zz_9211;
  wire       [35:0]   _zz_9212;
  wire       [17:0]   _zz_9213;
  wire       [35:0]   _zz_9214;
  wire       [35:0]   _zz_9215;
  wire       [35:0]   _zz_9216;
  wire       [35:0]   _zz_9217;
  wire       [35:0]   _zz_9218;
  wire       [35:0]   _zz_9219;
  wire       [26:0]   _zz_9220;
  wire       [35:0]   _zz_9221;
  wire       [17:0]   _zz_9222;
  wire       [35:0]   _zz_9223;
  wire       [35:0]   _zz_9224;
  wire       [35:0]   _zz_9225;
  wire       [35:0]   _zz_9226;
  wire       [35:0]   _zz_9227;
  wire       [26:0]   _zz_9228;
  wire       [35:0]   _zz_9229;
  wire       [17:0]   _zz_9230;
  wire       [35:0]   _zz_9231;
  wire       [35:0]   _zz_9232;
  wire       [35:0]   _zz_9233;
  wire       [35:0]   _zz_9234;
  wire       [35:0]   _zz_9235;
  wire       [26:0]   _zz_9236;
  wire       [35:0]   _zz_9237;
  wire       [17:0]   _zz_9238;
  wire       [35:0]   _zz_9239;
  wire       [35:0]   _zz_9240;
  wire       [35:0]   _zz_9241;
  wire       [35:0]   _zz_9242;
  wire       [35:0]   _zz_9243;
  wire       [26:0]   _zz_9244;
  wire       [35:0]   _zz_9245;
  wire       [17:0]   _zz_9246;
  wire       [17:0]   _zz_9247;
  wire       [35:0]   _zz_9248;
  wire       [35:0]   _zz_9249;
  wire       [17:0]   _zz_9250;
  wire       [35:0]   _zz_9251;
  wire       [35:0]   _zz_9252;
  wire       [35:0]   _zz_9253;
  wire       [17:0]   _zz_9254;
  wire       [35:0]   _zz_9255;
  wire       [35:0]   _zz_9256;
  wire       [35:0]   _zz_9257;
  wire       [35:0]   _zz_9258;
  wire       [35:0]   _zz_9259;
  wire       [35:0]   _zz_9260;
  wire       [26:0]   _zz_9261;
  wire       [35:0]   _zz_9262;
  wire       [17:0]   _zz_9263;
  wire       [35:0]   _zz_9264;
  wire       [35:0]   _zz_9265;
  wire       [35:0]   _zz_9266;
  wire       [35:0]   _zz_9267;
  wire       [35:0]   _zz_9268;
  wire       [26:0]   _zz_9269;
  wire       [35:0]   _zz_9270;
  wire       [17:0]   _zz_9271;
  wire       [35:0]   _zz_9272;
  wire       [35:0]   _zz_9273;
  wire       [35:0]   _zz_9274;
  wire       [35:0]   _zz_9275;
  wire       [35:0]   _zz_9276;
  wire       [26:0]   _zz_9277;
  wire       [35:0]   _zz_9278;
  wire       [17:0]   _zz_9279;
  wire       [35:0]   _zz_9280;
  wire       [35:0]   _zz_9281;
  wire       [35:0]   _zz_9282;
  wire       [35:0]   _zz_9283;
  wire       [35:0]   _zz_9284;
  wire       [26:0]   _zz_9285;
  wire       [35:0]   _zz_9286;
  wire       [17:0]   _zz_9287;
  wire       [17:0]   _zz_9288;
  wire       [35:0]   _zz_9289;
  wire       [35:0]   _zz_9290;
  wire       [17:0]   _zz_9291;
  wire       [35:0]   _zz_9292;
  wire       [35:0]   _zz_9293;
  wire       [35:0]   _zz_9294;
  wire       [17:0]   _zz_9295;
  wire       [35:0]   _zz_9296;
  wire       [35:0]   _zz_9297;
  wire       [35:0]   _zz_9298;
  wire       [35:0]   _zz_9299;
  wire       [35:0]   _zz_9300;
  wire       [35:0]   _zz_9301;
  wire       [26:0]   _zz_9302;
  wire       [35:0]   _zz_9303;
  wire       [17:0]   _zz_9304;
  wire       [35:0]   _zz_9305;
  wire       [35:0]   _zz_9306;
  wire       [35:0]   _zz_9307;
  wire       [35:0]   _zz_9308;
  wire       [35:0]   _zz_9309;
  wire       [26:0]   _zz_9310;
  wire       [35:0]   _zz_9311;
  wire       [17:0]   _zz_9312;
  wire       [35:0]   _zz_9313;
  wire       [35:0]   _zz_9314;
  wire       [35:0]   _zz_9315;
  wire       [35:0]   _zz_9316;
  wire       [35:0]   _zz_9317;
  wire       [26:0]   _zz_9318;
  wire       [35:0]   _zz_9319;
  wire       [17:0]   _zz_9320;
  wire       [35:0]   _zz_9321;
  wire       [35:0]   _zz_9322;
  wire       [35:0]   _zz_9323;
  wire       [35:0]   _zz_9324;
  wire       [35:0]   _zz_9325;
  wire       [26:0]   _zz_9326;
  wire       [35:0]   _zz_9327;
  wire       [17:0]   _zz_9328;
  wire       [17:0]   _zz_9329;
  wire       [35:0]   _zz_9330;
  wire       [35:0]   _zz_9331;
  wire       [17:0]   _zz_9332;
  wire       [35:0]   _zz_9333;
  wire       [35:0]   _zz_9334;
  wire       [35:0]   _zz_9335;
  wire       [17:0]   _zz_9336;
  wire       [35:0]   _zz_9337;
  wire       [35:0]   _zz_9338;
  wire       [35:0]   _zz_9339;
  wire       [35:0]   _zz_9340;
  wire       [35:0]   _zz_9341;
  wire       [35:0]   _zz_9342;
  wire       [26:0]   _zz_9343;
  wire       [35:0]   _zz_9344;
  wire       [17:0]   _zz_9345;
  wire       [35:0]   _zz_9346;
  wire       [35:0]   _zz_9347;
  wire       [35:0]   _zz_9348;
  wire       [35:0]   _zz_9349;
  wire       [35:0]   _zz_9350;
  wire       [26:0]   _zz_9351;
  wire       [35:0]   _zz_9352;
  wire       [17:0]   _zz_9353;
  wire       [35:0]   _zz_9354;
  wire       [35:0]   _zz_9355;
  wire       [35:0]   _zz_9356;
  wire       [35:0]   _zz_9357;
  wire       [35:0]   _zz_9358;
  wire       [26:0]   _zz_9359;
  wire       [35:0]   _zz_9360;
  wire       [17:0]   _zz_9361;
  wire       [35:0]   _zz_9362;
  wire       [35:0]   _zz_9363;
  wire       [35:0]   _zz_9364;
  wire       [35:0]   _zz_9365;
  wire       [35:0]   _zz_9366;
  wire       [26:0]   _zz_9367;
  wire       [35:0]   _zz_9368;
  wire       [17:0]   _zz_9369;
  wire       [17:0]   _zz_9370;
  wire       [35:0]   _zz_9371;
  wire       [35:0]   _zz_9372;
  wire       [17:0]   _zz_9373;
  wire       [35:0]   _zz_9374;
  wire       [35:0]   _zz_9375;
  wire       [35:0]   _zz_9376;
  wire       [17:0]   _zz_9377;
  wire       [35:0]   _zz_9378;
  wire       [35:0]   _zz_9379;
  wire       [35:0]   _zz_9380;
  wire       [35:0]   _zz_9381;
  wire       [35:0]   _zz_9382;
  wire       [35:0]   _zz_9383;
  wire       [26:0]   _zz_9384;
  wire       [35:0]   _zz_9385;
  wire       [17:0]   _zz_9386;
  wire       [35:0]   _zz_9387;
  wire       [35:0]   _zz_9388;
  wire       [35:0]   _zz_9389;
  wire       [35:0]   _zz_9390;
  wire       [35:0]   _zz_9391;
  wire       [26:0]   _zz_9392;
  wire       [35:0]   _zz_9393;
  wire       [17:0]   _zz_9394;
  wire       [35:0]   _zz_9395;
  wire       [35:0]   _zz_9396;
  wire       [35:0]   _zz_9397;
  wire       [35:0]   _zz_9398;
  wire       [35:0]   _zz_9399;
  wire       [26:0]   _zz_9400;
  wire       [35:0]   _zz_9401;
  wire       [17:0]   _zz_9402;
  wire       [35:0]   _zz_9403;
  wire       [35:0]   _zz_9404;
  wire       [35:0]   _zz_9405;
  wire       [35:0]   _zz_9406;
  wire       [35:0]   _zz_9407;
  wire       [26:0]   _zz_9408;
  wire       [35:0]   _zz_9409;
  wire       [17:0]   _zz_9410;
  wire       [17:0]   _zz_9411;
  wire       [35:0]   _zz_9412;
  wire       [35:0]   _zz_9413;
  wire       [17:0]   _zz_9414;
  wire       [35:0]   _zz_9415;
  wire       [35:0]   _zz_9416;
  wire       [35:0]   _zz_9417;
  wire       [17:0]   _zz_9418;
  wire       [35:0]   _zz_9419;
  wire       [35:0]   _zz_9420;
  wire       [35:0]   _zz_9421;
  wire       [35:0]   _zz_9422;
  wire       [35:0]   _zz_9423;
  wire       [35:0]   _zz_9424;
  wire       [26:0]   _zz_9425;
  wire       [35:0]   _zz_9426;
  wire       [17:0]   _zz_9427;
  wire       [35:0]   _zz_9428;
  wire       [35:0]   _zz_9429;
  wire       [35:0]   _zz_9430;
  wire       [35:0]   _zz_9431;
  wire       [35:0]   _zz_9432;
  wire       [26:0]   _zz_9433;
  wire       [35:0]   _zz_9434;
  wire       [17:0]   _zz_9435;
  wire       [35:0]   _zz_9436;
  wire       [35:0]   _zz_9437;
  wire       [35:0]   _zz_9438;
  wire       [35:0]   _zz_9439;
  wire       [35:0]   _zz_9440;
  wire       [26:0]   _zz_9441;
  wire       [35:0]   _zz_9442;
  wire       [17:0]   _zz_9443;
  wire       [35:0]   _zz_9444;
  wire       [35:0]   _zz_9445;
  wire       [35:0]   _zz_9446;
  wire       [35:0]   _zz_9447;
  wire       [35:0]   _zz_9448;
  wire       [26:0]   _zz_9449;
  wire       [35:0]   _zz_9450;
  wire       [17:0]   _zz_9451;
  wire       [17:0]   _zz_9452;
  wire       [35:0]   _zz_9453;
  wire       [35:0]   _zz_9454;
  wire       [17:0]   _zz_9455;
  wire       [35:0]   _zz_9456;
  wire       [35:0]   _zz_9457;
  wire       [35:0]   _zz_9458;
  wire       [17:0]   _zz_9459;
  wire       [35:0]   _zz_9460;
  wire       [35:0]   _zz_9461;
  wire       [35:0]   _zz_9462;
  wire       [35:0]   _zz_9463;
  wire       [35:0]   _zz_9464;
  wire       [35:0]   _zz_9465;
  wire       [26:0]   _zz_9466;
  wire       [35:0]   _zz_9467;
  wire       [17:0]   _zz_9468;
  wire       [35:0]   _zz_9469;
  wire       [35:0]   _zz_9470;
  wire       [35:0]   _zz_9471;
  wire       [35:0]   _zz_9472;
  wire       [35:0]   _zz_9473;
  wire       [26:0]   _zz_9474;
  wire       [35:0]   _zz_9475;
  wire       [17:0]   _zz_9476;
  wire       [35:0]   _zz_9477;
  wire       [35:0]   _zz_9478;
  wire       [35:0]   _zz_9479;
  wire       [35:0]   _zz_9480;
  wire       [35:0]   _zz_9481;
  wire       [26:0]   _zz_9482;
  wire       [35:0]   _zz_9483;
  wire       [17:0]   _zz_9484;
  wire       [35:0]   _zz_9485;
  wire       [35:0]   _zz_9486;
  wire       [35:0]   _zz_9487;
  wire       [35:0]   _zz_9488;
  wire       [35:0]   _zz_9489;
  wire       [26:0]   _zz_9490;
  wire       [35:0]   _zz_9491;
  wire       [17:0]   _zz_9492;
  wire       [17:0]   _zz_9493;
  wire       [35:0]   _zz_9494;
  wire       [35:0]   _zz_9495;
  wire       [17:0]   _zz_9496;
  wire       [35:0]   _zz_9497;
  wire       [35:0]   _zz_9498;
  wire       [35:0]   _zz_9499;
  wire       [17:0]   _zz_9500;
  wire       [35:0]   _zz_9501;
  wire       [35:0]   _zz_9502;
  wire       [35:0]   _zz_9503;
  wire       [35:0]   _zz_9504;
  wire       [35:0]   _zz_9505;
  wire       [35:0]   _zz_9506;
  wire       [26:0]   _zz_9507;
  wire       [35:0]   _zz_9508;
  wire       [17:0]   _zz_9509;
  wire       [35:0]   _zz_9510;
  wire       [35:0]   _zz_9511;
  wire       [35:0]   _zz_9512;
  wire       [35:0]   _zz_9513;
  wire       [35:0]   _zz_9514;
  wire       [26:0]   _zz_9515;
  wire       [35:0]   _zz_9516;
  wire       [17:0]   _zz_9517;
  wire       [35:0]   _zz_9518;
  wire       [35:0]   _zz_9519;
  wire       [35:0]   _zz_9520;
  wire       [35:0]   _zz_9521;
  wire       [35:0]   _zz_9522;
  wire       [26:0]   _zz_9523;
  wire       [35:0]   _zz_9524;
  wire       [17:0]   _zz_9525;
  wire       [35:0]   _zz_9526;
  wire       [35:0]   _zz_9527;
  wire       [35:0]   _zz_9528;
  wire       [35:0]   _zz_9529;
  wire       [35:0]   _zz_9530;
  wire       [26:0]   _zz_9531;
  wire       [35:0]   _zz_9532;
  wire       [17:0]   _zz_9533;
  wire       [17:0]   _zz_9534;
  wire       [35:0]   _zz_9535;
  wire       [35:0]   _zz_9536;
  wire       [17:0]   _zz_9537;
  wire       [35:0]   _zz_9538;
  wire       [35:0]   _zz_9539;
  wire       [35:0]   _zz_9540;
  wire       [17:0]   _zz_9541;
  wire       [35:0]   _zz_9542;
  wire       [35:0]   _zz_9543;
  wire       [35:0]   _zz_9544;
  wire       [35:0]   _zz_9545;
  wire       [35:0]   _zz_9546;
  wire       [35:0]   _zz_9547;
  wire       [26:0]   _zz_9548;
  wire       [35:0]   _zz_9549;
  wire       [17:0]   _zz_9550;
  wire       [35:0]   _zz_9551;
  wire       [35:0]   _zz_9552;
  wire       [35:0]   _zz_9553;
  wire       [35:0]   _zz_9554;
  wire       [35:0]   _zz_9555;
  wire       [26:0]   _zz_9556;
  wire       [35:0]   _zz_9557;
  wire       [17:0]   _zz_9558;
  wire       [35:0]   _zz_9559;
  wire       [35:0]   _zz_9560;
  wire       [35:0]   _zz_9561;
  wire       [35:0]   _zz_9562;
  wire       [35:0]   _zz_9563;
  wire       [26:0]   _zz_9564;
  wire       [35:0]   _zz_9565;
  wire       [17:0]   _zz_9566;
  wire       [35:0]   _zz_9567;
  wire       [35:0]   _zz_9568;
  wire       [35:0]   _zz_9569;
  wire       [35:0]   _zz_9570;
  wire       [35:0]   _zz_9571;
  wire       [26:0]   _zz_9572;
  wire       [35:0]   _zz_9573;
  wire       [17:0]   _zz_9574;
  wire       [17:0]   _zz_9575;
  wire       [35:0]   _zz_9576;
  wire       [35:0]   _zz_9577;
  wire       [17:0]   _zz_9578;
  wire       [35:0]   _zz_9579;
  wire       [35:0]   _zz_9580;
  wire       [35:0]   _zz_9581;
  wire       [17:0]   _zz_9582;
  wire       [35:0]   _zz_9583;
  wire       [35:0]   _zz_9584;
  wire       [35:0]   _zz_9585;
  wire       [35:0]   _zz_9586;
  wire       [35:0]   _zz_9587;
  wire       [35:0]   _zz_9588;
  wire       [26:0]   _zz_9589;
  wire       [35:0]   _zz_9590;
  wire       [17:0]   _zz_9591;
  wire       [35:0]   _zz_9592;
  wire       [35:0]   _zz_9593;
  wire       [35:0]   _zz_9594;
  wire       [35:0]   _zz_9595;
  wire       [35:0]   _zz_9596;
  wire       [26:0]   _zz_9597;
  wire       [35:0]   _zz_9598;
  wire       [17:0]   _zz_9599;
  wire       [35:0]   _zz_9600;
  wire       [35:0]   _zz_9601;
  wire       [35:0]   _zz_9602;
  wire       [35:0]   _zz_9603;
  wire       [35:0]   _zz_9604;
  wire       [26:0]   _zz_9605;
  wire       [35:0]   _zz_9606;
  wire       [17:0]   _zz_9607;
  wire       [35:0]   _zz_9608;
  wire       [35:0]   _zz_9609;
  wire       [35:0]   _zz_9610;
  wire       [35:0]   _zz_9611;
  wire       [35:0]   _zz_9612;
  wire       [26:0]   _zz_9613;
  wire       [35:0]   _zz_9614;
  wire       [17:0]   _zz_9615;
  wire       [17:0]   _zz_9616;
  wire       [35:0]   _zz_9617;
  wire       [35:0]   _zz_9618;
  wire       [17:0]   _zz_9619;
  wire       [35:0]   _zz_9620;
  wire       [35:0]   _zz_9621;
  wire       [35:0]   _zz_9622;
  wire       [17:0]   _zz_9623;
  wire       [35:0]   _zz_9624;
  wire       [35:0]   _zz_9625;
  wire       [35:0]   _zz_9626;
  wire       [35:0]   _zz_9627;
  wire       [35:0]   _zz_9628;
  wire       [35:0]   _zz_9629;
  wire       [26:0]   _zz_9630;
  wire       [35:0]   _zz_9631;
  wire       [17:0]   _zz_9632;
  wire       [35:0]   _zz_9633;
  wire       [35:0]   _zz_9634;
  wire       [35:0]   _zz_9635;
  wire       [35:0]   _zz_9636;
  wire       [35:0]   _zz_9637;
  wire       [26:0]   _zz_9638;
  wire       [35:0]   _zz_9639;
  wire       [17:0]   _zz_9640;
  wire       [35:0]   _zz_9641;
  wire       [35:0]   _zz_9642;
  wire       [35:0]   _zz_9643;
  wire       [35:0]   _zz_9644;
  wire       [35:0]   _zz_9645;
  wire       [26:0]   _zz_9646;
  wire       [35:0]   _zz_9647;
  wire       [17:0]   _zz_9648;
  wire       [35:0]   _zz_9649;
  wire       [35:0]   _zz_9650;
  wire       [35:0]   _zz_9651;
  wire       [35:0]   _zz_9652;
  wire       [35:0]   _zz_9653;
  wire       [26:0]   _zz_9654;
  wire       [35:0]   _zz_9655;
  wire       [17:0]   _zz_9656;
  wire       [17:0]   _zz_9657;
  wire       [35:0]   _zz_9658;
  wire       [35:0]   _zz_9659;
  wire       [17:0]   _zz_9660;
  wire       [35:0]   _zz_9661;
  wire       [35:0]   _zz_9662;
  wire       [35:0]   _zz_9663;
  wire       [17:0]   _zz_9664;
  wire       [35:0]   _zz_9665;
  wire       [35:0]   _zz_9666;
  wire       [35:0]   _zz_9667;
  wire       [35:0]   _zz_9668;
  wire       [35:0]   _zz_9669;
  wire       [35:0]   _zz_9670;
  wire       [26:0]   _zz_9671;
  wire       [35:0]   _zz_9672;
  wire       [17:0]   _zz_9673;
  wire       [35:0]   _zz_9674;
  wire       [35:0]   _zz_9675;
  wire       [35:0]   _zz_9676;
  wire       [35:0]   _zz_9677;
  wire       [35:0]   _zz_9678;
  wire       [26:0]   _zz_9679;
  wire       [35:0]   _zz_9680;
  wire       [17:0]   _zz_9681;
  wire       [35:0]   _zz_9682;
  wire       [35:0]   _zz_9683;
  wire       [35:0]   _zz_9684;
  wire       [35:0]   _zz_9685;
  wire       [35:0]   _zz_9686;
  wire       [26:0]   _zz_9687;
  wire       [35:0]   _zz_9688;
  wire       [17:0]   _zz_9689;
  wire       [35:0]   _zz_9690;
  wire       [35:0]   _zz_9691;
  wire       [35:0]   _zz_9692;
  wire       [35:0]   _zz_9693;
  wire       [35:0]   _zz_9694;
  wire       [26:0]   _zz_9695;
  wire       [35:0]   _zz_9696;
  wire       [17:0]   _zz_9697;
  wire       [17:0]   _zz_9698;
  wire       [35:0]   _zz_9699;
  wire       [35:0]   _zz_9700;
  wire       [17:0]   _zz_9701;
  wire       [35:0]   _zz_9702;
  wire       [35:0]   _zz_9703;
  wire       [35:0]   _zz_9704;
  wire       [17:0]   _zz_9705;
  wire       [35:0]   _zz_9706;
  wire       [35:0]   _zz_9707;
  wire       [35:0]   _zz_9708;
  wire       [35:0]   _zz_9709;
  wire       [35:0]   _zz_9710;
  wire       [35:0]   _zz_9711;
  wire       [26:0]   _zz_9712;
  wire       [35:0]   _zz_9713;
  wire       [17:0]   _zz_9714;
  wire       [35:0]   _zz_9715;
  wire       [35:0]   _zz_9716;
  wire       [35:0]   _zz_9717;
  wire       [35:0]   _zz_9718;
  wire       [35:0]   _zz_9719;
  wire       [26:0]   _zz_9720;
  wire       [35:0]   _zz_9721;
  wire       [17:0]   _zz_9722;
  wire       [35:0]   _zz_9723;
  wire       [35:0]   _zz_9724;
  wire       [35:0]   _zz_9725;
  wire       [35:0]   _zz_9726;
  wire       [35:0]   _zz_9727;
  wire       [26:0]   _zz_9728;
  wire       [35:0]   _zz_9729;
  wire       [17:0]   _zz_9730;
  wire       [35:0]   _zz_9731;
  wire       [35:0]   _zz_9732;
  wire       [35:0]   _zz_9733;
  wire       [35:0]   _zz_9734;
  wire       [35:0]   _zz_9735;
  wire       [26:0]   _zz_9736;
  wire       [35:0]   _zz_9737;
  wire       [17:0]   _zz_9738;
  wire       [17:0]   _zz_9739;
  wire       [35:0]   _zz_9740;
  wire       [35:0]   _zz_9741;
  wire       [17:0]   _zz_9742;
  wire       [35:0]   _zz_9743;
  wire       [35:0]   _zz_9744;
  wire       [35:0]   _zz_9745;
  wire       [17:0]   _zz_9746;
  wire       [35:0]   _zz_9747;
  wire       [35:0]   _zz_9748;
  wire       [35:0]   _zz_9749;
  wire       [35:0]   _zz_9750;
  wire       [35:0]   _zz_9751;
  wire       [35:0]   _zz_9752;
  wire       [26:0]   _zz_9753;
  wire       [35:0]   _zz_9754;
  wire       [17:0]   _zz_9755;
  wire       [35:0]   _zz_9756;
  wire       [35:0]   _zz_9757;
  wire       [35:0]   _zz_9758;
  wire       [35:0]   _zz_9759;
  wire       [35:0]   _zz_9760;
  wire       [26:0]   _zz_9761;
  wire       [35:0]   _zz_9762;
  wire       [17:0]   _zz_9763;
  wire       [35:0]   _zz_9764;
  wire       [35:0]   _zz_9765;
  wire       [35:0]   _zz_9766;
  wire       [35:0]   _zz_9767;
  wire       [35:0]   _zz_9768;
  wire       [26:0]   _zz_9769;
  wire       [35:0]   _zz_9770;
  wire       [17:0]   _zz_9771;
  wire       [35:0]   _zz_9772;
  wire       [35:0]   _zz_9773;
  wire       [35:0]   _zz_9774;
  wire       [35:0]   _zz_9775;
  wire       [35:0]   _zz_9776;
  wire       [26:0]   _zz_9777;
  wire       [35:0]   _zz_9778;
  wire       [17:0]   _zz_9779;
  wire       [17:0]   _zz_9780;
  wire       [35:0]   _zz_9781;
  wire       [35:0]   _zz_9782;
  wire       [17:0]   _zz_9783;
  wire       [35:0]   _zz_9784;
  wire       [35:0]   _zz_9785;
  wire       [35:0]   _zz_9786;
  wire       [17:0]   _zz_9787;
  wire       [35:0]   _zz_9788;
  wire       [35:0]   _zz_9789;
  wire       [35:0]   _zz_9790;
  wire       [35:0]   _zz_9791;
  wire       [35:0]   _zz_9792;
  wire       [35:0]   _zz_9793;
  wire       [26:0]   _zz_9794;
  wire       [35:0]   _zz_9795;
  wire       [17:0]   _zz_9796;
  wire       [35:0]   _zz_9797;
  wire       [35:0]   _zz_9798;
  wire       [35:0]   _zz_9799;
  wire       [35:0]   _zz_9800;
  wire       [35:0]   _zz_9801;
  wire       [26:0]   _zz_9802;
  wire       [35:0]   _zz_9803;
  wire       [17:0]   _zz_9804;
  wire       [35:0]   _zz_9805;
  wire       [35:0]   _zz_9806;
  wire       [35:0]   _zz_9807;
  wire       [35:0]   _zz_9808;
  wire       [35:0]   _zz_9809;
  wire       [26:0]   _zz_9810;
  wire       [35:0]   _zz_9811;
  wire       [17:0]   _zz_9812;
  wire       [35:0]   _zz_9813;
  wire       [35:0]   _zz_9814;
  wire       [35:0]   _zz_9815;
  wire       [35:0]   _zz_9816;
  wire       [35:0]   _zz_9817;
  wire       [26:0]   _zz_9818;
  wire       [35:0]   _zz_9819;
  wire       [17:0]   _zz_9820;
  wire       [17:0]   _zz_9821;
  wire       [35:0]   _zz_9822;
  wire       [35:0]   _zz_9823;
  wire       [17:0]   _zz_9824;
  wire       [35:0]   _zz_9825;
  wire       [35:0]   _zz_9826;
  wire       [35:0]   _zz_9827;
  wire       [17:0]   _zz_9828;
  wire       [35:0]   _zz_9829;
  wire       [35:0]   _zz_9830;
  wire       [35:0]   _zz_9831;
  wire       [35:0]   _zz_9832;
  wire       [35:0]   _zz_9833;
  wire       [35:0]   _zz_9834;
  wire       [26:0]   _zz_9835;
  wire       [35:0]   _zz_9836;
  wire       [17:0]   _zz_9837;
  wire       [35:0]   _zz_9838;
  wire       [35:0]   _zz_9839;
  wire       [35:0]   _zz_9840;
  wire       [35:0]   _zz_9841;
  wire       [35:0]   _zz_9842;
  wire       [26:0]   _zz_9843;
  wire       [35:0]   _zz_9844;
  wire       [17:0]   _zz_9845;
  wire       [35:0]   _zz_9846;
  wire       [35:0]   _zz_9847;
  wire       [35:0]   _zz_9848;
  wire       [35:0]   _zz_9849;
  wire       [35:0]   _zz_9850;
  wire       [26:0]   _zz_9851;
  wire       [35:0]   _zz_9852;
  wire       [17:0]   _zz_9853;
  wire       [35:0]   _zz_9854;
  wire       [35:0]   _zz_9855;
  wire       [35:0]   _zz_9856;
  wire       [35:0]   _zz_9857;
  wire       [35:0]   _zz_9858;
  wire       [26:0]   _zz_9859;
  wire       [35:0]   _zz_9860;
  wire       [17:0]   _zz_9861;
  wire       [17:0]   _zz_9862;
  wire       [35:0]   _zz_9863;
  wire       [35:0]   _zz_9864;
  wire       [17:0]   _zz_9865;
  wire       [35:0]   _zz_9866;
  wire       [35:0]   _zz_9867;
  wire       [35:0]   _zz_9868;
  wire       [17:0]   _zz_9869;
  wire       [35:0]   _zz_9870;
  wire       [35:0]   _zz_9871;
  wire       [35:0]   _zz_9872;
  wire       [35:0]   _zz_9873;
  wire       [35:0]   _zz_9874;
  wire       [35:0]   _zz_9875;
  wire       [26:0]   _zz_9876;
  wire       [35:0]   _zz_9877;
  wire       [17:0]   _zz_9878;
  wire       [35:0]   _zz_9879;
  wire       [35:0]   _zz_9880;
  wire       [35:0]   _zz_9881;
  wire       [35:0]   _zz_9882;
  wire       [35:0]   _zz_9883;
  wire       [26:0]   _zz_9884;
  wire       [35:0]   _zz_9885;
  wire       [17:0]   _zz_9886;
  wire       [35:0]   _zz_9887;
  wire       [35:0]   _zz_9888;
  wire       [35:0]   _zz_9889;
  wire       [35:0]   _zz_9890;
  wire       [35:0]   _zz_9891;
  wire       [26:0]   _zz_9892;
  wire       [35:0]   _zz_9893;
  wire       [17:0]   _zz_9894;
  wire       [35:0]   _zz_9895;
  wire       [35:0]   _zz_9896;
  wire       [35:0]   _zz_9897;
  wire       [35:0]   _zz_9898;
  wire       [35:0]   _zz_9899;
  wire       [26:0]   _zz_9900;
  wire       [35:0]   _zz_9901;
  wire       [17:0]   _zz_9902;
  wire       [17:0]   _zz_9903;
  wire       [35:0]   _zz_9904;
  wire       [35:0]   _zz_9905;
  wire       [17:0]   _zz_9906;
  wire       [35:0]   _zz_9907;
  wire       [35:0]   _zz_9908;
  wire       [35:0]   _zz_9909;
  wire       [17:0]   _zz_9910;
  wire       [35:0]   _zz_9911;
  wire       [35:0]   _zz_9912;
  wire       [35:0]   _zz_9913;
  wire       [35:0]   _zz_9914;
  wire       [35:0]   _zz_9915;
  wire       [35:0]   _zz_9916;
  wire       [26:0]   _zz_9917;
  wire       [35:0]   _zz_9918;
  wire       [17:0]   _zz_9919;
  wire       [35:0]   _zz_9920;
  wire       [35:0]   _zz_9921;
  wire       [35:0]   _zz_9922;
  wire       [35:0]   _zz_9923;
  wire       [35:0]   _zz_9924;
  wire       [26:0]   _zz_9925;
  wire       [35:0]   _zz_9926;
  wire       [17:0]   _zz_9927;
  wire       [35:0]   _zz_9928;
  wire       [35:0]   _zz_9929;
  wire       [35:0]   _zz_9930;
  wire       [35:0]   _zz_9931;
  wire       [35:0]   _zz_9932;
  wire       [26:0]   _zz_9933;
  wire       [35:0]   _zz_9934;
  wire       [17:0]   _zz_9935;
  wire       [35:0]   _zz_9936;
  wire       [35:0]   _zz_9937;
  wire       [35:0]   _zz_9938;
  wire       [35:0]   _zz_9939;
  wire       [35:0]   _zz_9940;
  wire       [26:0]   _zz_9941;
  wire       [35:0]   _zz_9942;
  wire       [17:0]   _zz_9943;
  wire       [17:0]   _zz_9944;
  wire       [35:0]   _zz_9945;
  wire       [35:0]   _zz_9946;
  wire       [17:0]   _zz_9947;
  wire       [35:0]   _zz_9948;
  wire       [35:0]   _zz_9949;
  wire       [35:0]   _zz_9950;
  wire       [17:0]   _zz_9951;
  wire       [35:0]   _zz_9952;
  wire       [35:0]   _zz_9953;
  wire       [35:0]   _zz_9954;
  wire       [35:0]   _zz_9955;
  wire       [35:0]   _zz_9956;
  wire       [35:0]   _zz_9957;
  wire       [26:0]   _zz_9958;
  wire       [35:0]   _zz_9959;
  wire       [17:0]   _zz_9960;
  wire       [35:0]   _zz_9961;
  wire       [35:0]   _zz_9962;
  wire       [35:0]   _zz_9963;
  wire       [35:0]   _zz_9964;
  wire       [35:0]   _zz_9965;
  wire       [26:0]   _zz_9966;
  wire       [35:0]   _zz_9967;
  wire       [17:0]   _zz_9968;
  wire       [35:0]   _zz_9969;
  wire       [35:0]   _zz_9970;
  wire       [35:0]   _zz_9971;
  wire       [35:0]   _zz_9972;
  wire       [35:0]   _zz_9973;
  wire       [26:0]   _zz_9974;
  wire       [35:0]   _zz_9975;
  wire       [17:0]   _zz_9976;
  wire       [35:0]   _zz_9977;
  wire       [35:0]   _zz_9978;
  wire       [35:0]   _zz_9979;
  wire       [35:0]   _zz_9980;
  wire       [35:0]   _zz_9981;
  wire       [26:0]   _zz_9982;
  wire       [35:0]   _zz_9983;
  wire       [17:0]   _zz_9984;
  reg        [17:0]   data_in_0_real;
  reg        [17:0]   data_in_0_imag;
  reg        [17:0]   data_in_1_real;
  reg        [17:0]   data_in_1_imag;
  reg        [17:0]   data_in_2_real;
  reg        [17:0]   data_in_2_imag;
  reg        [17:0]   data_in_3_real;
  reg        [17:0]   data_in_3_imag;
  reg        [17:0]   data_in_4_real;
  reg        [17:0]   data_in_4_imag;
  reg        [17:0]   data_in_5_real;
  reg        [17:0]   data_in_5_imag;
  reg        [17:0]   data_in_6_real;
  reg        [17:0]   data_in_6_imag;
  reg        [17:0]   data_in_7_real;
  reg        [17:0]   data_in_7_imag;
  reg        [17:0]   data_in_8_real;
  reg        [17:0]   data_in_8_imag;
  reg        [17:0]   data_in_9_real;
  reg        [17:0]   data_in_9_imag;
  reg        [17:0]   data_in_10_real;
  reg        [17:0]   data_in_10_imag;
  reg        [17:0]   data_in_11_real;
  reg        [17:0]   data_in_11_imag;
  reg        [17:0]   data_in_12_real;
  reg        [17:0]   data_in_12_imag;
  reg        [17:0]   data_in_13_real;
  reg        [17:0]   data_in_13_imag;
  reg        [17:0]   data_in_14_real;
  reg        [17:0]   data_in_14_imag;
  reg        [17:0]   data_in_15_real;
  reg        [17:0]   data_in_15_imag;
  reg        [17:0]   data_in_16_real;
  reg        [17:0]   data_in_16_imag;
  reg        [17:0]   data_in_17_real;
  reg        [17:0]   data_in_17_imag;
  reg        [17:0]   data_in_18_real;
  reg        [17:0]   data_in_18_imag;
  reg        [17:0]   data_in_19_real;
  reg        [17:0]   data_in_19_imag;
  reg        [17:0]   data_in_20_real;
  reg        [17:0]   data_in_20_imag;
  reg        [17:0]   data_in_21_real;
  reg        [17:0]   data_in_21_imag;
  reg        [17:0]   data_in_22_real;
  reg        [17:0]   data_in_22_imag;
  reg        [17:0]   data_in_23_real;
  reg        [17:0]   data_in_23_imag;
  reg        [17:0]   data_in_24_real;
  reg        [17:0]   data_in_24_imag;
  reg        [17:0]   data_in_25_real;
  reg        [17:0]   data_in_25_imag;
  reg        [17:0]   data_in_26_real;
  reg        [17:0]   data_in_26_imag;
  reg        [17:0]   data_in_27_real;
  reg        [17:0]   data_in_27_imag;
  reg        [17:0]   data_in_28_real;
  reg        [17:0]   data_in_28_imag;
  reg        [17:0]   data_in_29_real;
  reg        [17:0]   data_in_29_imag;
  reg        [17:0]   data_in_30_real;
  reg        [17:0]   data_in_30_imag;
  reg        [17:0]   data_in_31_real;
  reg        [17:0]   data_in_31_imag;
  reg        [17:0]   data_in_32_real;
  reg        [17:0]   data_in_32_imag;
  reg        [17:0]   data_in_33_real;
  reg        [17:0]   data_in_33_imag;
  reg        [17:0]   data_in_34_real;
  reg        [17:0]   data_in_34_imag;
  reg        [17:0]   data_in_35_real;
  reg        [17:0]   data_in_35_imag;
  reg        [17:0]   data_in_36_real;
  reg        [17:0]   data_in_36_imag;
  reg        [17:0]   data_in_37_real;
  reg        [17:0]   data_in_37_imag;
  reg        [17:0]   data_in_38_real;
  reg        [17:0]   data_in_38_imag;
  reg        [17:0]   data_in_39_real;
  reg        [17:0]   data_in_39_imag;
  reg        [17:0]   data_in_40_real;
  reg        [17:0]   data_in_40_imag;
  reg        [17:0]   data_in_41_real;
  reg        [17:0]   data_in_41_imag;
  reg        [17:0]   data_in_42_real;
  reg        [17:0]   data_in_42_imag;
  reg        [17:0]   data_in_43_real;
  reg        [17:0]   data_in_43_imag;
  reg        [17:0]   data_in_44_real;
  reg        [17:0]   data_in_44_imag;
  reg        [17:0]   data_in_45_real;
  reg        [17:0]   data_in_45_imag;
  reg        [17:0]   data_in_46_real;
  reg        [17:0]   data_in_46_imag;
  reg        [17:0]   data_in_47_real;
  reg        [17:0]   data_in_47_imag;
  reg        [17:0]   data_in_48_real;
  reg        [17:0]   data_in_48_imag;
  reg        [17:0]   data_in_49_real;
  reg        [17:0]   data_in_49_imag;
  reg        [17:0]   data_in_50_real;
  reg        [17:0]   data_in_50_imag;
  reg        [17:0]   data_in_51_real;
  reg        [17:0]   data_in_51_imag;
  reg        [17:0]   data_in_52_real;
  reg        [17:0]   data_in_52_imag;
  reg        [17:0]   data_in_53_real;
  reg        [17:0]   data_in_53_imag;
  reg        [17:0]   data_in_54_real;
  reg        [17:0]   data_in_54_imag;
  reg        [17:0]   data_in_55_real;
  reg        [17:0]   data_in_55_imag;
  reg        [17:0]   data_in_56_real;
  reg        [17:0]   data_in_56_imag;
  reg        [17:0]   data_in_57_real;
  reg        [17:0]   data_in_57_imag;
  reg        [17:0]   data_in_58_real;
  reg        [17:0]   data_in_58_imag;
  reg        [17:0]   data_in_59_real;
  reg        [17:0]   data_in_59_imag;
  reg        [17:0]   data_in_60_real;
  reg        [17:0]   data_in_60_imag;
  reg        [17:0]   data_in_61_real;
  reg        [17:0]   data_in_61_imag;
  reg        [17:0]   data_in_62_real;
  reg        [17:0]   data_in_62_imag;
  reg        [17:0]   data_in_63_real;
  reg        [17:0]   data_in_63_imag;
  wire       [17:0]   twiddle_factor_table_0_real;
  wire       [17:0]   twiddle_factor_table_0_imag;
  wire       [17:0]   twiddle_factor_table_1_real;
  wire       [17:0]   twiddle_factor_table_1_imag;
  wire       [17:0]   twiddle_factor_table_2_real;
  wire       [17:0]   twiddle_factor_table_2_imag;
  wire       [17:0]   twiddle_factor_table_3_real;
  wire       [17:0]   twiddle_factor_table_3_imag;
  wire       [17:0]   twiddle_factor_table_4_real;
  wire       [17:0]   twiddle_factor_table_4_imag;
  wire       [17:0]   twiddle_factor_table_5_real;
  wire       [17:0]   twiddle_factor_table_5_imag;
  wire       [17:0]   twiddle_factor_table_6_real;
  wire       [17:0]   twiddle_factor_table_6_imag;
  wire       [17:0]   twiddle_factor_table_7_real;
  wire       [17:0]   twiddle_factor_table_7_imag;
  wire       [17:0]   twiddle_factor_table_8_real;
  wire       [17:0]   twiddle_factor_table_8_imag;
  wire       [17:0]   twiddle_factor_table_9_real;
  wire       [17:0]   twiddle_factor_table_9_imag;
  wire       [17:0]   twiddle_factor_table_10_real;
  wire       [17:0]   twiddle_factor_table_10_imag;
  wire       [17:0]   twiddle_factor_table_11_real;
  wire       [17:0]   twiddle_factor_table_11_imag;
  wire       [17:0]   twiddle_factor_table_12_real;
  wire       [17:0]   twiddle_factor_table_12_imag;
  wire       [17:0]   twiddle_factor_table_13_real;
  wire       [17:0]   twiddle_factor_table_13_imag;
  wire       [17:0]   twiddle_factor_table_14_real;
  wire       [17:0]   twiddle_factor_table_14_imag;
  wire       [17:0]   twiddle_factor_table_15_real;
  wire       [17:0]   twiddle_factor_table_15_imag;
  wire       [17:0]   twiddle_factor_table_16_real;
  wire       [17:0]   twiddle_factor_table_16_imag;
  wire       [17:0]   twiddle_factor_table_17_real;
  wire       [17:0]   twiddle_factor_table_17_imag;
  wire       [17:0]   twiddle_factor_table_18_real;
  wire       [17:0]   twiddle_factor_table_18_imag;
  wire       [17:0]   twiddle_factor_table_19_real;
  wire       [17:0]   twiddle_factor_table_19_imag;
  wire       [17:0]   twiddle_factor_table_20_real;
  wire       [17:0]   twiddle_factor_table_20_imag;
  wire       [17:0]   twiddle_factor_table_21_real;
  wire       [17:0]   twiddle_factor_table_21_imag;
  wire       [17:0]   twiddle_factor_table_22_real;
  wire       [17:0]   twiddle_factor_table_22_imag;
  wire       [17:0]   twiddle_factor_table_23_real;
  wire       [17:0]   twiddle_factor_table_23_imag;
  wire       [17:0]   twiddle_factor_table_24_real;
  wire       [17:0]   twiddle_factor_table_24_imag;
  wire       [17:0]   twiddle_factor_table_25_real;
  wire       [17:0]   twiddle_factor_table_25_imag;
  wire       [17:0]   twiddle_factor_table_26_real;
  wire       [17:0]   twiddle_factor_table_26_imag;
  wire       [17:0]   twiddle_factor_table_27_real;
  wire       [17:0]   twiddle_factor_table_27_imag;
  wire       [17:0]   twiddle_factor_table_28_real;
  wire       [17:0]   twiddle_factor_table_28_imag;
  wire       [17:0]   twiddle_factor_table_29_real;
  wire       [17:0]   twiddle_factor_table_29_imag;
  wire       [17:0]   twiddle_factor_table_30_real;
  wire       [17:0]   twiddle_factor_table_30_imag;
  wire       [17:0]   twiddle_factor_table_31_real;
  wire       [17:0]   twiddle_factor_table_31_imag;
  wire       [17:0]   twiddle_factor_table_32_real;
  wire       [17:0]   twiddle_factor_table_32_imag;
  wire       [17:0]   twiddle_factor_table_33_real;
  wire       [17:0]   twiddle_factor_table_33_imag;
  wire       [17:0]   twiddle_factor_table_34_real;
  wire       [17:0]   twiddle_factor_table_34_imag;
  wire       [17:0]   twiddle_factor_table_35_real;
  wire       [17:0]   twiddle_factor_table_35_imag;
  wire       [17:0]   twiddle_factor_table_36_real;
  wire       [17:0]   twiddle_factor_table_36_imag;
  wire       [17:0]   twiddle_factor_table_37_real;
  wire       [17:0]   twiddle_factor_table_37_imag;
  wire       [17:0]   twiddle_factor_table_38_real;
  wire       [17:0]   twiddle_factor_table_38_imag;
  wire       [17:0]   twiddle_factor_table_39_real;
  wire       [17:0]   twiddle_factor_table_39_imag;
  wire       [17:0]   twiddle_factor_table_40_real;
  wire       [17:0]   twiddle_factor_table_40_imag;
  wire       [17:0]   twiddle_factor_table_41_real;
  wire       [17:0]   twiddle_factor_table_41_imag;
  wire       [17:0]   twiddle_factor_table_42_real;
  wire       [17:0]   twiddle_factor_table_42_imag;
  wire       [17:0]   twiddle_factor_table_43_real;
  wire       [17:0]   twiddle_factor_table_43_imag;
  wire       [17:0]   twiddle_factor_table_44_real;
  wire       [17:0]   twiddle_factor_table_44_imag;
  wire       [17:0]   twiddle_factor_table_45_real;
  wire       [17:0]   twiddle_factor_table_45_imag;
  wire       [17:0]   twiddle_factor_table_46_real;
  wire       [17:0]   twiddle_factor_table_46_imag;
  wire       [17:0]   twiddle_factor_table_47_real;
  wire       [17:0]   twiddle_factor_table_47_imag;
  wire       [17:0]   twiddle_factor_table_48_real;
  wire       [17:0]   twiddle_factor_table_48_imag;
  wire       [17:0]   twiddle_factor_table_49_real;
  wire       [17:0]   twiddle_factor_table_49_imag;
  wire       [17:0]   twiddle_factor_table_50_real;
  wire       [17:0]   twiddle_factor_table_50_imag;
  wire       [17:0]   twiddle_factor_table_51_real;
  wire       [17:0]   twiddle_factor_table_51_imag;
  wire       [17:0]   twiddle_factor_table_52_real;
  wire       [17:0]   twiddle_factor_table_52_imag;
  wire       [17:0]   twiddle_factor_table_53_real;
  wire       [17:0]   twiddle_factor_table_53_imag;
  wire       [17:0]   twiddle_factor_table_54_real;
  wire       [17:0]   twiddle_factor_table_54_imag;
  wire       [17:0]   twiddle_factor_table_55_real;
  wire       [17:0]   twiddle_factor_table_55_imag;
  wire       [17:0]   twiddle_factor_table_56_real;
  wire       [17:0]   twiddle_factor_table_56_imag;
  wire       [17:0]   twiddle_factor_table_57_real;
  wire       [17:0]   twiddle_factor_table_57_imag;
  wire       [17:0]   twiddle_factor_table_58_real;
  wire       [17:0]   twiddle_factor_table_58_imag;
  wire       [17:0]   twiddle_factor_table_59_real;
  wire       [17:0]   twiddle_factor_table_59_imag;
  wire       [17:0]   twiddle_factor_table_60_real;
  wire       [17:0]   twiddle_factor_table_60_imag;
  wire       [17:0]   twiddle_factor_table_61_real;
  wire       [17:0]   twiddle_factor_table_61_imag;
  wire       [17:0]   twiddle_factor_table_62_real;
  wire       [17:0]   twiddle_factor_table_62_imag;
  wire       [17:0]   data_reorder_0_real;
  wire       [17:0]   data_reorder_0_imag;
  wire       [17:0]   data_reorder_1_real;
  wire       [17:0]   data_reorder_1_imag;
  wire       [17:0]   data_reorder_2_real;
  wire       [17:0]   data_reorder_2_imag;
  wire       [17:0]   data_reorder_3_real;
  wire       [17:0]   data_reorder_3_imag;
  wire       [17:0]   data_reorder_4_real;
  wire       [17:0]   data_reorder_4_imag;
  wire       [17:0]   data_reorder_5_real;
  wire       [17:0]   data_reorder_5_imag;
  wire       [17:0]   data_reorder_6_real;
  wire       [17:0]   data_reorder_6_imag;
  wire       [17:0]   data_reorder_7_real;
  wire       [17:0]   data_reorder_7_imag;
  wire       [17:0]   data_reorder_8_real;
  wire       [17:0]   data_reorder_8_imag;
  wire       [17:0]   data_reorder_9_real;
  wire       [17:0]   data_reorder_9_imag;
  wire       [17:0]   data_reorder_10_real;
  wire       [17:0]   data_reorder_10_imag;
  wire       [17:0]   data_reorder_11_real;
  wire       [17:0]   data_reorder_11_imag;
  wire       [17:0]   data_reorder_12_real;
  wire       [17:0]   data_reorder_12_imag;
  wire       [17:0]   data_reorder_13_real;
  wire       [17:0]   data_reorder_13_imag;
  wire       [17:0]   data_reorder_14_real;
  wire       [17:0]   data_reorder_14_imag;
  wire       [17:0]   data_reorder_15_real;
  wire       [17:0]   data_reorder_15_imag;
  wire       [17:0]   data_reorder_16_real;
  wire       [17:0]   data_reorder_16_imag;
  wire       [17:0]   data_reorder_17_real;
  wire       [17:0]   data_reorder_17_imag;
  wire       [17:0]   data_reorder_18_real;
  wire       [17:0]   data_reorder_18_imag;
  wire       [17:0]   data_reorder_19_real;
  wire       [17:0]   data_reorder_19_imag;
  wire       [17:0]   data_reorder_20_real;
  wire       [17:0]   data_reorder_20_imag;
  wire       [17:0]   data_reorder_21_real;
  wire       [17:0]   data_reorder_21_imag;
  wire       [17:0]   data_reorder_22_real;
  wire       [17:0]   data_reorder_22_imag;
  wire       [17:0]   data_reorder_23_real;
  wire       [17:0]   data_reorder_23_imag;
  wire       [17:0]   data_reorder_24_real;
  wire       [17:0]   data_reorder_24_imag;
  wire       [17:0]   data_reorder_25_real;
  wire       [17:0]   data_reorder_25_imag;
  wire       [17:0]   data_reorder_26_real;
  wire       [17:0]   data_reorder_26_imag;
  wire       [17:0]   data_reorder_27_real;
  wire       [17:0]   data_reorder_27_imag;
  wire       [17:0]   data_reorder_28_real;
  wire       [17:0]   data_reorder_28_imag;
  wire       [17:0]   data_reorder_29_real;
  wire       [17:0]   data_reorder_29_imag;
  wire       [17:0]   data_reorder_30_real;
  wire       [17:0]   data_reorder_30_imag;
  wire       [17:0]   data_reorder_31_real;
  wire       [17:0]   data_reorder_31_imag;
  wire       [17:0]   data_reorder_32_real;
  wire       [17:0]   data_reorder_32_imag;
  wire       [17:0]   data_reorder_33_real;
  wire       [17:0]   data_reorder_33_imag;
  wire       [17:0]   data_reorder_34_real;
  wire       [17:0]   data_reorder_34_imag;
  wire       [17:0]   data_reorder_35_real;
  wire       [17:0]   data_reorder_35_imag;
  wire       [17:0]   data_reorder_36_real;
  wire       [17:0]   data_reorder_36_imag;
  wire       [17:0]   data_reorder_37_real;
  wire       [17:0]   data_reorder_37_imag;
  wire       [17:0]   data_reorder_38_real;
  wire       [17:0]   data_reorder_38_imag;
  wire       [17:0]   data_reorder_39_real;
  wire       [17:0]   data_reorder_39_imag;
  wire       [17:0]   data_reorder_40_real;
  wire       [17:0]   data_reorder_40_imag;
  wire       [17:0]   data_reorder_41_real;
  wire       [17:0]   data_reorder_41_imag;
  wire       [17:0]   data_reorder_42_real;
  wire       [17:0]   data_reorder_42_imag;
  wire       [17:0]   data_reorder_43_real;
  wire       [17:0]   data_reorder_43_imag;
  wire       [17:0]   data_reorder_44_real;
  wire       [17:0]   data_reorder_44_imag;
  wire       [17:0]   data_reorder_45_real;
  wire       [17:0]   data_reorder_45_imag;
  wire       [17:0]   data_reorder_46_real;
  wire       [17:0]   data_reorder_46_imag;
  wire       [17:0]   data_reorder_47_real;
  wire       [17:0]   data_reorder_47_imag;
  wire       [17:0]   data_reorder_48_real;
  wire       [17:0]   data_reorder_48_imag;
  wire       [17:0]   data_reorder_49_real;
  wire       [17:0]   data_reorder_49_imag;
  wire       [17:0]   data_reorder_50_real;
  wire       [17:0]   data_reorder_50_imag;
  wire       [17:0]   data_reorder_51_real;
  wire       [17:0]   data_reorder_51_imag;
  wire       [17:0]   data_reorder_52_real;
  wire       [17:0]   data_reorder_52_imag;
  wire       [17:0]   data_reorder_53_real;
  wire       [17:0]   data_reorder_53_imag;
  wire       [17:0]   data_reorder_54_real;
  wire       [17:0]   data_reorder_54_imag;
  wire       [17:0]   data_reorder_55_real;
  wire       [17:0]   data_reorder_55_imag;
  wire       [17:0]   data_reorder_56_real;
  wire       [17:0]   data_reorder_56_imag;
  wire       [17:0]   data_reorder_57_real;
  wire       [17:0]   data_reorder_57_imag;
  wire       [17:0]   data_reorder_58_real;
  wire       [17:0]   data_reorder_58_imag;
  wire       [17:0]   data_reorder_59_real;
  wire       [17:0]   data_reorder_59_imag;
  wire       [17:0]   data_reorder_60_real;
  wire       [17:0]   data_reorder_60_imag;
  wire       [17:0]   data_reorder_61_real;
  wire       [17:0]   data_reorder_61_imag;
  wire       [17:0]   data_reorder_62_real;
  wire       [17:0]   data_reorder_62_imag;
  wire       [17:0]   data_reorder_63_real;
  wire       [17:0]   data_reorder_63_imag;
  reg        [17:0]   data_mid_0_0_real;
  reg        [17:0]   data_mid_0_0_imag;
  reg        [17:0]   data_mid_0_1_real;
  reg        [17:0]   data_mid_0_1_imag;
  reg        [17:0]   data_mid_0_2_real;
  reg        [17:0]   data_mid_0_2_imag;
  reg        [17:0]   data_mid_0_3_real;
  reg        [17:0]   data_mid_0_3_imag;
  reg        [17:0]   data_mid_0_4_real;
  reg        [17:0]   data_mid_0_4_imag;
  reg        [17:0]   data_mid_0_5_real;
  reg        [17:0]   data_mid_0_5_imag;
  reg        [17:0]   data_mid_0_6_real;
  reg        [17:0]   data_mid_0_6_imag;
  reg        [17:0]   data_mid_0_7_real;
  reg        [17:0]   data_mid_0_7_imag;
  reg        [17:0]   data_mid_0_8_real;
  reg        [17:0]   data_mid_0_8_imag;
  reg        [17:0]   data_mid_0_9_real;
  reg        [17:0]   data_mid_0_9_imag;
  reg        [17:0]   data_mid_0_10_real;
  reg        [17:0]   data_mid_0_10_imag;
  reg        [17:0]   data_mid_0_11_real;
  reg        [17:0]   data_mid_0_11_imag;
  reg        [17:0]   data_mid_0_12_real;
  reg        [17:0]   data_mid_0_12_imag;
  reg        [17:0]   data_mid_0_13_real;
  reg        [17:0]   data_mid_0_13_imag;
  reg        [17:0]   data_mid_0_14_real;
  reg        [17:0]   data_mid_0_14_imag;
  reg        [17:0]   data_mid_0_15_real;
  reg        [17:0]   data_mid_0_15_imag;
  reg        [17:0]   data_mid_0_16_real;
  reg        [17:0]   data_mid_0_16_imag;
  reg        [17:0]   data_mid_0_17_real;
  reg        [17:0]   data_mid_0_17_imag;
  reg        [17:0]   data_mid_0_18_real;
  reg        [17:0]   data_mid_0_18_imag;
  reg        [17:0]   data_mid_0_19_real;
  reg        [17:0]   data_mid_0_19_imag;
  reg        [17:0]   data_mid_0_20_real;
  reg        [17:0]   data_mid_0_20_imag;
  reg        [17:0]   data_mid_0_21_real;
  reg        [17:0]   data_mid_0_21_imag;
  reg        [17:0]   data_mid_0_22_real;
  reg        [17:0]   data_mid_0_22_imag;
  reg        [17:0]   data_mid_0_23_real;
  reg        [17:0]   data_mid_0_23_imag;
  reg        [17:0]   data_mid_0_24_real;
  reg        [17:0]   data_mid_0_24_imag;
  reg        [17:0]   data_mid_0_25_real;
  reg        [17:0]   data_mid_0_25_imag;
  reg        [17:0]   data_mid_0_26_real;
  reg        [17:0]   data_mid_0_26_imag;
  reg        [17:0]   data_mid_0_27_real;
  reg        [17:0]   data_mid_0_27_imag;
  reg        [17:0]   data_mid_0_28_real;
  reg        [17:0]   data_mid_0_28_imag;
  reg        [17:0]   data_mid_0_29_real;
  reg        [17:0]   data_mid_0_29_imag;
  reg        [17:0]   data_mid_0_30_real;
  reg        [17:0]   data_mid_0_30_imag;
  reg        [17:0]   data_mid_0_31_real;
  reg        [17:0]   data_mid_0_31_imag;
  reg        [17:0]   data_mid_0_32_real;
  reg        [17:0]   data_mid_0_32_imag;
  reg        [17:0]   data_mid_0_33_real;
  reg        [17:0]   data_mid_0_33_imag;
  reg        [17:0]   data_mid_0_34_real;
  reg        [17:0]   data_mid_0_34_imag;
  reg        [17:0]   data_mid_0_35_real;
  reg        [17:0]   data_mid_0_35_imag;
  reg        [17:0]   data_mid_0_36_real;
  reg        [17:0]   data_mid_0_36_imag;
  reg        [17:0]   data_mid_0_37_real;
  reg        [17:0]   data_mid_0_37_imag;
  reg        [17:0]   data_mid_0_38_real;
  reg        [17:0]   data_mid_0_38_imag;
  reg        [17:0]   data_mid_0_39_real;
  reg        [17:0]   data_mid_0_39_imag;
  reg        [17:0]   data_mid_0_40_real;
  reg        [17:0]   data_mid_0_40_imag;
  reg        [17:0]   data_mid_0_41_real;
  reg        [17:0]   data_mid_0_41_imag;
  reg        [17:0]   data_mid_0_42_real;
  reg        [17:0]   data_mid_0_42_imag;
  reg        [17:0]   data_mid_0_43_real;
  reg        [17:0]   data_mid_0_43_imag;
  reg        [17:0]   data_mid_0_44_real;
  reg        [17:0]   data_mid_0_44_imag;
  reg        [17:0]   data_mid_0_45_real;
  reg        [17:0]   data_mid_0_45_imag;
  reg        [17:0]   data_mid_0_46_real;
  reg        [17:0]   data_mid_0_46_imag;
  reg        [17:0]   data_mid_0_47_real;
  reg        [17:0]   data_mid_0_47_imag;
  reg        [17:0]   data_mid_0_48_real;
  reg        [17:0]   data_mid_0_48_imag;
  reg        [17:0]   data_mid_0_49_real;
  reg        [17:0]   data_mid_0_49_imag;
  reg        [17:0]   data_mid_0_50_real;
  reg        [17:0]   data_mid_0_50_imag;
  reg        [17:0]   data_mid_0_51_real;
  reg        [17:0]   data_mid_0_51_imag;
  reg        [17:0]   data_mid_0_52_real;
  reg        [17:0]   data_mid_0_52_imag;
  reg        [17:0]   data_mid_0_53_real;
  reg        [17:0]   data_mid_0_53_imag;
  reg        [17:0]   data_mid_0_54_real;
  reg        [17:0]   data_mid_0_54_imag;
  reg        [17:0]   data_mid_0_55_real;
  reg        [17:0]   data_mid_0_55_imag;
  reg        [17:0]   data_mid_0_56_real;
  reg        [17:0]   data_mid_0_56_imag;
  reg        [17:0]   data_mid_0_57_real;
  reg        [17:0]   data_mid_0_57_imag;
  reg        [17:0]   data_mid_0_58_real;
  reg        [17:0]   data_mid_0_58_imag;
  reg        [17:0]   data_mid_0_59_real;
  reg        [17:0]   data_mid_0_59_imag;
  reg        [17:0]   data_mid_0_60_real;
  reg        [17:0]   data_mid_0_60_imag;
  reg        [17:0]   data_mid_0_61_real;
  reg        [17:0]   data_mid_0_61_imag;
  reg        [17:0]   data_mid_0_62_real;
  reg        [17:0]   data_mid_0_62_imag;
  reg        [17:0]   data_mid_0_63_real;
  reg        [17:0]   data_mid_0_63_imag;
  reg        [17:0]   data_mid_1_0_real;
  reg        [17:0]   data_mid_1_0_imag;
  reg        [17:0]   data_mid_1_1_real;
  reg        [17:0]   data_mid_1_1_imag;
  reg        [17:0]   data_mid_1_2_real;
  reg        [17:0]   data_mid_1_2_imag;
  reg        [17:0]   data_mid_1_3_real;
  reg        [17:0]   data_mid_1_3_imag;
  reg        [17:0]   data_mid_1_4_real;
  reg        [17:0]   data_mid_1_4_imag;
  reg        [17:0]   data_mid_1_5_real;
  reg        [17:0]   data_mid_1_5_imag;
  reg        [17:0]   data_mid_1_6_real;
  reg        [17:0]   data_mid_1_6_imag;
  reg        [17:0]   data_mid_1_7_real;
  reg        [17:0]   data_mid_1_7_imag;
  reg        [17:0]   data_mid_1_8_real;
  reg        [17:0]   data_mid_1_8_imag;
  reg        [17:0]   data_mid_1_9_real;
  reg        [17:0]   data_mid_1_9_imag;
  reg        [17:0]   data_mid_1_10_real;
  reg        [17:0]   data_mid_1_10_imag;
  reg        [17:0]   data_mid_1_11_real;
  reg        [17:0]   data_mid_1_11_imag;
  reg        [17:0]   data_mid_1_12_real;
  reg        [17:0]   data_mid_1_12_imag;
  reg        [17:0]   data_mid_1_13_real;
  reg        [17:0]   data_mid_1_13_imag;
  reg        [17:0]   data_mid_1_14_real;
  reg        [17:0]   data_mid_1_14_imag;
  reg        [17:0]   data_mid_1_15_real;
  reg        [17:0]   data_mid_1_15_imag;
  reg        [17:0]   data_mid_1_16_real;
  reg        [17:0]   data_mid_1_16_imag;
  reg        [17:0]   data_mid_1_17_real;
  reg        [17:0]   data_mid_1_17_imag;
  reg        [17:0]   data_mid_1_18_real;
  reg        [17:0]   data_mid_1_18_imag;
  reg        [17:0]   data_mid_1_19_real;
  reg        [17:0]   data_mid_1_19_imag;
  reg        [17:0]   data_mid_1_20_real;
  reg        [17:0]   data_mid_1_20_imag;
  reg        [17:0]   data_mid_1_21_real;
  reg        [17:0]   data_mid_1_21_imag;
  reg        [17:0]   data_mid_1_22_real;
  reg        [17:0]   data_mid_1_22_imag;
  reg        [17:0]   data_mid_1_23_real;
  reg        [17:0]   data_mid_1_23_imag;
  reg        [17:0]   data_mid_1_24_real;
  reg        [17:0]   data_mid_1_24_imag;
  reg        [17:0]   data_mid_1_25_real;
  reg        [17:0]   data_mid_1_25_imag;
  reg        [17:0]   data_mid_1_26_real;
  reg        [17:0]   data_mid_1_26_imag;
  reg        [17:0]   data_mid_1_27_real;
  reg        [17:0]   data_mid_1_27_imag;
  reg        [17:0]   data_mid_1_28_real;
  reg        [17:0]   data_mid_1_28_imag;
  reg        [17:0]   data_mid_1_29_real;
  reg        [17:0]   data_mid_1_29_imag;
  reg        [17:0]   data_mid_1_30_real;
  reg        [17:0]   data_mid_1_30_imag;
  reg        [17:0]   data_mid_1_31_real;
  reg        [17:0]   data_mid_1_31_imag;
  reg        [17:0]   data_mid_1_32_real;
  reg        [17:0]   data_mid_1_32_imag;
  reg        [17:0]   data_mid_1_33_real;
  reg        [17:0]   data_mid_1_33_imag;
  reg        [17:0]   data_mid_1_34_real;
  reg        [17:0]   data_mid_1_34_imag;
  reg        [17:0]   data_mid_1_35_real;
  reg        [17:0]   data_mid_1_35_imag;
  reg        [17:0]   data_mid_1_36_real;
  reg        [17:0]   data_mid_1_36_imag;
  reg        [17:0]   data_mid_1_37_real;
  reg        [17:0]   data_mid_1_37_imag;
  reg        [17:0]   data_mid_1_38_real;
  reg        [17:0]   data_mid_1_38_imag;
  reg        [17:0]   data_mid_1_39_real;
  reg        [17:0]   data_mid_1_39_imag;
  reg        [17:0]   data_mid_1_40_real;
  reg        [17:0]   data_mid_1_40_imag;
  reg        [17:0]   data_mid_1_41_real;
  reg        [17:0]   data_mid_1_41_imag;
  reg        [17:0]   data_mid_1_42_real;
  reg        [17:0]   data_mid_1_42_imag;
  reg        [17:0]   data_mid_1_43_real;
  reg        [17:0]   data_mid_1_43_imag;
  reg        [17:0]   data_mid_1_44_real;
  reg        [17:0]   data_mid_1_44_imag;
  reg        [17:0]   data_mid_1_45_real;
  reg        [17:0]   data_mid_1_45_imag;
  reg        [17:0]   data_mid_1_46_real;
  reg        [17:0]   data_mid_1_46_imag;
  reg        [17:0]   data_mid_1_47_real;
  reg        [17:0]   data_mid_1_47_imag;
  reg        [17:0]   data_mid_1_48_real;
  reg        [17:0]   data_mid_1_48_imag;
  reg        [17:0]   data_mid_1_49_real;
  reg        [17:0]   data_mid_1_49_imag;
  reg        [17:0]   data_mid_1_50_real;
  reg        [17:0]   data_mid_1_50_imag;
  reg        [17:0]   data_mid_1_51_real;
  reg        [17:0]   data_mid_1_51_imag;
  reg        [17:0]   data_mid_1_52_real;
  reg        [17:0]   data_mid_1_52_imag;
  reg        [17:0]   data_mid_1_53_real;
  reg        [17:0]   data_mid_1_53_imag;
  reg        [17:0]   data_mid_1_54_real;
  reg        [17:0]   data_mid_1_54_imag;
  reg        [17:0]   data_mid_1_55_real;
  reg        [17:0]   data_mid_1_55_imag;
  reg        [17:0]   data_mid_1_56_real;
  reg        [17:0]   data_mid_1_56_imag;
  reg        [17:0]   data_mid_1_57_real;
  reg        [17:0]   data_mid_1_57_imag;
  reg        [17:0]   data_mid_1_58_real;
  reg        [17:0]   data_mid_1_58_imag;
  reg        [17:0]   data_mid_1_59_real;
  reg        [17:0]   data_mid_1_59_imag;
  reg        [17:0]   data_mid_1_60_real;
  reg        [17:0]   data_mid_1_60_imag;
  reg        [17:0]   data_mid_1_61_real;
  reg        [17:0]   data_mid_1_61_imag;
  reg        [17:0]   data_mid_1_62_real;
  reg        [17:0]   data_mid_1_62_imag;
  reg        [17:0]   data_mid_1_63_real;
  reg        [17:0]   data_mid_1_63_imag;
  reg        [17:0]   data_mid_2_0_real;
  reg        [17:0]   data_mid_2_0_imag;
  reg        [17:0]   data_mid_2_1_real;
  reg        [17:0]   data_mid_2_1_imag;
  reg        [17:0]   data_mid_2_2_real;
  reg        [17:0]   data_mid_2_2_imag;
  reg        [17:0]   data_mid_2_3_real;
  reg        [17:0]   data_mid_2_3_imag;
  reg        [17:0]   data_mid_2_4_real;
  reg        [17:0]   data_mid_2_4_imag;
  reg        [17:0]   data_mid_2_5_real;
  reg        [17:0]   data_mid_2_5_imag;
  reg        [17:0]   data_mid_2_6_real;
  reg        [17:0]   data_mid_2_6_imag;
  reg        [17:0]   data_mid_2_7_real;
  reg        [17:0]   data_mid_2_7_imag;
  reg        [17:0]   data_mid_2_8_real;
  reg        [17:0]   data_mid_2_8_imag;
  reg        [17:0]   data_mid_2_9_real;
  reg        [17:0]   data_mid_2_9_imag;
  reg        [17:0]   data_mid_2_10_real;
  reg        [17:0]   data_mid_2_10_imag;
  reg        [17:0]   data_mid_2_11_real;
  reg        [17:0]   data_mid_2_11_imag;
  reg        [17:0]   data_mid_2_12_real;
  reg        [17:0]   data_mid_2_12_imag;
  reg        [17:0]   data_mid_2_13_real;
  reg        [17:0]   data_mid_2_13_imag;
  reg        [17:0]   data_mid_2_14_real;
  reg        [17:0]   data_mid_2_14_imag;
  reg        [17:0]   data_mid_2_15_real;
  reg        [17:0]   data_mid_2_15_imag;
  reg        [17:0]   data_mid_2_16_real;
  reg        [17:0]   data_mid_2_16_imag;
  reg        [17:0]   data_mid_2_17_real;
  reg        [17:0]   data_mid_2_17_imag;
  reg        [17:0]   data_mid_2_18_real;
  reg        [17:0]   data_mid_2_18_imag;
  reg        [17:0]   data_mid_2_19_real;
  reg        [17:0]   data_mid_2_19_imag;
  reg        [17:0]   data_mid_2_20_real;
  reg        [17:0]   data_mid_2_20_imag;
  reg        [17:0]   data_mid_2_21_real;
  reg        [17:0]   data_mid_2_21_imag;
  reg        [17:0]   data_mid_2_22_real;
  reg        [17:0]   data_mid_2_22_imag;
  reg        [17:0]   data_mid_2_23_real;
  reg        [17:0]   data_mid_2_23_imag;
  reg        [17:0]   data_mid_2_24_real;
  reg        [17:0]   data_mid_2_24_imag;
  reg        [17:0]   data_mid_2_25_real;
  reg        [17:0]   data_mid_2_25_imag;
  reg        [17:0]   data_mid_2_26_real;
  reg        [17:0]   data_mid_2_26_imag;
  reg        [17:0]   data_mid_2_27_real;
  reg        [17:0]   data_mid_2_27_imag;
  reg        [17:0]   data_mid_2_28_real;
  reg        [17:0]   data_mid_2_28_imag;
  reg        [17:0]   data_mid_2_29_real;
  reg        [17:0]   data_mid_2_29_imag;
  reg        [17:0]   data_mid_2_30_real;
  reg        [17:0]   data_mid_2_30_imag;
  reg        [17:0]   data_mid_2_31_real;
  reg        [17:0]   data_mid_2_31_imag;
  reg        [17:0]   data_mid_2_32_real;
  reg        [17:0]   data_mid_2_32_imag;
  reg        [17:0]   data_mid_2_33_real;
  reg        [17:0]   data_mid_2_33_imag;
  reg        [17:0]   data_mid_2_34_real;
  reg        [17:0]   data_mid_2_34_imag;
  reg        [17:0]   data_mid_2_35_real;
  reg        [17:0]   data_mid_2_35_imag;
  reg        [17:0]   data_mid_2_36_real;
  reg        [17:0]   data_mid_2_36_imag;
  reg        [17:0]   data_mid_2_37_real;
  reg        [17:0]   data_mid_2_37_imag;
  reg        [17:0]   data_mid_2_38_real;
  reg        [17:0]   data_mid_2_38_imag;
  reg        [17:0]   data_mid_2_39_real;
  reg        [17:0]   data_mid_2_39_imag;
  reg        [17:0]   data_mid_2_40_real;
  reg        [17:0]   data_mid_2_40_imag;
  reg        [17:0]   data_mid_2_41_real;
  reg        [17:0]   data_mid_2_41_imag;
  reg        [17:0]   data_mid_2_42_real;
  reg        [17:0]   data_mid_2_42_imag;
  reg        [17:0]   data_mid_2_43_real;
  reg        [17:0]   data_mid_2_43_imag;
  reg        [17:0]   data_mid_2_44_real;
  reg        [17:0]   data_mid_2_44_imag;
  reg        [17:0]   data_mid_2_45_real;
  reg        [17:0]   data_mid_2_45_imag;
  reg        [17:0]   data_mid_2_46_real;
  reg        [17:0]   data_mid_2_46_imag;
  reg        [17:0]   data_mid_2_47_real;
  reg        [17:0]   data_mid_2_47_imag;
  reg        [17:0]   data_mid_2_48_real;
  reg        [17:0]   data_mid_2_48_imag;
  reg        [17:0]   data_mid_2_49_real;
  reg        [17:0]   data_mid_2_49_imag;
  reg        [17:0]   data_mid_2_50_real;
  reg        [17:0]   data_mid_2_50_imag;
  reg        [17:0]   data_mid_2_51_real;
  reg        [17:0]   data_mid_2_51_imag;
  reg        [17:0]   data_mid_2_52_real;
  reg        [17:0]   data_mid_2_52_imag;
  reg        [17:0]   data_mid_2_53_real;
  reg        [17:0]   data_mid_2_53_imag;
  reg        [17:0]   data_mid_2_54_real;
  reg        [17:0]   data_mid_2_54_imag;
  reg        [17:0]   data_mid_2_55_real;
  reg        [17:0]   data_mid_2_55_imag;
  reg        [17:0]   data_mid_2_56_real;
  reg        [17:0]   data_mid_2_56_imag;
  reg        [17:0]   data_mid_2_57_real;
  reg        [17:0]   data_mid_2_57_imag;
  reg        [17:0]   data_mid_2_58_real;
  reg        [17:0]   data_mid_2_58_imag;
  reg        [17:0]   data_mid_2_59_real;
  reg        [17:0]   data_mid_2_59_imag;
  reg        [17:0]   data_mid_2_60_real;
  reg        [17:0]   data_mid_2_60_imag;
  reg        [17:0]   data_mid_2_61_real;
  reg        [17:0]   data_mid_2_61_imag;
  reg        [17:0]   data_mid_2_62_real;
  reg        [17:0]   data_mid_2_62_imag;
  reg        [17:0]   data_mid_2_63_real;
  reg        [17:0]   data_mid_2_63_imag;
  reg        [17:0]   data_mid_3_0_real;
  reg        [17:0]   data_mid_3_0_imag;
  reg        [17:0]   data_mid_3_1_real;
  reg        [17:0]   data_mid_3_1_imag;
  reg        [17:0]   data_mid_3_2_real;
  reg        [17:0]   data_mid_3_2_imag;
  reg        [17:0]   data_mid_3_3_real;
  reg        [17:0]   data_mid_3_3_imag;
  reg        [17:0]   data_mid_3_4_real;
  reg        [17:0]   data_mid_3_4_imag;
  reg        [17:0]   data_mid_3_5_real;
  reg        [17:0]   data_mid_3_5_imag;
  reg        [17:0]   data_mid_3_6_real;
  reg        [17:0]   data_mid_3_6_imag;
  reg        [17:0]   data_mid_3_7_real;
  reg        [17:0]   data_mid_3_7_imag;
  reg        [17:0]   data_mid_3_8_real;
  reg        [17:0]   data_mid_3_8_imag;
  reg        [17:0]   data_mid_3_9_real;
  reg        [17:0]   data_mid_3_9_imag;
  reg        [17:0]   data_mid_3_10_real;
  reg        [17:0]   data_mid_3_10_imag;
  reg        [17:0]   data_mid_3_11_real;
  reg        [17:0]   data_mid_3_11_imag;
  reg        [17:0]   data_mid_3_12_real;
  reg        [17:0]   data_mid_3_12_imag;
  reg        [17:0]   data_mid_3_13_real;
  reg        [17:0]   data_mid_3_13_imag;
  reg        [17:0]   data_mid_3_14_real;
  reg        [17:0]   data_mid_3_14_imag;
  reg        [17:0]   data_mid_3_15_real;
  reg        [17:0]   data_mid_3_15_imag;
  reg        [17:0]   data_mid_3_16_real;
  reg        [17:0]   data_mid_3_16_imag;
  reg        [17:0]   data_mid_3_17_real;
  reg        [17:0]   data_mid_3_17_imag;
  reg        [17:0]   data_mid_3_18_real;
  reg        [17:0]   data_mid_3_18_imag;
  reg        [17:0]   data_mid_3_19_real;
  reg        [17:0]   data_mid_3_19_imag;
  reg        [17:0]   data_mid_3_20_real;
  reg        [17:0]   data_mid_3_20_imag;
  reg        [17:0]   data_mid_3_21_real;
  reg        [17:0]   data_mid_3_21_imag;
  reg        [17:0]   data_mid_3_22_real;
  reg        [17:0]   data_mid_3_22_imag;
  reg        [17:0]   data_mid_3_23_real;
  reg        [17:0]   data_mid_3_23_imag;
  reg        [17:0]   data_mid_3_24_real;
  reg        [17:0]   data_mid_3_24_imag;
  reg        [17:0]   data_mid_3_25_real;
  reg        [17:0]   data_mid_3_25_imag;
  reg        [17:0]   data_mid_3_26_real;
  reg        [17:0]   data_mid_3_26_imag;
  reg        [17:0]   data_mid_3_27_real;
  reg        [17:0]   data_mid_3_27_imag;
  reg        [17:0]   data_mid_3_28_real;
  reg        [17:0]   data_mid_3_28_imag;
  reg        [17:0]   data_mid_3_29_real;
  reg        [17:0]   data_mid_3_29_imag;
  reg        [17:0]   data_mid_3_30_real;
  reg        [17:0]   data_mid_3_30_imag;
  reg        [17:0]   data_mid_3_31_real;
  reg        [17:0]   data_mid_3_31_imag;
  reg        [17:0]   data_mid_3_32_real;
  reg        [17:0]   data_mid_3_32_imag;
  reg        [17:0]   data_mid_3_33_real;
  reg        [17:0]   data_mid_3_33_imag;
  reg        [17:0]   data_mid_3_34_real;
  reg        [17:0]   data_mid_3_34_imag;
  reg        [17:0]   data_mid_3_35_real;
  reg        [17:0]   data_mid_3_35_imag;
  reg        [17:0]   data_mid_3_36_real;
  reg        [17:0]   data_mid_3_36_imag;
  reg        [17:0]   data_mid_3_37_real;
  reg        [17:0]   data_mid_3_37_imag;
  reg        [17:0]   data_mid_3_38_real;
  reg        [17:0]   data_mid_3_38_imag;
  reg        [17:0]   data_mid_3_39_real;
  reg        [17:0]   data_mid_3_39_imag;
  reg        [17:0]   data_mid_3_40_real;
  reg        [17:0]   data_mid_3_40_imag;
  reg        [17:0]   data_mid_3_41_real;
  reg        [17:0]   data_mid_3_41_imag;
  reg        [17:0]   data_mid_3_42_real;
  reg        [17:0]   data_mid_3_42_imag;
  reg        [17:0]   data_mid_3_43_real;
  reg        [17:0]   data_mid_3_43_imag;
  reg        [17:0]   data_mid_3_44_real;
  reg        [17:0]   data_mid_3_44_imag;
  reg        [17:0]   data_mid_3_45_real;
  reg        [17:0]   data_mid_3_45_imag;
  reg        [17:0]   data_mid_3_46_real;
  reg        [17:0]   data_mid_3_46_imag;
  reg        [17:0]   data_mid_3_47_real;
  reg        [17:0]   data_mid_3_47_imag;
  reg        [17:0]   data_mid_3_48_real;
  reg        [17:0]   data_mid_3_48_imag;
  reg        [17:0]   data_mid_3_49_real;
  reg        [17:0]   data_mid_3_49_imag;
  reg        [17:0]   data_mid_3_50_real;
  reg        [17:0]   data_mid_3_50_imag;
  reg        [17:0]   data_mid_3_51_real;
  reg        [17:0]   data_mid_3_51_imag;
  reg        [17:0]   data_mid_3_52_real;
  reg        [17:0]   data_mid_3_52_imag;
  reg        [17:0]   data_mid_3_53_real;
  reg        [17:0]   data_mid_3_53_imag;
  reg        [17:0]   data_mid_3_54_real;
  reg        [17:0]   data_mid_3_54_imag;
  reg        [17:0]   data_mid_3_55_real;
  reg        [17:0]   data_mid_3_55_imag;
  reg        [17:0]   data_mid_3_56_real;
  reg        [17:0]   data_mid_3_56_imag;
  reg        [17:0]   data_mid_3_57_real;
  reg        [17:0]   data_mid_3_57_imag;
  reg        [17:0]   data_mid_3_58_real;
  reg        [17:0]   data_mid_3_58_imag;
  reg        [17:0]   data_mid_3_59_real;
  reg        [17:0]   data_mid_3_59_imag;
  reg        [17:0]   data_mid_3_60_real;
  reg        [17:0]   data_mid_3_60_imag;
  reg        [17:0]   data_mid_3_61_real;
  reg        [17:0]   data_mid_3_61_imag;
  reg        [17:0]   data_mid_3_62_real;
  reg        [17:0]   data_mid_3_62_imag;
  reg        [17:0]   data_mid_3_63_real;
  reg        [17:0]   data_mid_3_63_imag;
  reg        [17:0]   data_mid_4_0_real;
  reg        [17:0]   data_mid_4_0_imag;
  reg        [17:0]   data_mid_4_1_real;
  reg        [17:0]   data_mid_4_1_imag;
  reg        [17:0]   data_mid_4_2_real;
  reg        [17:0]   data_mid_4_2_imag;
  reg        [17:0]   data_mid_4_3_real;
  reg        [17:0]   data_mid_4_3_imag;
  reg        [17:0]   data_mid_4_4_real;
  reg        [17:0]   data_mid_4_4_imag;
  reg        [17:0]   data_mid_4_5_real;
  reg        [17:0]   data_mid_4_5_imag;
  reg        [17:0]   data_mid_4_6_real;
  reg        [17:0]   data_mid_4_6_imag;
  reg        [17:0]   data_mid_4_7_real;
  reg        [17:0]   data_mid_4_7_imag;
  reg        [17:0]   data_mid_4_8_real;
  reg        [17:0]   data_mid_4_8_imag;
  reg        [17:0]   data_mid_4_9_real;
  reg        [17:0]   data_mid_4_9_imag;
  reg        [17:0]   data_mid_4_10_real;
  reg        [17:0]   data_mid_4_10_imag;
  reg        [17:0]   data_mid_4_11_real;
  reg        [17:0]   data_mid_4_11_imag;
  reg        [17:0]   data_mid_4_12_real;
  reg        [17:0]   data_mid_4_12_imag;
  reg        [17:0]   data_mid_4_13_real;
  reg        [17:0]   data_mid_4_13_imag;
  reg        [17:0]   data_mid_4_14_real;
  reg        [17:0]   data_mid_4_14_imag;
  reg        [17:0]   data_mid_4_15_real;
  reg        [17:0]   data_mid_4_15_imag;
  reg        [17:0]   data_mid_4_16_real;
  reg        [17:0]   data_mid_4_16_imag;
  reg        [17:0]   data_mid_4_17_real;
  reg        [17:0]   data_mid_4_17_imag;
  reg        [17:0]   data_mid_4_18_real;
  reg        [17:0]   data_mid_4_18_imag;
  reg        [17:0]   data_mid_4_19_real;
  reg        [17:0]   data_mid_4_19_imag;
  reg        [17:0]   data_mid_4_20_real;
  reg        [17:0]   data_mid_4_20_imag;
  reg        [17:0]   data_mid_4_21_real;
  reg        [17:0]   data_mid_4_21_imag;
  reg        [17:0]   data_mid_4_22_real;
  reg        [17:0]   data_mid_4_22_imag;
  reg        [17:0]   data_mid_4_23_real;
  reg        [17:0]   data_mid_4_23_imag;
  reg        [17:0]   data_mid_4_24_real;
  reg        [17:0]   data_mid_4_24_imag;
  reg        [17:0]   data_mid_4_25_real;
  reg        [17:0]   data_mid_4_25_imag;
  reg        [17:0]   data_mid_4_26_real;
  reg        [17:0]   data_mid_4_26_imag;
  reg        [17:0]   data_mid_4_27_real;
  reg        [17:0]   data_mid_4_27_imag;
  reg        [17:0]   data_mid_4_28_real;
  reg        [17:0]   data_mid_4_28_imag;
  reg        [17:0]   data_mid_4_29_real;
  reg        [17:0]   data_mid_4_29_imag;
  reg        [17:0]   data_mid_4_30_real;
  reg        [17:0]   data_mid_4_30_imag;
  reg        [17:0]   data_mid_4_31_real;
  reg        [17:0]   data_mid_4_31_imag;
  reg        [17:0]   data_mid_4_32_real;
  reg        [17:0]   data_mid_4_32_imag;
  reg        [17:0]   data_mid_4_33_real;
  reg        [17:0]   data_mid_4_33_imag;
  reg        [17:0]   data_mid_4_34_real;
  reg        [17:0]   data_mid_4_34_imag;
  reg        [17:0]   data_mid_4_35_real;
  reg        [17:0]   data_mid_4_35_imag;
  reg        [17:0]   data_mid_4_36_real;
  reg        [17:0]   data_mid_4_36_imag;
  reg        [17:0]   data_mid_4_37_real;
  reg        [17:0]   data_mid_4_37_imag;
  reg        [17:0]   data_mid_4_38_real;
  reg        [17:0]   data_mid_4_38_imag;
  reg        [17:0]   data_mid_4_39_real;
  reg        [17:0]   data_mid_4_39_imag;
  reg        [17:0]   data_mid_4_40_real;
  reg        [17:0]   data_mid_4_40_imag;
  reg        [17:0]   data_mid_4_41_real;
  reg        [17:0]   data_mid_4_41_imag;
  reg        [17:0]   data_mid_4_42_real;
  reg        [17:0]   data_mid_4_42_imag;
  reg        [17:0]   data_mid_4_43_real;
  reg        [17:0]   data_mid_4_43_imag;
  reg        [17:0]   data_mid_4_44_real;
  reg        [17:0]   data_mid_4_44_imag;
  reg        [17:0]   data_mid_4_45_real;
  reg        [17:0]   data_mid_4_45_imag;
  reg        [17:0]   data_mid_4_46_real;
  reg        [17:0]   data_mid_4_46_imag;
  reg        [17:0]   data_mid_4_47_real;
  reg        [17:0]   data_mid_4_47_imag;
  reg        [17:0]   data_mid_4_48_real;
  reg        [17:0]   data_mid_4_48_imag;
  reg        [17:0]   data_mid_4_49_real;
  reg        [17:0]   data_mid_4_49_imag;
  reg        [17:0]   data_mid_4_50_real;
  reg        [17:0]   data_mid_4_50_imag;
  reg        [17:0]   data_mid_4_51_real;
  reg        [17:0]   data_mid_4_51_imag;
  reg        [17:0]   data_mid_4_52_real;
  reg        [17:0]   data_mid_4_52_imag;
  reg        [17:0]   data_mid_4_53_real;
  reg        [17:0]   data_mid_4_53_imag;
  reg        [17:0]   data_mid_4_54_real;
  reg        [17:0]   data_mid_4_54_imag;
  reg        [17:0]   data_mid_4_55_real;
  reg        [17:0]   data_mid_4_55_imag;
  reg        [17:0]   data_mid_4_56_real;
  reg        [17:0]   data_mid_4_56_imag;
  reg        [17:0]   data_mid_4_57_real;
  reg        [17:0]   data_mid_4_57_imag;
  reg        [17:0]   data_mid_4_58_real;
  reg        [17:0]   data_mid_4_58_imag;
  reg        [17:0]   data_mid_4_59_real;
  reg        [17:0]   data_mid_4_59_imag;
  reg        [17:0]   data_mid_4_60_real;
  reg        [17:0]   data_mid_4_60_imag;
  reg        [17:0]   data_mid_4_61_real;
  reg        [17:0]   data_mid_4_61_imag;
  reg        [17:0]   data_mid_4_62_real;
  reg        [17:0]   data_mid_4_62_imag;
  reg        [17:0]   data_mid_4_63_real;
  reg        [17:0]   data_mid_4_63_imag;
  reg        [17:0]   data_mid_5_0_real;
  reg        [17:0]   data_mid_5_0_imag;
  reg        [17:0]   data_mid_5_1_real;
  reg        [17:0]   data_mid_5_1_imag;
  reg        [17:0]   data_mid_5_2_real;
  reg        [17:0]   data_mid_5_2_imag;
  reg        [17:0]   data_mid_5_3_real;
  reg        [17:0]   data_mid_5_3_imag;
  reg        [17:0]   data_mid_5_4_real;
  reg        [17:0]   data_mid_5_4_imag;
  reg        [17:0]   data_mid_5_5_real;
  reg        [17:0]   data_mid_5_5_imag;
  reg        [17:0]   data_mid_5_6_real;
  reg        [17:0]   data_mid_5_6_imag;
  reg        [17:0]   data_mid_5_7_real;
  reg        [17:0]   data_mid_5_7_imag;
  reg        [17:0]   data_mid_5_8_real;
  reg        [17:0]   data_mid_5_8_imag;
  reg        [17:0]   data_mid_5_9_real;
  reg        [17:0]   data_mid_5_9_imag;
  reg        [17:0]   data_mid_5_10_real;
  reg        [17:0]   data_mid_5_10_imag;
  reg        [17:0]   data_mid_5_11_real;
  reg        [17:0]   data_mid_5_11_imag;
  reg        [17:0]   data_mid_5_12_real;
  reg        [17:0]   data_mid_5_12_imag;
  reg        [17:0]   data_mid_5_13_real;
  reg        [17:0]   data_mid_5_13_imag;
  reg        [17:0]   data_mid_5_14_real;
  reg        [17:0]   data_mid_5_14_imag;
  reg        [17:0]   data_mid_5_15_real;
  reg        [17:0]   data_mid_5_15_imag;
  reg        [17:0]   data_mid_5_16_real;
  reg        [17:0]   data_mid_5_16_imag;
  reg        [17:0]   data_mid_5_17_real;
  reg        [17:0]   data_mid_5_17_imag;
  reg        [17:0]   data_mid_5_18_real;
  reg        [17:0]   data_mid_5_18_imag;
  reg        [17:0]   data_mid_5_19_real;
  reg        [17:0]   data_mid_5_19_imag;
  reg        [17:0]   data_mid_5_20_real;
  reg        [17:0]   data_mid_5_20_imag;
  reg        [17:0]   data_mid_5_21_real;
  reg        [17:0]   data_mid_5_21_imag;
  reg        [17:0]   data_mid_5_22_real;
  reg        [17:0]   data_mid_5_22_imag;
  reg        [17:0]   data_mid_5_23_real;
  reg        [17:0]   data_mid_5_23_imag;
  reg        [17:0]   data_mid_5_24_real;
  reg        [17:0]   data_mid_5_24_imag;
  reg        [17:0]   data_mid_5_25_real;
  reg        [17:0]   data_mid_5_25_imag;
  reg        [17:0]   data_mid_5_26_real;
  reg        [17:0]   data_mid_5_26_imag;
  reg        [17:0]   data_mid_5_27_real;
  reg        [17:0]   data_mid_5_27_imag;
  reg        [17:0]   data_mid_5_28_real;
  reg        [17:0]   data_mid_5_28_imag;
  reg        [17:0]   data_mid_5_29_real;
  reg        [17:0]   data_mid_5_29_imag;
  reg        [17:0]   data_mid_5_30_real;
  reg        [17:0]   data_mid_5_30_imag;
  reg        [17:0]   data_mid_5_31_real;
  reg        [17:0]   data_mid_5_31_imag;
  reg        [17:0]   data_mid_5_32_real;
  reg        [17:0]   data_mid_5_32_imag;
  reg        [17:0]   data_mid_5_33_real;
  reg        [17:0]   data_mid_5_33_imag;
  reg        [17:0]   data_mid_5_34_real;
  reg        [17:0]   data_mid_5_34_imag;
  reg        [17:0]   data_mid_5_35_real;
  reg        [17:0]   data_mid_5_35_imag;
  reg        [17:0]   data_mid_5_36_real;
  reg        [17:0]   data_mid_5_36_imag;
  reg        [17:0]   data_mid_5_37_real;
  reg        [17:0]   data_mid_5_37_imag;
  reg        [17:0]   data_mid_5_38_real;
  reg        [17:0]   data_mid_5_38_imag;
  reg        [17:0]   data_mid_5_39_real;
  reg        [17:0]   data_mid_5_39_imag;
  reg        [17:0]   data_mid_5_40_real;
  reg        [17:0]   data_mid_5_40_imag;
  reg        [17:0]   data_mid_5_41_real;
  reg        [17:0]   data_mid_5_41_imag;
  reg        [17:0]   data_mid_5_42_real;
  reg        [17:0]   data_mid_5_42_imag;
  reg        [17:0]   data_mid_5_43_real;
  reg        [17:0]   data_mid_5_43_imag;
  reg        [17:0]   data_mid_5_44_real;
  reg        [17:0]   data_mid_5_44_imag;
  reg        [17:0]   data_mid_5_45_real;
  reg        [17:0]   data_mid_5_45_imag;
  reg        [17:0]   data_mid_5_46_real;
  reg        [17:0]   data_mid_5_46_imag;
  reg        [17:0]   data_mid_5_47_real;
  reg        [17:0]   data_mid_5_47_imag;
  reg        [17:0]   data_mid_5_48_real;
  reg        [17:0]   data_mid_5_48_imag;
  reg        [17:0]   data_mid_5_49_real;
  reg        [17:0]   data_mid_5_49_imag;
  reg        [17:0]   data_mid_5_50_real;
  reg        [17:0]   data_mid_5_50_imag;
  reg        [17:0]   data_mid_5_51_real;
  reg        [17:0]   data_mid_5_51_imag;
  reg        [17:0]   data_mid_5_52_real;
  reg        [17:0]   data_mid_5_52_imag;
  reg        [17:0]   data_mid_5_53_real;
  reg        [17:0]   data_mid_5_53_imag;
  reg        [17:0]   data_mid_5_54_real;
  reg        [17:0]   data_mid_5_54_imag;
  reg        [17:0]   data_mid_5_55_real;
  reg        [17:0]   data_mid_5_55_imag;
  reg        [17:0]   data_mid_5_56_real;
  reg        [17:0]   data_mid_5_56_imag;
  reg        [17:0]   data_mid_5_57_real;
  reg        [17:0]   data_mid_5_57_imag;
  reg        [17:0]   data_mid_5_58_real;
  reg        [17:0]   data_mid_5_58_imag;
  reg        [17:0]   data_mid_5_59_real;
  reg        [17:0]   data_mid_5_59_imag;
  reg        [17:0]   data_mid_5_60_real;
  reg        [17:0]   data_mid_5_60_imag;
  reg        [17:0]   data_mid_5_61_real;
  reg        [17:0]   data_mid_5_61_imag;
  reg        [17:0]   data_mid_5_62_real;
  reg        [17:0]   data_mid_5_62_imag;
  reg        [17:0]   data_mid_5_63_real;
  reg        [17:0]   data_mid_5_63_imag;
  reg        [17:0]   data_mid_6_0_real;
  reg        [17:0]   data_mid_6_0_imag;
  reg        [17:0]   data_mid_6_1_real;
  reg        [17:0]   data_mid_6_1_imag;
  reg        [17:0]   data_mid_6_2_real;
  reg        [17:0]   data_mid_6_2_imag;
  reg        [17:0]   data_mid_6_3_real;
  reg        [17:0]   data_mid_6_3_imag;
  reg        [17:0]   data_mid_6_4_real;
  reg        [17:0]   data_mid_6_4_imag;
  reg        [17:0]   data_mid_6_5_real;
  reg        [17:0]   data_mid_6_5_imag;
  reg        [17:0]   data_mid_6_6_real;
  reg        [17:0]   data_mid_6_6_imag;
  reg        [17:0]   data_mid_6_7_real;
  reg        [17:0]   data_mid_6_7_imag;
  reg        [17:0]   data_mid_6_8_real;
  reg        [17:0]   data_mid_6_8_imag;
  reg        [17:0]   data_mid_6_9_real;
  reg        [17:0]   data_mid_6_9_imag;
  reg        [17:0]   data_mid_6_10_real;
  reg        [17:0]   data_mid_6_10_imag;
  reg        [17:0]   data_mid_6_11_real;
  reg        [17:0]   data_mid_6_11_imag;
  reg        [17:0]   data_mid_6_12_real;
  reg        [17:0]   data_mid_6_12_imag;
  reg        [17:0]   data_mid_6_13_real;
  reg        [17:0]   data_mid_6_13_imag;
  reg        [17:0]   data_mid_6_14_real;
  reg        [17:0]   data_mid_6_14_imag;
  reg        [17:0]   data_mid_6_15_real;
  reg        [17:0]   data_mid_6_15_imag;
  reg        [17:0]   data_mid_6_16_real;
  reg        [17:0]   data_mid_6_16_imag;
  reg        [17:0]   data_mid_6_17_real;
  reg        [17:0]   data_mid_6_17_imag;
  reg        [17:0]   data_mid_6_18_real;
  reg        [17:0]   data_mid_6_18_imag;
  reg        [17:0]   data_mid_6_19_real;
  reg        [17:0]   data_mid_6_19_imag;
  reg        [17:0]   data_mid_6_20_real;
  reg        [17:0]   data_mid_6_20_imag;
  reg        [17:0]   data_mid_6_21_real;
  reg        [17:0]   data_mid_6_21_imag;
  reg        [17:0]   data_mid_6_22_real;
  reg        [17:0]   data_mid_6_22_imag;
  reg        [17:0]   data_mid_6_23_real;
  reg        [17:0]   data_mid_6_23_imag;
  reg        [17:0]   data_mid_6_24_real;
  reg        [17:0]   data_mid_6_24_imag;
  reg        [17:0]   data_mid_6_25_real;
  reg        [17:0]   data_mid_6_25_imag;
  reg        [17:0]   data_mid_6_26_real;
  reg        [17:0]   data_mid_6_26_imag;
  reg        [17:0]   data_mid_6_27_real;
  reg        [17:0]   data_mid_6_27_imag;
  reg        [17:0]   data_mid_6_28_real;
  reg        [17:0]   data_mid_6_28_imag;
  reg        [17:0]   data_mid_6_29_real;
  reg        [17:0]   data_mid_6_29_imag;
  reg        [17:0]   data_mid_6_30_real;
  reg        [17:0]   data_mid_6_30_imag;
  reg        [17:0]   data_mid_6_31_real;
  reg        [17:0]   data_mid_6_31_imag;
  reg        [17:0]   data_mid_6_32_real;
  reg        [17:0]   data_mid_6_32_imag;
  reg        [17:0]   data_mid_6_33_real;
  reg        [17:0]   data_mid_6_33_imag;
  reg        [17:0]   data_mid_6_34_real;
  reg        [17:0]   data_mid_6_34_imag;
  reg        [17:0]   data_mid_6_35_real;
  reg        [17:0]   data_mid_6_35_imag;
  reg        [17:0]   data_mid_6_36_real;
  reg        [17:0]   data_mid_6_36_imag;
  reg        [17:0]   data_mid_6_37_real;
  reg        [17:0]   data_mid_6_37_imag;
  reg        [17:0]   data_mid_6_38_real;
  reg        [17:0]   data_mid_6_38_imag;
  reg        [17:0]   data_mid_6_39_real;
  reg        [17:0]   data_mid_6_39_imag;
  reg        [17:0]   data_mid_6_40_real;
  reg        [17:0]   data_mid_6_40_imag;
  reg        [17:0]   data_mid_6_41_real;
  reg        [17:0]   data_mid_6_41_imag;
  reg        [17:0]   data_mid_6_42_real;
  reg        [17:0]   data_mid_6_42_imag;
  reg        [17:0]   data_mid_6_43_real;
  reg        [17:0]   data_mid_6_43_imag;
  reg        [17:0]   data_mid_6_44_real;
  reg        [17:0]   data_mid_6_44_imag;
  reg        [17:0]   data_mid_6_45_real;
  reg        [17:0]   data_mid_6_45_imag;
  reg        [17:0]   data_mid_6_46_real;
  reg        [17:0]   data_mid_6_46_imag;
  reg        [17:0]   data_mid_6_47_real;
  reg        [17:0]   data_mid_6_47_imag;
  reg        [17:0]   data_mid_6_48_real;
  reg        [17:0]   data_mid_6_48_imag;
  reg        [17:0]   data_mid_6_49_real;
  reg        [17:0]   data_mid_6_49_imag;
  reg        [17:0]   data_mid_6_50_real;
  reg        [17:0]   data_mid_6_50_imag;
  reg        [17:0]   data_mid_6_51_real;
  reg        [17:0]   data_mid_6_51_imag;
  reg        [17:0]   data_mid_6_52_real;
  reg        [17:0]   data_mid_6_52_imag;
  reg        [17:0]   data_mid_6_53_real;
  reg        [17:0]   data_mid_6_53_imag;
  reg        [17:0]   data_mid_6_54_real;
  reg        [17:0]   data_mid_6_54_imag;
  reg        [17:0]   data_mid_6_55_real;
  reg        [17:0]   data_mid_6_55_imag;
  reg        [17:0]   data_mid_6_56_real;
  reg        [17:0]   data_mid_6_56_imag;
  reg        [17:0]   data_mid_6_57_real;
  reg        [17:0]   data_mid_6_57_imag;
  reg        [17:0]   data_mid_6_58_real;
  reg        [17:0]   data_mid_6_58_imag;
  reg        [17:0]   data_mid_6_59_real;
  reg        [17:0]   data_mid_6_59_imag;
  reg        [17:0]   data_mid_6_60_real;
  reg        [17:0]   data_mid_6_60_imag;
  reg        [17:0]   data_mid_6_61_real;
  reg        [17:0]   data_mid_6_61_imag;
  reg        [17:0]   data_mid_6_62_real;
  reg        [17:0]   data_mid_6_62_imag;
  reg        [17:0]   data_mid_6_63_real;
  reg        [17:0]   data_mid_6_63_imag;
  wire       [35:0]   _zz_1;
  wire       [35:0]   _zz_2;
  wire       [35:0]   _zz_3;
  wire       [0:0]    _zz_4;
  wire       [0:0]    _zz_5;
  wire       [35:0]   _zz_6;
  wire       [35:0]   _zz_7;
  wire       [35:0]   _zz_8;
  wire       [0:0]    _zz_9;
  wire       [0:0]    _zz_10;
  wire       [35:0]   _zz_11;
  wire       [35:0]   _zz_12;
  wire       [35:0]   _zz_13;
  wire       [0:0]    _zz_14;
  wire       [0:0]    _zz_15;
  wire       [35:0]   _zz_16;
  wire       [35:0]   _zz_17;
  wire       [35:0]   _zz_18;
  wire       [0:0]    _zz_19;
  wire       [0:0]    _zz_20;
  wire       [35:0]   _zz_21;
  wire       [35:0]   _zz_22;
  wire       [35:0]   _zz_23;
  wire       [0:0]    _zz_24;
  wire       [0:0]    _zz_25;
  wire       [35:0]   _zz_26;
  wire       [35:0]   _zz_27;
  wire       [35:0]   _zz_28;
  wire       [0:0]    _zz_29;
  wire       [0:0]    _zz_30;
  wire       [35:0]   _zz_31;
  wire       [35:0]   _zz_32;
  wire       [35:0]   _zz_33;
  wire       [0:0]    _zz_34;
  wire       [0:0]    _zz_35;
  wire       [35:0]   _zz_36;
  wire       [35:0]   _zz_37;
  wire       [35:0]   _zz_38;
  wire       [0:0]    _zz_39;
  wire       [0:0]    _zz_40;
  wire       [35:0]   _zz_41;
  wire       [35:0]   _zz_42;
  wire       [35:0]   _zz_43;
  wire       [0:0]    _zz_44;
  wire       [0:0]    _zz_45;
  wire       [35:0]   _zz_46;
  wire       [35:0]   _zz_47;
  wire       [35:0]   _zz_48;
  wire       [0:0]    _zz_49;
  wire       [0:0]    _zz_50;
  wire       [35:0]   _zz_51;
  wire       [35:0]   _zz_52;
  wire       [35:0]   _zz_53;
  wire       [0:0]    _zz_54;
  wire       [0:0]    _zz_55;
  wire       [35:0]   _zz_56;
  wire       [35:0]   _zz_57;
  wire       [35:0]   _zz_58;
  wire       [0:0]    _zz_59;
  wire       [0:0]    _zz_60;
  wire       [35:0]   _zz_61;
  wire       [35:0]   _zz_62;
  wire       [35:0]   _zz_63;
  wire       [0:0]    _zz_64;
  wire       [0:0]    _zz_65;
  wire       [35:0]   _zz_66;
  wire       [35:0]   _zz_67;
  wire       [35:0]   _zz_68;
  wire       [0:0]    _zz_69;
  wire       [0:0]    _zz_70;
  wire       [35:0]   _zz_71;
  wire       [35:0]   _zz_72;
  wire       [35:0]   _zz_73;
  wire       [0:0]    _zz_74;
  wire       [0:0]    _zz_75;
  wire       [35:0]   _zz_76;
  wire       [35:0]   _zz_77;
  wire       [35:0]   _zz_78;
  wire       [0:0]    _zz_79;
  wire       [0:0]    _zz_80;
  wire       [35:0]   _zz_81;
  wire       [35:0]   _zz_82;
  wire       [35:0]   _zz_83;
  wire       [0:0]    _zz_84;
  wire       [0:0]    _zz_85;
  wire       [35:0]   _zz_86;
  wire       [35:0]   _zz_87;
  wire       [35:0]   _zz_88;
  wire       [0:0]    _zz_89;
  wire       [0:0]    _zz_90;
  wire       [35:0]   _zz_91;
  wire       [35:0]   _zz_92;
  wire       [35:0]   _zz_93;
  wire       [0:0]    _zz_94;
  wire       [0:0]    _zz_95;
  wire       [35:0]   _zz_96;
  wire       [35:0]   _zz_97;
  wire       [35:0]   _zz_98;
  wire       [0:0]    _zz_99;
  wire       [0:0]    _zz_100;
  wire       [35:0]   _zz_101;
  wire       [35:0]   _zz_102;
  wire       [35:0]   _zz_103;
  wire       [0:0]    _zz_104;
  wire       [0:0]    _zz_105;
  wire       [35:0]   _zz_106;
  wire       [35:0]   _zz_107;
  wire       [35:0]   _zz_108;
  wire       [0:0]    _zz_109;
  wire       [0:0]    _zz_110;
  wire       [35:0]   _zz_111;
  wire       [35:0]   _zz_112;
  wire       [35:0]   _zz_113;
  wire       [0:0]    _zz_114;
  wire       [0:0]    _zz_115;
  wire       [35:0]   _zz_116;
  wire       [35:0]   _zz_117;
  wire       [35:0]   _zz_118;
  wire       [0:0]    _zz_119;
  wire       [0:0]    _zz_120;
  wire       [35:0]   _zz_121;
  wire       [35:0]   _zz_122;
  wire       [35:0]   _zz_123;
  wire       [0:0]    _zz_124;
  wire       [0:0]    _zz_125;
  wire       [35:0]   _zz_126;
  wire       [35:0]   _zz_127;
  wire       [35:0]   _zz_128;
  wire       [0:0]    _zz_129;
  wire       [0:0]    _zz_130;
  wire       [35:0]   _zz_131;
  wire       [35:0]   _zz_132;
  wire       [35:0]   _zz_133;
  wire       [0:0]    _zz_134;
  wire       [0:0]    _zz_135;
  wire       [35:0]   _zz_136;
  wire       [35:0]   _zz_137;
  wire       [35:0]   _zz_138;
  wire       [0:0]    _zz_139;
  wire       [0:0]    _zz_140;
  wire       [35:0]   _zz_141;
  wire       [35:0]   _zz_142;
  wire       [35:0]   _zz_143;
  wire       [0:0]    _zz_144;
  wire       [0:0]    _zz_145;
  wire       [35:0]   _zz_146;
  wire       [35:0]   _zz_147;
  wire       [35:0]   _zz_148;
  wire       [0:0]    _zz_149;
  wire       [0:0]    _zz_150;
  wire       [35:0]   _zz_151;
  wire       [35:0]   _zz_152;
  wire       [35:0]   _zz_153;
  wire       [0:0]    _zz_154;
  wire       [0:0]    _zz_155;
  wire       [35:0]   _zz_156;
  wire       [35:0]   _zz_157;
  wire       [35:0]   _zz_158;
  wire       [0:0]    _zz_159;
  wire       [0:0]    _zz_160;
  wire       [35:0]   _zz_161;
  wire       [35:0]   _zz_162;
  wire       [35:0]   _zz_163;
  wire       [0:0]    _zz_164;
  wire       [0:0]    _zz_165;
  wire       [35:0]   _zz_166;
  wire       [35:0]   _zz_167;
  wire       [35:0]   _zz_168;
  wire       [0:0]    _zz_169;
  wire       [0:0]    _zz_170;
  wire       [35:0]   _zz_171;
  wire       [35:0]   _zz_172;
  wire       [35:0]   _zz_173;
  wire       [0:0]    _zz_174;
  wire       [0:0]    _zz_175;
  wire       [35:0]   _zz_176;
  wire       [35:0]   _zz_177;
  wire       [35:0]   _zz_178;
  wire       [0:0]    _zz_179;
  wire       [0:0]    _zz_180;
  wire       [35:0]   _zz_181;
  wire       [35:0]   _zz_182;
  wire       [35:0]   _zz_183;
  wire       [0:0]    _zz_184;
  wire       [0:0]    _zz_185;
  wire       [35:0]   _zz_186;
  wire       [35:0]   _zz_187;
  wire       [35:0]   _zz_188;
  wire       [0:0]    _zz_189;
  wire       [0:0]    _zz_190;
  wire       [35:0]   _zz_191;
  wire       [35:0]   _zz_192;
  wire       [35:0]   _zz_193;
  wire       [0:0]    _zz_194;
  wire       [0:0]    _zz_195;
  wire       [35:0]   _zz_196;
  wire       [35:0]   _zz_197;
  wire       [35:0]   _zz_198;
  wire       [0:0]    _zz_199;
  wire       [0:0]    _zz_200;
  wire       [35:0]   _zz_201;
  wire       [35:0]   _zz_202;
  wire       [35:0]   _zz_203;
  wire       [0:0]    _zz_204;
  wire       [0:0]    _zz_205;
  wire       [35:0]   _zz_206;
  wire       [35:0]   _zz_207;
  wire       [35:0]   _zz_208;
  wire       [0:0]    _zz_209;
  wire       [0:0]    _zz_210;
  wire       [35:0]   _zz_211;
  wire       [35:0]   _zz_212;
  wire       [35:0]   _zz_213;
  wire       [0:0]    _zz_214;
  wire       [0:0]    _zz_215;
  wire       [35:0]   _zz_216;
  wire       [35:0]   _zz_217;
  wire       [35:0]   _zz_218;
  wire       [0:0]    _zz_219;
  wire       [0:0]    _zz_220;
  wire       [35:0]   _zz_221;
  wire       [35:0]   _zz_222;
  wire       [35:0]   _zz_223;
  wire       [0:0]    _zz_224;
  wire       [0:0]    _zz_225;
  wire       [35:0]   _zz_226;
  wire       [35:0]   _zz_227;
  wire       [35:0]   _zz_228;
  wire       [0:0]    _zz_229;
  wire       [0:0]    _zz_230;
  wire       [35:0]   _zz_231;
  wire       [35:0]   _zz_232;
  wire       [35:0]   _zz_233;
  wire       [0:0]    _zz_234;
  wire       [0:0]    _zz_235;
  wire       [35:0]   _zz_236;
  wire       [35:0]   _zz_237;
  wire       [35:0]   _zz_238;
  wire       [0:0]    _zz_239;
  wire       [0:0]    _zz_240;
  wire       [35:0]   _zz_241;
  wire       [35:0]   _zz_242;
  wire       [35:0]   _zz_243;
  wire       [0:0]    _zz_244;
  wire       [0:0]    _zz_245;
  wire       [35:0]   _zz_246;
  wire       [35:0]   _zz_247;
  wire       [35:0]   _zz_248;
  wire       [0:0]    _zz_249;
  wire       [0:0]    _zz_250;
  wire       [35:0]   _zz_251;
  wire       [35:0]   _zz_252;
  wire       [35:0]   _zz_253;
  wire       [0:0]    _zz_254;
  wire       [0:0]    _zz_255;
  wire       [35:0]   _zz_256;
  wire       [35:0]   _zz_257;
  wire       [35:0]   _zz_258;
  wire       [0:0]    _zz_259;
  wire       [0:0]    _zz_260;
  wire       [35:0]   _zz_261;
  wire       [35:0]   _zz_262;
  wire       [35:0]   _zz_263;
  wire       [0:0]    _zz_264;
  wire       [0:0]    _zz_265;
  wire       [35:0]   _zz_266;
  wire       [35:0]   _zz_267;
  wire       [35:0]   _zz_268;
  wire       [0:0]    _zz_269;
  wire       [0:0]    _zz_270;
  wire       [35:0]   _zz_271;
  wire       [35:0]   _zz_272;
  wire       [35:0]   _zz_273;
  wire       [0:0]    _zz_274;
  wire       [0:0]    _zz_275;
  wire       [35:0]   _zz_276;
  wire       [35:0]   _zz_277;
  wire       [35:0]   _zz_278;
  wire       [0:0]    _zz_279;
  wire       [0:0]    _zz_280;
  wire       [35:0]   _zz_281;
  wire       [35:0]   _zz_282;
  wire       [35:0]   _zz_283;
  wire       [0:0]    _zz_284;
  wire       [0:0]    _zz_285;
  wire       [35:0]   _zz_286;
  wire       [35:0]   _zz_287;
  wire       [35:0]   _zz_288;
  wire       [0:0]    _zz_289;
  wire       [0:0]    _zz_290;
  wire       [35:0]   _zz_291;
  wire       [35:0]   _zz_292;
  wire       [35:0]   _zz_293;
  wire       [0:0]    _zz_294;
  wire       [0:0]    _zz_295;
  wire       [35:0]   _zz_296;
  wire       [35:0]   _zz_297;
  wire       [35:0]   _zz_298;
  wire       [0:0]    _zz_299;
  wire       [0:0]    _zz_300;
  wire       [35:0]   _zz_301;
  wire       [35:0]   _zz_302;
  wire       [35:0]   _zz_303;
  wire       [0:0]    _zz_304;
  wire       [0:0]    _zz_305;
  wire       [35:0]   _zz_306;
  wire       [35:0]   _zz_307;
  wire       [35:0]   _zz_308;
  wire       [0:0]    _zz_309;
  wire       [0:0]    _zz_310;
  wire       [35:0]   _zz_311;
  wire       [35:0]   _zz_312;
  wire       [35:0]   _zz_313;
  wire       [0:0]    _zz_314;
  wire       [0:0]    _zz_315;
  wire       [35:0]   _zz_316;
  wire       [35:0]   _zz_317;
  wire       [35:0]   _zz_318;
  wire       [0:0]    _zz_319;
  wire       [0:0]    _zz_320;
  wire       [35:0]   _zz_321;
  wire       [35:0]   _zz_322;
  wire       [35:0]   _zz_323;
  wire       [0:0]    _zz_324;
  wire       [0:0]    _zz_325;
  wire       [35:0]   _zz_326;
  wire       [35:0]   _zz_327;
  wire       [35:0]   _zz_328;
  wire       [0:0]    _zz_329;
  wire       [0:0]    _zz_330;
  wire       [35:0]   _zz_331;
  wire       [35:0]   _zz_332;
  wire       [35:0]   _zz_333;
  wire       [0:0]    _zz_334;
  wire       [0:0]    _zz_335;
  wire       [35:0]   _zz_336;
  wire       [35:0]   _zz_337;
  wire       [35:0]   _zz_338;
  wire       [0:0]    _zz_339;
  wire       [0:0]    _zz_340;
  wire       [35:0]   _zz_341;
  wire       [35:0]   _zz_342;
  wire       [35:0]   _zz_343;
  wire       [0:0]    _zz_344;
  wire       [0:0]    _zz_345;
  wire       [35:0]   _zz_346;
  wire       [35:0]   _zz_347;
  wire       [35:0]   _zz_348;
  wire       [0:0]    _zz_349;
  wire       [0:0]    _zz_350;
  wire       [35:0]   _zz_351;
  wire       [35:0]   _zz_352;
  wire       [35:0]   _zz_353;
  wire       [0:0]    _zz_354;
  wire       [0:0]    _zz_355;
  wire       [35:0]   _zz_356;
  wire       [35:0]   _zz_357;
  wire       [35:0]   _zz_358;
  wire       [0:0]    _zz_359;
  wire       [0:0]    _zz_360;
  wire       [35:0]   _zz_361;
  wire       [35:0]   _zz_362;
  wire       [35:0]   _zz_363;
  wire       [0:0]    _zz_364;
  wire       [0:0]    _zz_365;
  wire       [35:0]   _zz_366;
  wire       [35:0]   _zz_367;
  wire       [35:0]   _zz_368;
  wire       [0:0]    _zz_369;
  wire       [0:0]    _zz_370;
  wire       [35:0]   _zz_371;
  wire       [35:0]   _zz_372;
  wire       [35:0]   _zz_373;
  wire       [0:0]    _zz_374;
  wire       [0:0]    _zz_375;
  wire       [35:0]   _zz_376;
  wire       [35:0]   _zz_377;
  wire       [35:0]   _zz_378;
  wire       [0:0]    _zz_379;
  wire       [0:0]    _zz_380;
  wire       [35:0]   _zz_381;
  wire       [35:0]   _zz_382;
  wire       [35:0]   _zz_383;
  wire       [0:0]    _zz_384;
  wire       [0:0]    _zz_385;
  wire       [35:0]   _zz_386;
  wire       [35:0]   _zz_387;
  wire       [35:0]   _zz_388;
  wire       [0:0]    _zz_389;
  wire       [0:0]    _zz_390;
  wire       [35:0]   _zz_391;
  wire       [35:0]   _zz_392;
  wire       [35:0]   _zz_393;
  wire       [0:0]    _zz_394;
  wire       [0:0]    _zz_395;
  wire       [35:0]   _zz_396;
  wire       [35:0]   _zz_397;
  wire       [35:0]   _zz_398;
  wire       [0:0]    _zz_399;
  wire       [0:0]    _zz_400;
  wire       [35:0]   _zz_401;
  wire       [35:0]   _zz_402;
  wire       [35:0]   _zz_403;
  wire       [0:0]    _zz_404;
  wire       [0:0]    _zz_405;
  wire       [35:0]   _zz_406;
  wire       [35:0]   _zz_407;
  wire       [35:0]   _zz_408;
  wire       [0:0]    _zz_409;
  wire       [0:0]    _zz_410;
  wire       [35:0]   _zz_411;
  wire       [35:0]   _zz_412;
  wire       [35:0]   _zz_413;
  wire       [0:0]    _zz_414;
  wire       [0:0]    _zz_415;
  wire       [35:0]   _zz_416;
  wire       [35:0]   _zz_417;
  wire       [35:0]   _zz_418;
  wire       [0:0]    _zz_419;
  wire       [0:0]    _zz_420;
  wire       [35:0]   _zz_421;
  wire       [35:0]   _zz_422;
  wire       [35:0]   _zz_423;
  wire       [0:0]    _zz_424;
  wire       [0:0]    _zz_425;
  wire       [35:0]   _zz_426;
  wire       [35:0]   _zz_427;
  wire       [35:0]   _zz_428;
  wire       [0:0]    _zz_429;
  wire       [0:0]    _zz_430;
  wire       [35:0]   _zz_431;
  wire       [35:0]   _zz_432;
  wire       [35:0]   _zz_433;
  wire       [0:0]    _zz_434;
  wire       [0:0]    _zz_435;
  wire       [35:0]   _zz_436;
  wire       [35:0]   _zz_437;
  wire       [35:0]   _zz_438;
  wire       [0:0]    _zz_439;
  wire       [0:0]    _zz_440;
  wire       [35:0]   _zz_441;
  wire       [35:0]   _zz_442;
  wire       [35:0]   _zz_443;
  wire       [0:0]    _zz_444;
  wire       [0:0]    _zz_445;
  wire       [35:0]   _zz_446;
  wire       [35:0]   _zz_447;
  wire       [35:0]   _zz_448;
  wire       [0:0]    _zz_449;
  wire       [0:0]    _zz_450;
  wire       [35:0]   _zz_451;
  wire       [35:0]   _zz_452;
  wire       [35:0]   _zz_453;
  wire       [0:0]    _zz_454;
  wire       [0:0]    _zz_455;
  wire       [35:0]   _zz_456;
  wire       [35:0]   _zz_457;
  wire       [35:0]   _zz_458;
  wire       [0:0]    _zz_459;
  wire       [0:0]    _zz_460;
  wire       [35:0]   _zz_461;
  wire       [35:0]   _zz_462;
  wire       [35:0]   _zz_463;
  wire       [0:0]    _zz_464;
  wire       [0:0]    _zz_465;
  wire       [35:0]   _zz_466;
  wire       [35:0]   _zz_467;
  wire       [35:0]   _zz_468;
  wire       [0:0]    _zz_469;
  wire       [0:0]    _zz_470;
  wire       [35:0]   _zz_471;
  wire       [35:0]   _zz_472;
  wire       [35:0]   _zz_473;
  wire       [0:0]    _zz_474;
  wire       [0:0]    _zz_475;
  wire       [35:0]   _zz_476;
  wire       [35:0]   _zz_477;
  wire       [35:0]   _zz_478;
  wire       [0:0]    _zz_479;
  wire       [0:0]    _zz_480;
  wire       [35:0]   _zz_481;
  wire       [35:0]   _zz_482;
  wire       [35:0]   _zz_483;
  wire       [0:0]    _zz_484;
  wire       [0:0]    _zz_485;
  wire       [35:0]   _zz_486;
  wire       [35:0]   _zz_487;
  wire       [35:0]   _zz_488;
  wire       [0:0]    _zz_489;
  wire       [0:0]    _zz_490;
  wire       [35:0]   _zz_491;
  wire       [35:0]   _zz_492;
  wire       [35:0]   _zz_493;
  wire       [0:0]    _zz_494;
  wire       [0:0]    _zz_495;
  wire       [35:0]   _zz_496;
  wire       [35:0]   _zz_497;
  wire       [35:0]   _zz_498;
  wire       [0:0]    _zz_499;
  wire       [0:0]    _zz_500;
  wire       [35:0]   _zz_501;
  wire       [35:0]   _zz_502;
  wire       [35:0]   _zz_503;
  wire       [0:0]    _zz_504;
  wire       [0:0]    _zz_505;
  wire       [35:0]   _zz_506;
  wire       [35:0]   _zz_507;
  wire       [35:0]   _zz_508;
  wire       [0:0]    _zz_509;
  wire       [0:0]    _zz_510;
  wire       [35:0]   _zz_511;
  wire       [35:0]   _zz_512;
  wire       [35:0]   _zz_513;
  wire       [0:0]    _zz_514;
  wire       [0:0]    _zz_515;
  wire       [35:0]   _zz_516;
  wire       [35:0]   _zz_517;
  wire       [35:0]   _zz_518;
  wire       [0:0]    _zz_519;
  wire       [0:0]    _zz_520;
  wire       [35:0]   _zz_521;
  wire       [35:0]   _zz_522;
  wire       [35:0]   _zz_523;
  wire       [0:0]    _zz_524;
  wire       [0:0]    _zz_525;
  wire       [35:0]   _zz_526;
  wire       [35:0]   _zz_527;
  wire       [35:0]   _zz_528;
  wire       [0:0]    _zz_529;
  wire       [0:0]    _zz_530;
  wire       [35:0]   _zz_531;
  wire       [35:0]   _zz_532;
  wire       [35:0]   _zz_533;
  wire       [0:0]    _zz_534;
  wire       [0:0]    _zz_535;
  wire       [35:0]   _zz_536;
  wire       [35:0]   _zz_537;
  wire       [35:0]   _zz_538;
  wire       [0:0]    _zz_539;
  wire       [0:0]    _zz_540;
  wire       [35:0]   _zz_541;
  wire       [35:0]   _zz_542;
  wire       [35:0]   _zz_543;
  wire       [0:0]    _zz_544;
  wire       [0:0]    _zz_545;
  wire       [35:0]   _zz_546;
  wire       [35:0]   _zz_547;
  wire       [35:0]   _zz_548;
  wire       [0:0]    _zz_549;
  wire       [0:0]    _zz_550;
  wire       [35:0]   _zz_551;
  wire       [35:0]   _zz_552;
  wire       [35:0]   _zz_553;
  wire       [0:0]    _zz_554;
  wire       [0:0]    _zz_555;
  wire       [35:0]   _zz_556;
  wire       [35:0]   _zz_557;
  wire       [35:0]   _zz_558;
  wire       [0:0]    _zz_559;
  wire       [0:0]    _zz_560;
  wire       [35:0]   _zz_561;
  wire       [35:0]   _zz_562;
  wire       [35:0]   _zz_563;
  wire       [0:0]    _zz_564;
  wire       [0:0]    _zz_565;
  wire       [35:0]   _zz_566;
  wire       [35:0]   _zz_567;
  wire       [35:0]   _zz_568;
  wire       [0:0]    _zz_569;
  wire       [0:0]    _zz_570;
  wire       [35:0]   _zz_571;
  wire       [35:0]   _zz_572;
  wire       [35:0]   _zz_573;
  wire       [0:0]    _zz_574;
  wire       [0:0]    _zz_575;
  wire       [35:0]   _zz_576;
  wire       [35:0]   _zz_577;
  wire       [35:0]   _zz_578;
  wire       [0:0]    _zz_579;
  wire       [0:0]    _zz_580;
  wire       [35:0]   _zz_581;
  wire       [35:0]   _zz_582;
  wire       [35:0]   _zz_583;
  wire       [0:0]    _zz_584;
  wire       [0:0]    _zz_585;
  wire       [35:0]   _zz_586;
  wire       [35:0]   _zz_587;
  wire       [35:0]   _zz_588;
  wire       [0:0]    _zz_589;
  wire       [0:0]    _zz_590;
  wire       [35:0]   _zz_591;
  wire       [35:0]   _zz_592;
  wire       [35:0]   _zz_593;
  wire       [0:0]    _zz_594;
  wire       [0:0]    _zz_595;
  wire       [35:0]   _zz_596;
  wire       [35:0]   _zz_597;
  wire       [35:0]   _zz_598;
  wire       [0:0]    _zz_599;
  wire       [0:0]    _zz_600;
  wire       [35:0]   _zz_601;
  wire       [35:0]   _zz_602;
  wire       [35:0]   _zz_603;
  wire       [0:0]    _zz_604;
  wire       [0:0]    _zz_605;
  wire       [35:0]   _zz_606;
  wire       [35:0]   _zz_607;
  wire       [35:0]   _zz_608;
  wire       [0:0]    _zz_609;
  wire       [0:0]    _zz_610;
  wire       [35:0]   _zz_611;
  wire       [35:0]   _zz_612;
  wire       [35:0]   _zz_613;
  wire       [0:0]    _zz_614;
  wire       [0:0]    _zz_615;
  wire       [35:0]   _zz_616;
  wire       [35:0]   _zz_617;
  wire       [35:0]   _zz_618;
  wire       [0:0]    _zz_619;
  wire       [0:0]    _zz_620;
  wire       [35:0]   _zz_621;
  wire       [35:0]   _zz_622;
  wire       [35:0]   _zz_623;
  wire       [0:0]    _zz_624;
  wire       [0:0]    _zz_625;
  wire       [35:0]   _zz_626;
  wire       [35:0]   _zz_627;
  wire       [35:0]   _zz_628;
  wire       [0:0]    _zz_629;
  wire       [0:0]    _zz_630;
  wire       [35:0]   _zz_631;
  wire       [35:0]   _zz_632;
  wire       [35:0]   _zz_633;
  wire       [0:0]    _zz_634;
  wire       [0:0]    _zz_635;
  wire       [35:0]   _zz_636;
  wire       [35:0]   _zz_637;
  wire       [35:0]   _zz_638;
  wire       [0:0]    _zz_639;
  wire       [0:0]    _zz_640;
  wire       [35:0]   _zz_641;
  wire       [35:0]   _zz_642;
  wire       [35:0]   _zz_643;
  wire       [0:0]    _zz_644;
  wire       [0:0]    _zz_645;
  wire       [35:0]   _zz_646;
  wire       [35:0]   _zz_647;
  wire       [35:0]   _zz_648;
  wire       [0:0]    _zz_649;
  wire       [0:0]    _zz_650;
  wire       [35:0]   _zz_651;
  wire       [35:0]   _zz_652;
  wire       [35:0]   _zz_653;
  wire       [0:0]    _zz_654;
  wire       [0:0]    _zz_655;
  wire       [35:0]   _zz_656;
  wire       [35:0]   _zz_657;
  wire       [35:0]   _zz_658;
  wire       [0:0]    _zz_659;
  wire       [0:0]    _zz_660;
  wire       [35:0]   _zz_661;
  wire       [35:0]   _zz_662;
  wire       [35:0]   _zz_663;
  wire       [0:0]    _zz_664;
  wire       [0:0]    _zz_665;
  wire       [35:0]   _zz_666;
  wire       [35:0]   _zz_667;
  wire       [35:0]   _zz_668;
  wire       [0:0]    _zz_669;
  wire       [0:0]    _zz_670;
  wire       [35:0]   _zz_671;
  wire       [35:0]   _zz_672;
  wire       [35:0]   _zz_673;
  wire       [0:0]    _zz_674;
  wire       [0:0]    _zz_675;
  wire       [35:0]   _zz_676;
  wire       [35:0]   _zz_677;
  wire       [35:0]   _zz_678;
  wire       [0:0]    _zz_679;
  wire       [0:0]    _zz_680;
  wire       [35:0]   _zz_681;
  wire       [35:0]   _zz_682;
  wire       [35:0]   _zz_683;
  wire       [0:0]    _zz_684;
  wire       [0:0]    _zz_685;
  wire       [35:0]   _zz_686;
  wire       [35:0]   _zz_687;
  wire       [35:0]   _zz_688;
  wire       [0:0]    _zz_689;
  wire       [0:0]    _zz_690;
  wire       [35:0]   _zz_691;
  wire       [35:0]   _zz_692;
  wire       [35:0]   _zz_693;
  wire       [0:0]    _zz_694;
  wire       [0:0]    _zz_695;
  wire       [35:0]   _zz_696;
  wire       [35:0]   _zz_697;
  wire       [35:0]   _zz_698;
  wire       [0:0]    _zz_699;
  wire       [0:0]    _zz_700;
  wire       [35:0]   _zz_701;
  wire       [35:0]   _zz_702;
  wire       [35:0]   _zz_703;
  wire       [0:0]    _zz_704;
  wire       [0:0]    _zz_705;
  wire       [35:0]   _zz_706;
  wire       [35:0]   _zz_707;
  wire       [35:0]   _zz_708;
  wire       [0:0]    _zz_709;
  wire       [0:0]    _zz_710;
  wire       [35:0]   _zz_711;
  wire       [35:0]   _zz_712;
  wire       [35:0]   _zz_713;
  wire       [0:0]    _zz_714;
  wire       [0:0]    _zz_715;
  wire       [35:0]   _zz_716;
  wire       [35:0]   _zz_717;
  wire       [35:0]   _zz_718;
  wire       [0:0]    _zz_719;
  wire       [0:0]    _zz_720;
  wire       [35:0]   _zz_721;
  wire       [35:0]   _zz_722;
  wire       [35:0]   _zz_723;
  wire       [0:0]    _zz_724;
  wire       [0:0]    _zz_725;
  wire       [35:0]   _zz_726;
  wire       [35:0]   _zz_727;
  wire       [35:0]   _zz_728;
  wire       [0:0]    _zz_729;
  wire       [0:0]    _zz_730;
  wire       [35:0]   _zz_731;
  wire       [35:0]   _zz_732;
  wire       [35:0]   _zz_733;
  wire       [0:0]    _zz_734;
  wire       [0:0]    _zz_735;
  wire       [35:0]   _zz_736;
  wire       [35:0]   _zz_737;
  wire       [35:0]   _zz_738;
  wire       [0:0]    _zz_739;
  wire       [0:0]    _zz_740;
  wire       [35:0]   _zz_741;
  wire       [35:0]   _zz_742;
  wire       [35:0]   _zz_743;
  wire       [0:0]    _zz_744;
  wire       [0:0]    _zz_745;
  wire       [35:0]   _zz_746;
  wire       [35:0]   _zz_747;
  wire       [35:0]   _zz_748;
  wire       [0:0]    _zz_749;
  wire       [0:0]    _zz_750;
  wire       [35:0]   _zz_751;
  wire       [35:0]   _zz_752;
  wire       [35:0]   _zz_753;
  wire       [0:0]    _zz_754;
  wire       [0:0]    _zz_755;
  wire       [35:0]   _zz_756;
  wire       [35:0]   _zz_757;
  wire       [35:0]   _zz_758;
  wire       [0:0]    _zz_759;
  wire       [0:0]    _zz_760;
  wire       [35:0]   _zz_761;
  wire       [35:0]   _zz_762;
  wire       [35:0]   _zz_763;
  wire       [0:0]    _zz_764;
  wire       [0:0]    _zz_765;
  wire       [35:0]   _zz_766;
  wire       [35:0]   _zz_767;
  wire       [35:0]   _zz_768;
  wire       [0:0]    _zz_769;
  wire       [0:0]    _zz_770;
  wire       [35:0]   _zz_771;
  wire       [35:0]   _zz_772;
  wire       [35:0]   _zz_773;
  wire       [0:0]    _zz_774;
  wire       [0:0]    _zz_775;
  wire       [35:0]   _zz_776;
  wire       [35:0]   _zz_777;
  wire       [35:0]   _zz_778;
  wire       [0:0]    _zz_779;
  wire       [0:0]    _zz_780;
  wire       [35:0]   _zz_781;
  wire       [35:0]   _zz_782;
  wire       [35:0]   _zz_783;
  wire       [0:0]    _zz_784;
  wire       [0:0]    _zz_785;
  wire       [35:0]   _zz_786;
  wire       [35:0]   _zz_787;
  wire       [35:0]   _zz_788;
  wire       [0:0]    _zz_789;
  wire       [0:0]    _zz_790;
  wire       [35:0]   _zz_791;
  wire       [35:0]   _zz_792;
  wire       [35:0]   _zz_793;
  wire       [0:0]    _zz_794;
  wire       [0:0]    _zz_795;
  wire       [35:0]   _zz_796;
  wire       [35:0]   _zz_797;
  wire       [35:0]   _zz_798;
  wire       [0:0]    _zz_799;
  wire       [0:0]    _zz_800;
  wire       [35:0]   _zz_801;
  wire       [35:0]   _zz_802;
  wire       [35:0]   _zz_803;
  wire       [0:0]    _zz_804;
  wire       [0:0]    _zz_805;
  wire       [35:0]   _zz_806;
  wire       [35:0]   _zz_807;
  wire       [35:0]   _zz_808;
  wire       [0:0]    _zz_809;
  wire       [0:0]    _zz_810;
  wire       [35:0]   _zz_811;
  wire       [35:0]   _zz_812;
  wire       [35:0]   _zz_813;
  wire       [0:0]    _zz_814;
  wire       [0:0]    _zz_815;
  wire       [35:0]   _zz_816;
  wire       [35:0]   _zz_817;
  wire       [35:0]   _zz_818;
  wire       [0:0]    _zz_819;
  wire       [0:0]    _zz_820;
  wire       [35:0]   _zz_821;
  wire       [35:0]   _zz_822;
  wire       [35:0]   _zz_823;
  wire       [0:0]    _zz_824;
  wire       [0:0]    _zz_825;
  wire       [35:0]   _zz_826;
  wire       [35:0]   _zz_827;
  wire       [35:0]   _zz_828;
  wire       [0:0]    _zz_829;
  wire       [0:0]    _zz_830;
  wire       [35:0]   _zz_831;
  wire       [35:0]   _zz_832;
  wire       [35:0]   _zz_833;
  wire       [0:0]    _zz_834;
  wire       [0:0]    _zz_835;
  wire       [35:0]   _zz_836;
  wire       [35:0]   _zz_837;
  wire       [35:0]   _zz_838;
  wire       [0:0]    _zz_839;
  wire       [0:0]    _zz_840;
  wire       [35:0]   _zz_841;
  wire       [35:0]   _zz_842;
  wire       [35:0]   _zz_843;
  wire       [0:0]    _zz_844;
  wire       [0:0]    _zz_845;
  wire       [35:0]   _zz_846;
  wire       [35:0]   _zz_847;
  wire       [35:0]   _zz_848;
  wire       [0:0]    _zz_849;
  wire       [0:0]    _zz_850;
  wire       [35:0]   _zz_851;
  wire       [35:0]   _zz_852;
  wire       [35:0]   _zz_853;
  wire       [0:0]    _zz_854;
  wire       [0:0]    _zz_855;
  wire       [35:0]   _zz_856;
  wire       [35:0]   _zz_857;
  wire       [35:0]   _zz_858;
  wire       [0:0]    _zz_859;
  wire       [0:0]    _zz_860;
  wire       [35:0]   _zz_861;
  wire       [35:0]   _zz_862;
  wire       [35:0]   _zz_863;
  wire       [0:0]    _zz_864;
  wire       [0:0]    _zz_865;
  wire       [35:0]   _zz_866;
  wire       [35:0]   _zz_867;
  wire       [35:0]   _zz_868;
  wire       [0:0]    _zz_869;
  wire       [0:0]    _zz_870;
  wire       [35:0]   _zz_871;
  wire       [35:0]   _zz_872;
  wire       [35:0]   _zz_873;
  wire       [0:0]    _zz_874;
  wire       [0:0]    _zz_875;
  wire       [35:0]   _zz_876;
  wire       [35:0]   _zz_877;
  wire       [35:0]   _zz_878;
  wire       [0:0]    _zz_879;
  wire       [0:0]    _zz_880;
  wire       [35:0]   _zz_881;
  wire       [35:0]   _zz_882;
  wire       [35:0]   _zz_883;
  wire       [0:0]    _zz_884;
  wire       [0:0]    _zz_885;
  wire       [35:0]   _zz_886;
  wire       [35:0]   _zz_887;
  wire       [35:0]   _zz_888;
  wire       [0:0]    _zz_889;
  wire       [0:0]    _zz_890;
  wire       [35:0]   _zz_891;
  wire       [35:0]   _zz_892;
  wire       [35:0]   _zz_893;
  wire       [0:0]    _zz_894;
  wire       [0:0]    _zz_895;
  wire       [35:0]   _zz_896;
  wire       [35:0]   _zz_897;
  wire       [35:0]   _zz_898;
  wire       [0:0]    _zz_899;
  wire       [0:0]    _zz_900;
  wire       [35:0]   _zz_901;
  wire       [35:0]   _zz_902;
  wire       [35:0]   _zz_903;
  wire       [0:0]    _zz_904;
  wire       [0:0]    _zz_905;
  wire       [35:0]   _zz_906;
  wire       [35:0]   _zz_907;
  wire       [35:0]   _zz_908;
  wire       [0:0]    _zz_909;
  wire       [0:0]    _zz_910;
  wire       [35:0]   _zz_911;
  wire       [35:0]   _zz_912;
  wire       [35:0]   _zz_913;
  wire       [0:0]    _zz_914;
  wire       [0:0]    _zz_915;
  wire       [35:0]   _zz_916;
  wire       [35:0]   _zz_917;
  wire       [35:0]   _zz_918;
  wire       [0:0]    _zz_919;
  wire       [0:0]    _zz_920;
  wire       [35:0]   _zz_921;
  wire       [35:0]   _zz_922;
  wire       [35:0]   _zz_923;
  wire       [0:0]    _zz_924;
  wire       [0:0]    _zz_925;
  wire       [35:0]   _zz_926;
  wire       [35:0]   _zz_927;
  wire       [35:0]   _zz_928;
  wire       [0:0]    _zz_929;
  wire       [0:0]    _zz_930;
  wire       [35:0]   _zz_931;
  wire       [35:0]   _zz_932;
  wire       [35:0]   _zz_933;
  wire       [0:0]    _zz_934;
  wire       [0:0]    _zz_935;
  wire       [35:0]   _zz_936;
  wire       [35:0]   _zz_937;
  wire       [35:0]   _zz_938;
  wire       [0:0]    _zz_939;
  wire       [0:0]    _zz_940;
  wire       [35:0]   _zz_941;
  wire       [35:0]   _zz_942;
  wire       [35:0]   _zz_943;
  wire       [0:0]    _zz_944;
  wire       [0:0]    _zz_945;
  wire       [35:0]   _zz_946;
  wire       [35:0]   _zz_947;
  wire       [35:0]   _zz_948;
  wire       [0:0]    _zz_949;
  wire       [0:0]    _zz_950;
  wire       [35:0]   _zz_951;
  wire       [35:0]   _zz_952;
  wire       [35:0]   _zz_953;
  wire       [0:0]    _zz_954;
  wire       [0:0]    _zz_955;
  wire       [35:0]   _zz_956;
  wire       [35:0]   _zz_957;
  wire       [35:0]   _zz_958;
  wire       [0:0]    _zz_959;
  wire       [0:0]    _zz_960;
  reg                 io_data_in_valid_delay_1;
  reg                 io_data_in_valid_delay_2;
  reg                 io_data_in_valid_delay_3;
  reg                 io_data_in_valid_delay_4;
  reg                 io_data_in_valid_delay_5;
  reg                 io_data_in_valid_delay_6;
  reg                 io_data_in_valid_delay_7;
  reg                 io_data_in_valid_delay_8;

  assign _zz_2113 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2114 = ($signed(_zz_3) - $signed(_zz_2115));
  assign _zz_2115 = ($signed(_zz_2116) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2116 = ($signed(data_mid_0_1_real) + $signed(data_mid_0_1_imag));
  assign _zz_2117 = fixTo_dout;
  assign _zz_2118 = ($signed(_zz_3) + $signed(_zz_2119));
  assign _zz_2119 = ($signed(_zz_2120) * $signed(twiddle_factor_table_0_real));
  assign _zz_2120 = ($signed(data_mid_0_1_imag) - $signed(data_mid_0_1_real));
  assign _zz_2121 = fixTo_1_dout;
  assign _zz_2122 = _zz_2123[35 : 0];
  assign _zz_2123 = _zz_2124;
  assign _zz_2124 = ($signed(_zz_2125) >>> _zz_4);
  assign _zz_2125 = _zz_2126;
  assign _zz_2126 = ($signed(_zz_2128) - $signed(_zz_1));
  assign _zz_2127 = ({9'd0,data_mid_0_0_real} <<< 9);
  assign _zz_2128 = {{9{_zz_2127[26]}}, _zz_2127};
  assign _zz_2129 = fixTo_2_dout;
  assign _zz_2130 = _zz_2131[35 : 0];
  assign _zz_2131 = _zz_2132;
  assign _zz_2132 = ($signed(_zz_2133) >>> _zz_4);
  assign _zz_2133 = _zz_2134;
  assign _zz_2134 = ($signed(_zz_2136) - $signed(_zz_2));
  assign _zz_2135 = ({9'd0,data_mid_0_0_imag} <<< 9);
  assign _zz_2136 = {{9{_zz_2135[26]}}, _zz_2135};
  assign _zz_2137 = fixTo_3_dout;
  assign _zz_2138 = _zz_2139[35 : 0];
  assign _zz_2139 = _zz_2140;
  assign _zz_2140 = ($signed(_zz_2141) >>> _zz_5);
  assign _zz_2141 = _zz_2142;
  assign _zz_2142 = ($signed(_zz_2144) + $signed(_zz_1));
  assign _zz_2143 = ({9'd0,data_mid_0_0_real} <<< 9);
  assign _zz_2144 = {{9{_zz_2143[26]}}, _zz_2143};
  assign _zz_2145 = fixTo_4_dout;
  assign _zz_2146 = _zz_2147[35 : 0];
  assign _zz_2147 = _zz_2148;
  assign _zz_2148 = ($signed(_zz_2149) >>> _zz_5);
  assign _zz_2149 = _zz_2150;
  assign _zz_2150 = ($signed(_zz_2152) + $signed(_zz_2));
  assign _zz_2151 = ({9'd0,data_mid_0_0_imag} <<< 9);
  assign _zz_2152 = {{9{_zz_2151[26]}}, _zz_2151};
  assign _zz_2153 = fixTo_5_dout;
  assign _zz_2154 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2155 = ($signed(_zz_8) - $signed(_zz_2156));
  assign _zz_2156 = ($signed(_zz_2157) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2157 = ($signed(data_mid_0_3_real) + $signed(data_mid_0_3_imag));
  assign _zz_2158 = fixTo_6_dout;
  assign _zz_2159 = ($signed(_zz_8) + $signed(_zz_2160));
  assign _zz_2160 = ($signed(_zz_2161) * $signed(twiddle_factor_table_0_real));
  assign _zz_2161 = ($signed(data_mid_0_3_imag) - $signed(data_mid_0_3_real));
  assign _zz_2162 = fixTo_7_dout;
  assign _zz_2163 = _zz_2164[35 : 0];
  assign _zz_2164 = _zz_2165;
  assign _zz_2165 = ($signed(_zz_2166) >>> _zz_9);
  assign _zz_2166 = _zz_2167;
  assign _zz_2167 = ($signed(_zz_2169) - $signed(_zz_6));
  assign _zz_2168 = ({9'd0,data_mid_0_2_real} <<< 9);
  assign _zz_2169 = {{9{_zz_2168[26]}}, _zz_2168};
  assign _zz_2170 = fixTo_8_dout;
  assign _zz_2171 = _zz_2172[35 : 0];
  assign _zz_2172 = _zz_2173;
  assign _zz_2173 = ($signed(_zz_2174) >>> _zz_9);
  assign _zz_2174 = _zz_2175;
  assign _zz_2175 = ($signed(_zz_2177) - $signed(_zz_7));
  assign _zz_2176 = ({9'd0,data_mid_0_2_imag} <<< 9);
  assign _zz_2177 = {{9{_zz_2176[26]}}, _zz_2176};
  assign _zz_2178 = fixTo_9_dout;
  assign _zz_2179 = _zz_2180[35 : 0];
  assign _zz_2180 = _zz_2181;
  assign _zz_2181 = ($signed(_zz_2182) >>> _zz_10);
  assign _zz_2182 = _zz_2183;
  assign _zz_2183 = ($signed(_zz_2185) + $signed(_zz_6));
  assign _zz_2184 = ({9'd0,data_mid_0_2_real} <<< 9);
  assign _zz_2185 = {{9{_zz_2184[26]}}, _zz_2184};
  assign _zz_2186 = fixTo_10_dout;
  assign _zz_2187 = _zz_2188[35 : 0];
  assign _zz_2188 = _zz_2189;
  assign _zz_2189 = ($signed(_zz_2190) >>> _zz_10);
  assign _zz_2190 = _zz_2191;
  assign _zz_2191 = ($signed(_zz_2193) + $signed(_zz_7));
  assign _zz_2192 = ({9'd0,data_mid_0_2_imag} <<< 9);
  assign _zz_2193 = {{9{_zz_2192[26]}}, _zz_2192};
  assign _zz_2194 = fixTo_11_dout;
  assign _zz_2195 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2196 = ($signed(_zz_13) - $signed(_zz_2197));
  assign _zz_2197 = ($signed(_zz_2198) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2198 = ($signed(data_mid_0_5_real) + $signed(data_mid_0_5_imag));
  assign _zz_2199 = fixTo_12_dout;
  assign _zz_2200 = ($signed(_zz_13) + $signed(_zz_2201));
  assign _zz_2201 = ($signed(_zz_2202) * $signed(twiddle_factor_table_0_real));
  assign _zz_2202 = ($signed(data_mid_0_5_imag) - $signed(data_mid_0_5_real));
  assign _zz_2203 = fixTo_13_dout;
  assign _zz_2204 = _zz_2205[35 : 0];
  assign _zz_2205 = _zz_2206;
  assign _zz_2206 = ($signed(_zz_2207) >>> _zz_14);
  assign _zz_2207 = _zz_2208;
  assign _zz_2208 = ($signed(_zz_2210) - $signed(_zz_11));
  assign _zz_2209 = ({9'd0,data_mid_0_4_real} <<< 9);
  assign _zz_2210 = {{9{_zz_2209[26]}}, _zz_2209};
  assign _zz_2211 = fixTo_14_dout;
  assign _zz_2212 = _zz_2213[35 : 0];
  assign _zz_2213 = _zz_2214;
  assign _zz_2214 = ($signed(_zz_2215) >>> _zz_14);
  assign _zz_2215 = _zz_2216;
  assign _zz_2216 = ($signed(_zz_2218) - $signed(_zz_12));
  assign _zz_2217 = ({9'd0,data_mid_0_4_imag} <<< 9);
  assign _zz_2218 = {{9{_zz_2217[26]}}, _zz_2217};
  assign _zz_2219 = fixTo_15_dout;
  assign _zz_2220 = _zz_2221[35 : 0];
  assign _zz_2221 = _zz_2222;
  assign _zz_2222 = ($signed(_zz_2223) >>> _zz_15);
  assign _zz_2223 = _zz_2224;
  assign _zz_2224 = ($signed(_zz_2226) + $signed(_zz_11));
  assign _zz_2225 = ({9'd0,data_mid_0_4_real} <<< 9);
  assign _zz_2226 = {{9{_zz_2225[26]}}, _zz_2225};
  assign _zz_2227 = fixTo_16_dout;
  assign _zz_2228 = _zz_2229[35 : 0];
  assign _zz_2229 = _zz_2230;
  assign _zz_2230 = ($signed(_zz_2231) >>> _zz_15);
  assign _zz_2231 = _zz_2232;
  assign _zz_2232 = ($signed(_zz_2234) + $signed(_zz_12));
  assign _zz_2233 = ({9'd0,data_mid_0_4_imag} <<< 9);
  assign _zz_2234 = {{9{_zz_2233[26]}}, _zz_2233};
  assign _zz_2235 = fixTo_17_dout;
  assign _zz_2236 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2237 = ($signed(_zz_18) - $signed(_zz_2238));
  assign _zz_2238 = ($signed(_zz_2239) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2239 = ($signed(data_mid_0_7_real) + $signed(data_mid_0_7_imag));
  assign _zz_2240 = fixTo_18_dout;
  assign _zz_2241 = ($signed(_zz_18) + $signed(_zz_2242));
  assign _zz_2242 = ($signed(_zz_2243) * $signed(twiddle_factor_table_0_real));
  assign _zz_2243 = ($signed(data_mid_0_7_imag) - $signed(data_mid_0_7_real));
  assign _zz_2244 = fixTo_19_dout;
  assign _zz_2245 = _zz_2246[35 : 0];
  assign _zz_2246 = _zz_2247;
  assign _zz_2247 = ($signed(_zz_2248) >>> _zz_19);
  assign _zz_2248 = _zz_2249;
  assign _zz_2249 = ($signed(_zz_2251) - $signed(_zz_16));
  assign _zz_2250 = ({9'd0,data_mid_0_6_real} <<< 9);
  assign _zz_2251 = {{9{_zz_2250[26]}}, _zz_2250};
  assign _zz_2252 = fixTo_20_dout;
  assign _zz_2253 = _zz_2254[35 : 0];
  assign _zz_2254 = _zz_2255;
  assign _zz_2255 = ($signed(_zz_2256) >>> _zz_19);
  assign _zz_2256 = _zz_2257;
  assign _zz_2257 = ($signed(_zz_2259) - $signed(_zz_17));
  assign _zz_2258 = ({9'd0,data_mid_0_6_imag} <<< 9);
  assign _zz_2259 = {{9{_zz_2258[26]}}, _zz_2258};
  assign _zz_2260 = fixTo_21_dout;
  assign _zz_2261 = _zz_2262[35 : 0];
  assign _zz_2262 = _zz_2263;
  assign _zz_2263 = ($signed(_zz_2264) >>> _zz_20);
  assign _zz_2264 = _zz_2265;
  assign _zz_2265 = ($signed(_zz_2267) + $signed(_zz_16));
  assign _zz_2266 = ({9'd0,data_mid_0_6_real} <<< 9);
  assign _zz_2267 = {{9{_zz_2266[26]}}, _zz_2266};
  assign _zz_2268 = fixTo_22_dout;
  assign _zz_2269 = _zz_2270[35 : 0];
  assign _zz_2270 = _zz_2271;
  assign _zz_2271 = ($signed(_zz_2272) >>> _zz_20);
  assign _zz_2272 = _zz_2273;
  assign _zz_2273 = ($signed(_zz_2275) + $signed(_zz_17));
  assign _zz_2274 = ({9'd0,data_mid_0_6_imag} <<< 9);
  assign _zz_2275 = {{9{_zz_2274[26]}}, _zz_2274};
  assign _zz_2276 = fixTo_23_dout;
  assign _zz_2277 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2278 = ($signed(_zz_23) - $signed(_zz_2279));
  assign _zz_2279 = ($signed(_zz_2280) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2280 = ($signed(data_mid_0_9_real) + $signed(data_mid_0_9_imag));
  assign _zz_2281 = fixTo_24_dout;
  assign _zz_2282 = ($signed(_zz_23) + $signed(_zz_2283));
  assign _zz_2283 = ($signed(_zz_2284) * $signed(twiddle_factor_table_0_real));
  assign _zz_2284 = ($signed(data_mid_0_9_imag) - $signed(data_mid_0_9_real));
  assign _zz_2285 = fixTo_25_dout;
  assign _zz_2286 = _zz_2287[35 : 0];
  assign _zz_2287 = _zz_2288;
  assign _zz_2288 = ($signed(_zz_2289) >>> _zz_24);
  assign _zz_2289 = _zz_2290;
  assign _zz_2290 = ($signed(_zz_2292) - $signed(_zz_21));
  assign _zz_2291 = ({9'd0,data_mid_0_8_real} <<< 9);
  assign _zz_2292 = {{9{_zz_2291[26]}}, _zz_2291};
  assign _zz_2293 = fixTo_26_dout;
  assign _zz_2294 = _zz_2295[35 : 0];
  assign _zz_2295 = _zz_2296;
  assign _zz_2296 = ($signed(_zz_2297) >>> _zz_24);
  assign _zz_2297 = _zz_2298;
  assign _zz_2298 = ($signed(_zz_2300) - $signed(_zz_22));
  assign _zz_2299 = ({9'd0,data_mid_0_8_imag} <<< 9);
  assign _zz_2300 = {{9{_zz_2299[26]}}, _zz_2299};
  assign _zz_2301 = fixTo_27_dout;
  assign _zz_2302 = _zz_2303[35 : 0];
  assign _zz_2303 = _zz_2304;
  assign _zz_2304 = ($signed(_zz_2305) >>> _zz_25);
  assign _zz_2305 = _zz_2306;
  assign _zz_2306 = ($signed(_zz_2308) + $signed(_zz_21));
  assign _zz_2307 = ({9'd0,data_mid_0_8_real} <<< 9);
  assign _zz_2308 = {{9{_zz_2307[26]}}, _zz_2307};
  assign _zz_2309 = fixTo_28_dout;
  assign _zz_2310 = _zz_2311[35 : 0];
  assign _zz_2311 = _zz_2312;
  assign _zz_2312 = ($signed(_zz_2313) >>> _zz_25);
  assign _zz_2313 = _zz_2314;
  assign _zz_2314 = ($signed(_zz_2316) + $signed(_zz_22));
  assign _zz_2315 = ({9'd0,data_mid_0_8_imag} <<< 9);
  assign _zz_2316 = {{9{_zz_2315[26]}}, _zz_2315};
  assign _zz_2317 = fixTo_29_dout;
  assign _zz_2318 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2319 = ($signed(_zz_28) - $signed(_zz_2320));
  assign _zz_2320 = ($signed(_zz_2321) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2321 = ($signed(data_mid_0_11_real) + $signed(data_mid_0_11_imag));
  assign _zz_2322 = fixTo_30_dout;
  assign _zz_2323 = ($signed(_zz_28) + $signed(_zz_2324));
  assign _zz_2324 = ($signed(_zz_2325) * $signed(twiddle_factor_table_0_real));
  assign _zz_2325 = ($signed(data_mid_0_11_imag) - $signed(data_mid_0_11_real));
  assign _zz_2326 = fixTo_31_dout;
  assign _zz_2327 = _zz_2328[35 : 0];
  assign _zz_2328 = _zz_2329;
  assign _zz_2329 = ($signed(_zz_2330) >>> _zz_29);
  assign _zz_2330 = _zz_2331;
  assign _zz_2331 = ($signed(_zz_2333) - $signed(_zz_26));
  assign _zz_2332 = ({9'd0,data_mid_0_10_real} <<< 9);
  assign _zz_2333 = {{9{_zz_2332[26]}}, _zz_2332};
  assign _zz_2334 = fixTo_32_dout;
  assign _zz_2335 = _zz_2336[35 : 0];
  assign _zz_2336 = _zz_2337;
  assign _zz_2337 = ($signed(_zz_2338) >>> _zz_29);
  assign _zz_2338 = _zz_2339;
  assign _zz_2339 = ($signed(_zz_2341) - $signed(_zz_27));
  assign _zz_2340 = ({9'd0,data_mid_0_10_imag} <<< 9);
  assign _zz_2341 = {{9{_zz_2340[26]}}, _zz_2340};
  assign _zz_2342 = fixTo_33_dout;
  assign _zz_2343 = _zz_2344[35 : 0];
  assign _zz_2344 = _zz_2345;
  assign _zz_2345 = ($signed(_zz_2346) >>> _zz_30);
  assign _zz_2346 = _zz_2347;
  assign _zz_2347 = ($signed(_zz_2349) + $signed(_zz_26));
  assign _zz_2348 = ({9'd0,data_mid_0_10_real} <<< 9);
  assign _zz_2349 = {{9{_zz_2348[26]}}, _zz_2348};
  assign _zz_2350 = fixTo_34_dout;
  assign _zz_2351 = _zz_2352[35 : 0];
  assign _zz_2352 = _zz_2353;
  assign _zz_2353 = ($signed(_zz_2354) >>> _zz_30);
  assign _zz_2354 = _zz_2355;
  assign _zz_2355 = ($signed(_zz_2357) + $signed(_zz_27));
  assign _zz_2356 = ({9'd0,data_mid_0_10_imag} <<< 9);
  assign _zz_2357 = {{9{_zz_2356[26]}}, _zz_2356};
  assign _zz_2358 = fixTo_35_dout;
  assign _zz_2359 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2360 = ($signed(_zz_33) - $signed(_zz_2361));
  assign _zz_2361 = ($signed(_zz_2362) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2362 = ($signed(data_mid_0_13_real) + $signed(data_mid_0_13_imag));
  assign _zz_2363 = fixTo_36_dout;
  assign _zz_2364 = ($signed(_zz_33) + $signed(_zz_2365));
  assign _zz_2365 = ($signed(_zz_2366) * $signed(twiddle_factor_table_0_real));
  assign _zz_2366 = ($signed(data_mid_0_13_imag) - $signed(data_mid_0_13_real));
  assign _zz_2367 = fixTo_37_dout;
  assign _zz_2368 = _zz_2369[35 : 0];
  assign _zz_2369 = _zz_2370;
  assign _zz_2370 = ($signed(_zz_2371) >>> _zz_34);
  assign _zz_2371 = _zz_2372;
  assign _zz_2372 = ($signed(_zz_2374) - $signed(_zz_31));
  assign _zz_2373 = ({9'd0,data_mid_0_12_real} <<< 9);
  assign _zz_2374 = {{9{_zz_2373[26]}}, _zz_2373};
  assign _zz_2375 = fixTo_38_dout;
  assign _zz_2376 = _zz_2377[35 : 0];
  assign _zz_2377 = _zz_2378;
  assign _zz_2378 = ($signed(_zz_2379) >>> _zz_34);
  assign _zz_2379 = _zz_2380;
  assign _zz_2380 = ($signed(_zz_2382) - $signed(_zz_32));
  assign _zz_2381 = ({9'd0,data_mid_0_12_imag} <<< 9);
  assign _zz_2382 = {{9{_zz_2381[26]}}, _zz_2381};
  assign _zz_2383 = fixTo_39_dout;
  assign _zz_2384 = _zz_2385[35 : 0];
  assign _zz_2385 = _zz_2386;
  assign _zz_2386 = ($signed(_zz_2387) >>> _zz_35);
  assign _zz_2387 = _zz_2388;
  assign _zz_2388 = ($signed(_zz_2390) + $signed(_zz_31));
  assign _zz_2389 = ({9'd0,data_mid_0_12_real} <<< 9);
  assign _zz_2390 = {{9{_zz_2389[26]}}, _zz_2389};
  assign _zz_2391 = fixTo_40_dout;
  assign _zz_2392 = _zz_2393[35 : 0];
  assign _zz_2393 = _zz_2394;
  assign _zz_2394 = ($signed(_zz_2395) >>> _zz_35);
  assign _zz_2395 = _zz_2396;
  assign _zz_2396 = ($signed(_zz_2398) + $signed(_zz_32));
  assign _zz_2397 = ({9'd0,data_mid_0_12_imag} <<< 9);
  assign _zz_2398 = {{9{_zz_2397[26]}}, _zz_2397};
  assign _zz_2399 = fixTo_41_dout;
  assign _zz_2400 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2401 = ($signed(_zz_38) - $signed(_zz_2402));
  assign _zz_2402 = ($signed(_zz_2403) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2403 = ($signed(data_mid_0_15_real) + $signed(data_mid_0_15_imag));
  assign _zz_2404 = fixTo_42_dout;
  assign _zz_2405 = ($signed(_zz_38) + $signed(_zz_2406));
  assign _zz_2406 = ($signed(_zz_2407) * $signed(twiddle_factor_table_0_real));
  assign _zz_2407 = ($signed(data_mid_0_15_imag) - $signed(data_mid_0_15_real));
  assign _zz_2408 = fixTo_43_dout;
  assign _zz_2409 = _zz_2410[35 : 0];
  assign _zz_2410 = _zz_2411;
  assign _zz_2411 = ($signed(_zz_2412) >>> _zz_39);
  assign _zz_2412 = _zz_2413;
  assign _zz_2413 = ($signed(_zz_2415) - $signed(_zz_36));
  assign _zz_2414 = ({9'd0,data_mid_0_14_real} <<< 9);
  assign _zz_2415 = {{9{_zz_2414[26]}}, _zz_2414};
  assign _zz_2416 = fixTo_44_dout;
  assign _zz_2417 = _zz_2418[35 : 0];
  assign _zz_2418 = _zz_2419;
  assign _zz_2419 = ($signed(_zz_2420) >>> _zz_39);
  assign _zz_2420 = _zz_2421;
  assign _zz_2421 = ($signed(_zz_2423) - $signed(_zz_37));
  assign _zz_2422 = ({9'd0,data_mid_0_14_imag} <<< 9);
  assign _zz_2423 = {{9{_zz_2422[26]}}, _zz_2422};
  assign _zz_2424 = fixTo_45_dout;
  assign _zz_2425 = _zz_2426[35 : 0];
  assign _zz_2426 = _zz_2427;
  assign _zz_2427 = ($signed(_zz_2428) >>> _zz_40);
  assign _zz_2428 = _zz_2429;
  assign _zz_2429 = ($signed(_zz_2431) + $signed(_zz_36));
  assign _zz_2430 = ({9'd0,data_mid_0_14_real} <<< 9);
  assign _zz_2431 = {{9{_zz_2430[26]}}, _zz_2430};
  assign _zz_2432 = fixTo_46_dout;
  assign _zz_2433 = _zz_2434[35 : 0];
  assign _zz_2434 = _zz_2435;
  assign _zz_2435 = ($signed(_zz_2436) >>> _zz_40);
  assign _zz_2436 = _zz_2437;
  assign _zz_2437 = ($signed(_zz_2439) + $signed(_zz_37));
  assign _zz_2438 = ({9'd0,data_mid_0_14_imag} <<< 9);
  assign _zz_2439 = {{9{_zz_2438[26]}}, _zz_2438};
  assign _zz_2440 = fixTo_47_dout;
  assign _zz_2441 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2442 = ($signed(_zz_43) - $signed(_zz_2443));
  assign _zz_2443 = ($signed(_zz_2444) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2444 = ($signed(data_mid_0_17_real) + $signed(data_mid_0_17_imag));
  assign _zz_2445 = fixTo_48_dout;
  assign _zz_2446 = ($signed(_zz_43) + $signed(_zz_2447));
  assign _zz_2447 = ($signed(_zz_2448) * $signed(twiddle_factor_table_0_real));
  assign _zz_2448 = ($signed(data_mid_0_17_imag) - $signed(data_mid_0_17_real));
  assign _zz_2449 = fixTo_49_dout;
  assign _zz_2450 = _zz_2451[35 : 0];
  assign _zz_2451 = _zz_2452;
  assign _zz_2452 = ($signed(_zz_2453) >>> _zz_44);
  assign _zz_2453 = _zz_2454;
  assign _zz_2454 = ($signed(_zz_2456) - $signed(_zz_41));
  assign _zz_2455 = ({9'd0,data_mid_0_16_real} <<< 9);
  assign _zz_2456 = {{9{_zz_2455[26]}}, _zz_2455};
  assign _zz_2457 = fixTo_50_dout;
  assign _zz_2458 = _zz_2459[35 : 0];
  assign _zz_2459 = _zz_2460;
  assign _zz_2460 = ($signed(_zz_2461) >>> _zz_44);
  assign _zz_2461 = _zz_2462;
  assign _zz_2462 = ($signed(_zz_2464) - $signed(_zz_42));
  assign _zz_2463 = ({9'd0,data_mid_0_16_imag} <<< 9);
  assign _zz_2464 = {{9{_zz_2463[26]}}, _zz_2463};
  assign _zz_2465 = fixTo_51_dout;
  assign _zz_2466 = _zz_2467[35 : 0];
  assign _zz_2467 = _zz_2468;
  assign _zz_2468 = ($signed(_zz_2469) >>> _zz_45);
  assign _zz_2469 = _zz_2470;
  assign _zz_2470 = ($signed(_zz_2472) + $signed(_zz_41));
  assign _zz_2471 = ({9'd0,data_mid_0_16_real} <<< 9);
  assign _zz_2472 = {{9{_zz_2471[26]}}, _zz_2471};
  assign _zz_2473 = fixTo_52_dout;
  assign _zz_2474 = _zz_2475[35 : 0];
  assign _zz_2475 = _zz_2476;
  assign _zz_2476 = ($signed(_zz_2477) >>> _zz_45);
  assign _zz_2477 = _zz_2478;
  assign _zz_2478 = ($signed(_zz_2480) + $signed(_zz_42));
  assign _zz_2479 = ({9'd0,data_mid_0_16_imag} <<< 9);
  assign _zz_2480 = {{9{_zz_2479[26]}}, _zz_2479};
  assign _zz_2481 = fixTo_53_dout;
  assign _zz_2482 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2483 = ($signed(_zz_48) - $signed(_zz_2484));
  assign _zz_2484 = ($signed(_zz_2485) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2485 = ($signed(data_mid_0_19_real) + $signed(data_mid_0_19_imag));
  assign _zz_2486 = fixTo_54_dout;
  assign _zz_2487 = ($signed(_zz_48) + $signed(_zz_2488));
  assign _zz_2488 = ($signed(_zz_2489) * $signed(twiddle_factor_table_0_real));
  assign _zz_2489 = ($signed(data_mid_0_19_imag) - $signed(data_mid_0_19_real));
  assign _zz_2490 = fixTo_55_dout;
  assign _zz_2491 = _zz_2492[35 : 0];
  assign _zz_2492 = _zz_2493;
  assign _zz_2493 = ($signed(_zz_2494) >>> _zz_49);
  assign _zz_2494 = _zz_2495;
  assign _zz_2495 = ($signed(_zz_2497) - $signed(_zz_46));
  assign _zz_2496 = ({9'd0,data_mid_0_18_real} <<< 9);
  assign _zz_2497 = {{9{_zz_2496[26]}}, _zz_2496};
  assign _zz_2498 = fixTo_56_dout;
  assign _zz_2499 = _zz_2500[35 : 0];
  assign _zz_2500 = _zz_2501;
  assign _zz_2501 = ($signed(_zz_2502) >>> _zz_49);
  assign _zz_2502 = _zz_2503;
  assign _zz_2503 = ($signed(_zz_2505) - $signed(_zz_47));
  assign _zz_2504 = ({9'd0,data_mid_0_18_imag} <<< 9);
  assign _zz_2505 = {{9{_zz_2504[26]}}, _zz_2504};
  assign _zz_2506 = fixTo_57_dout;
  assign _zz_2507 = _zz_2508[35 : 0];
  assign _zz_2508 = _zz_2509;
  assign _zz_2509 = ($signed(_zz_2510) >>> _zz_50);
  assign _zz_2510 = _zz_2511;
  assign _zz_2511 = ($signed(_zz_2513) + $signed(_zz_46));
  assign _zz_2512 = ({9'd0,data_mid_0_18_real} <<< 9);
  assign _zz_2513 = {{9{_zz_2512[26]}}, _zz_2512};
  assign _zz_2514 = fixTo_58_dout;
  assign _zz_2515 = _zz_2516[35 : 0];
  assign _zz_2516 = _zz_2517;
  assign _zz_2517 = ($signed(_zz_2518) >>> _zz_50);
  assign _zz_2518 = _zz_2519;
  assign _zz_2519 = ($signed(_zz_2521) + $signed(_zz_47));
  assign _zz_2520 = ({9'd0,data_mid_0_18_imag} <<< 9);
  assign _zz_2521 = {{9{_zz_2520[26]}}, _zz_2520};
  assign _zz_2522 = fixTo_59_dout;
  assign _zz_2523 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2524 = ($signed(_zz_53) - $signed(_zz_2525));
  assign _zz_2525 = ($signed(_zz_2526) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2526 = ($signed(data_mid_0_21_real) + $signed(data_mid_0_21_imag));
  assign _zz_2527 = fixTo_60_dout;
  assign _zz_2528 = ($signed(_zz_53) + $signed(_zz_2529));
  assign _zz_2529 = ($signed(_zz_2530) * $signed(twiddle_factor_table_0_real));
  assign _zz_2530 = ($signed(data_mid_0_21_imag) - $signed(data_mid_0_21_real));
  assign _zz_2531 = fixTo_61_dout;
  assign _zz_2532 = _zz_2533[35 : 0];
  assign _zz_2533 = _zz_2534;
  assign _zz_2534 = ($signed(_zz_2535) >>> _zz_54);
  assign _zz_2535 = _zz_2536;
  assign _zz_2536 = ($signed(_zz_2538) - $signed(_zz_51));
  assign _zz_2537 = ({9'd0,data_mid_0_20_real} <<< 9);
  assign _zz_2538 = {{9{_zz_2537[26]}}, _zz_2537};
  assign _zz_2539 = fixTo_62_dout;
  assign _zz_2540 = _zz_2541[35 : 0];
  assign _zz_2541 = _zz_2542;
  assign _zz_2542 = ($signed(_zz_2543) >>> _zz_54);
  assign _zz_2543 = _zz_2544;
  assign _zz_2544 = ($signed(_zz_2546) - $signed(_zz_52));
  assign _zz_2545 = ({9'd0,data_mid_0_20_imag} <<< 9);
  assign _zz_2546 = {{9{_zz_2545[26]}}, _zz_2545};
  assign _zz_2547 = fixTo_63_dout;
  assign _zz_2548 = _zz_2549[35 : 0];
  assign _zz_2549 = _zz_2550;
  assign _zz_2550 = ($signed(_zz_2551) >>> _zz_55);
  assign _zz_2551 = _zz_2552;
  assign _zz_2552 = ($signed(_zz_2554) + $signed(_zz_51));
  assign _zz_2553 = ({9'd0,data_mid_0_20_real} <<< 9);
  assign _zz_2554 = {{9{_zz_2553[26]}}, _zz_2553};
  assign _zz_2555 = fixTo_64_dout;
  assign _zz_2556 = _zz_2557[35 : 0];
  assign _zz_2557 = _zz_2558;
  assign _zz_2558 = ($signed(_zz_2559) >>> _zz_55);
  assign _zz_2559 = _zz_2560;
  assign _zz_2560 = ($signed(_zz_2562) + $signed(_zz_52));
  assign _zz_2561 = ({9'd0,data_mid_0_20_imag} <<< 9);
  assign _zz_2562 = {{9{_zz_2561[26]}}, _zz_2561};
  assign _zz_2563 = fixTo_65_dout;
  assign _zz_2564 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2565 = ($signed(_zz_58) - $signed(_zz_2566));
  assign _zz_2566 = ($signed(_zz_2567) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2567 = ($signed(data_mid_0_23_real) + $signed(data_mid_0_23_imag));
  assign _zz_2568 = fixTo_66_dout;
  assign _zz_2569 = ($signed(_zz_58) + $signed(_zz_2570));
  assign _zz_2570 = ($signed(_zz_2571) * $signed(twiddle_factor_table_0_real));
  assign _zz_2571 = ($signed(data_mid_0_23_imag) - $signed(data_mid_0_23_real));
  assign _zz_2572 = fixTo_67_dout;
  assign _zz_2573 = _zz_2574[35 : 0];
  assign _zz_2574 = _zz_2575;
  assign _zz_2575 = ($signed(_zz_2576) >>> _zz_59);
  assign _zz_2576 = _zz_2577;
  assign _zz_2577 = ($signed(_zz_2579) - $signed(_zz_56));
  assign _zz_2578 = ({9'd0,data_mid_0_22_real} <<< 9);
  assign _zz_2579 = {{9{_zz_2578[26]}}, _zz_2578};
  assign _zz_2580 = fixTo_68_dout;
  assign _zz_2581 = _zz_2582[35 : 0];
  assign _zz_2582 = _zz_2583;
  assign _zz_2583 = ($signed(_zz_2584) >>> _zz_59);
  assign _zz_2584 = _zz_2585;
  assign _zz_2585 = ($signed(_zz_2587) - $signed(_zz_57));
  assign _zz_2586 = ({9'd0,data_mid_0_22_imag} <<< 9);
  assign _zz_2587 = {{9{_zz_2586[26]}}, _zz_2586};
  assign _zz_2588 = fixTo_69_dout;
  assign _zz_2589 = _zz_2590[35 : 0];
  assign _zz_2590 = _zz_2591;
  assign _zz_2591 = ($signed(_zz_2592) >>> _zz_60);
  assign _zz_2592 = _zz_2593;
  assign _zz_2593 = ($signed(_zz_2595) + $signed(_zz_56));
  assign _zz_2594 = ({9'd0,data_mid_0_22_real} <<< 9);
  assign _zz_2595 = {{9{_zz_2594[26]}}, _zz_2594};
  assign _zz_2596 = fixTo_70_dout;
  assign _zz_2597 = _zz_2598[35 : 0];
  assign _zz_2598 = _zz_2599;
  assign _zz_2599 = ($signed(_zz_2600) >>> _zz_60);
  assign _zz_2600 = _zz_2601;
  assign _zz_2601 = ($signed(_zz_2603) + $signed(_zz_57));
  assign _zz_2602 = ({9'd0,data_mid_0_22_imag} <<< 9);
  assign _zz_2603 = {{9{_zz_2602[26]}}, _zz_2602};
  assign _zz_2604 = fixTo_71_dout;
  assign _zz_2605 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2606 = ($signed(_zz_63) - $signed(_zz_2607));
  assign _zz_2607 = ($signed(_zz_2608) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2608 = ($signed(data_mid_0_25_real) + $signed(data_mid_0_25_imag));
  assign _zz_2609 = fixTo_72_dout;
  assign _zz_2610 = ($signed(_zz_63) + $signed(_zz_2611));
  assign _zz_2611 = ($signed(_zz_2612) * $signed(twiddle_factor_table_0_real));
  assign _zz_2612 = ($signed(data_mid_0_25_imag) - $signed(data_mid_0_25_real));
  assign _zz_2613 = fixTo_73_dout;
  assign _zz_2614 = _zz_2615[35 : 0];
  assign _zz_2615 = _zz_2616;
  assign _zz_2616 = ($signed(_zz_2617) >>> _zz_64);
  assign _zz_2617 = _zz_2618;
  assign _zz_2618 = ($signed(_zz_2620) - $signed(_zz_61));
  assign _zz_2619 = ({9'd0,data_mid_0_24_real} <<< 9);
  assign _zz_2620 = {{9{_zz_2619[26]}}, _zz_2619};
  assign _zz_2621 = fixTo_74_dout;
  assign _zz_2622 = _zz_2623[35 : 0];
  assign _zz_2623 = _zz_2624;
  assign _zz_2624 = ($signed(_zz_2625) >>> _zz_64);
  assign _zz_2625 = _zz_2626;
  assign _zz_2626 = ($signed(_zz_2628) - $signed(_zz_62));
  assign _zz_2627 = ({9'd0,data_mid_0_24_imag} <<< 9);
  assign _zz_2628 = {{9{_zz_2627[26]}}, _zz_2627};
  assign _zz_2629 = fixTo_75_dout;
  assign _zz_2630 = _zz_2631[35 : 0];
  assign _zz_2631 = _zz_2632;
  assign _zz_2632 = ($signed(_zz_2633) >>> _zz_65);
  assign _zz_2633 = _zz_2634;
  assign _zz_2634 = ($signed(_zz_2636) + $signed(_zz_61));
  assign _zz_2635 = ({9'd0,data_mid_0_24_real} <<< 9);
  assign _zz_2636 = {{9{_zz_2635[26]}}, _zz_2635};
  assign _zz_2637 = fixTo_76_dout;
  assign _zz_2638 = _zz_2639[35 : 0];
  assign _zz_2639 = _zz_2640;
  assign _zz_2640 = ($signed(_zz_2641) >>> _zz_65);
  assign _zz_2641 = _zz_2642;
  assign _zz_2642 = ($signed(_zz_2644) + $signed(_zz_62));
  assign _zz_2643 = ({9'd0,data_mid_0_24_imag} <<< 9);
  assign _zz_2644 = {{9{_zz_2643[26]}}, _zz_2643};
  assign _zz_2645 = fixTo_77_dout;
  assign _zz_2646 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2647 = ($signed(_zz_68) - $signed(_zz_2648));
  assign _zz_2648 = ($signed(_zz_2649) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2649 = ($signed(data_mid_0_27_real) + $signed(data_mid_0_27_imag));
  assign _zz_2650 = fixTo_78_dout;
  assign _zz_2651 = ($signed(_zz_68) + $signed(_zz_2652));
  assign _zz_2652 = ($signed(_zz_2653) * $signed(twiddle_factor_table_0_real));
  assign _zz_2653 = ($signed(data_mid_0_27_imag) - $signed(data_mid_0_27_real));
  assign _zz_2654 = fixTo_79_dout;
  assign _zz_2655 = _zz_2656[35 : 0];
  assign _zz_2656 = _zz_2657;
  assign _zz_2657 = ($signed(_zz_2658) >>> _zz_69);
  assign _zz_2658 = _zz_2659;
  assign _zz_2659 = ($signed(_zz_2661) - $signed(_zz_66));
  assign _zz_2660 = ({9'd0,data_mid_0_26_real} <<< 9);
  assign _zz_2661 = {{9{_zz_2660[26]}}, _zz_2660};
  assign _zz_2662 = fixTo_80_dout;
  assign _zz_2663 = _zz_2664[35 : 0];
  assign _zz_2664 = _zz_2665;
  assign _zz_2665 = ($signed(_zz_2666) >>> _zz_69);
  assign _zz_2666 = _zz_2667;
  assign _zz_2667 = ($signed(_zz_2669) - $signed(_zz_67));
  assign _zz_2668 = ({9'd0,data_mid_0_26_imag} <<< 9);
  assign _zz_2669 = {{9{_zz_2668[26]}}, _zz_2668};
  assign _zz_2670 = fixTo_81_dout;
  assign _zz_2671 = _zz_2672[35 : 0];
  assign _zz_2672 = _zz_2673;
  assign _zz_2673 = ($signed(_zz_2674) >>> _zz_70);
  assign _zz_2674 = _zz_2675;
  assign _zz_2675 = ($signed(_zz_2677) + $signed(_zz_66));
  assign _zz_2676 = ({9'd0,data_mid_0_26_real} <<< 9);
  assign _zz_2677 = {{9{_zz_2676[26]}}, _zz_2676};
  assign _zz_2678 = fixTo_82_dout;
  assign _zz_2679 = _zz_2680[35 : 0];
  assign _zz_2680 = _zz_2681;
  assign _zz_2681 = ($signed(_zz_2682) >>> _zz_70);
  assign _zz_2682 = _zz_2683;
  assign _zz_2683 = ($signed(_zz_2685) + $signed(_zz_67));
  assign _zz_2684 = ({9'd0,data_mid_0_26_imag} <<< 9);
  assign _zz_2685 = {{9{_zz_2684[26]}}, _zz_2684};
  assign _zz_2686 = fixTo_83_dout;
  assign _zz_2687 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2688 = ($signed(_zz_73) - $signed(_zz_2689));
  assign _zz_2689 = ($signed(_zz_2690) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2690 = ($signed(data_mid_0_29_real) + $signed(data_mid_0_29_imag));
  assign _zz_2691 = fixTo_84_dout;
  assign _zz_2692 = ($signed(_zz_73) + $signed(_zz_2693));
  assign _zz_2693 = ($signed(_zz_2694) * $signed(twiddle_factor_table_0_real));
  assign _zz_2694 = ($signed(data_mid_0_29_imag) - $signed(data_mid_0_29_real));
  assign _zz_2695 = fixTo_85_dout;
  assign _zz_2696 = _zz_2697[35 : 0];
  assign _zz_2697 = _zz_2698;
  assign _zz_2698 = ($signed(_zz_2699) >>> _zz_74);
  assign _zz_2699 = _zz_2700;
  assign _zz_2700 = ($signed(_zz_2702) - $signed(_zz_71));
  assign _zz_2701 = ({9'd0,data_mid_0_28_real} <<< 9);
  assign _zz_2702 = {{9{_zz_2701[26]}}, _zz_2701};
  assign _zz_2703 = fixTo_86_dout;
  assign _zz_2704 = _zz_2705[35 : 0];
  assign _zz_2705 = _zz_2706;
  assign _zz_2706 = ($signed(_zz_2707) >>> _zz_74);
  assign _zz_2707 = _zz_2708;
  assign _zz_2708 = ($signed(_zz_2710) - $signed(_zz_72));
  assign _zz_2709 = ({9'd0,data_mid_0_28_imag} <<< 9);
  assign _zz_2710 = {{9{_zz_2709[26]}}, _zz_2709};
  assign _zz_2711 = fixTo_87_dout;
  assign _zz_2712 = _zz_2713[35 : 0];
  assign _zz_2713 = _zz_2714;
  assign _zz_2714 = ($signed(_zz_2715) >>> _zz_75);
  assign _zz_2715 = _zz_2716;
  assign _zz_2716 = ($signed(_zz_2718) + $signed(_zz_71));
  assign _zz_2717 = ({9'd0,data_mid_0_28_real} <<< 9);
  assign _zz_2718 = {{9{_zz_2717[26]}}, _zz_2717};
  assign _zz_2719 = fixTo_88_dout;
  assign _zz_2720 = _zz_2721[35 : 0];
  assign _zz_2721 = _zz_2722;
  assign _zz_2722 = ($signed(_zz_2723) >>> _zz_75);
  assign _zz_2723 = _zz_2724;
  assign _zz_2724 = ($signed(_zz_2726) + $signed(_zz_72));
  assign _zz_2725 = ({9'd0,data_mid_0_28_imag} <<< 9);
  assign _zz_2726 = {{9{_zz_2725[26]}}, _zz_2725};
  assign _zz_2727 = fixTo_89_dout;
  assign _zz_2728 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2729 = ($signed(_zz_78) - $signed(_zz_2730));
  assign _zz_2730 = ($signed(_zz_2731) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2731 = ($signed(data_mid_0_31_real) + $signed(data_mid_0_31_imag));
  assign _zz_2732 = fixTo_90_dout;
  assign _zz_2733 = ($signed(_zz_78) + $signed(_zz_2734));
  assign _zz_2734 = ($signed(_zz_2735) * $signed(twiddle_factor_table_0_real));
  assign _zz_2735 = ($signed(data_mid_0_31_imag) - $signed(data_mid_0_31_real));
  assign _zz_2736 = fixTo_91_dout;
  assign _zz_2737 = _zz_2738[35 : 0];
  assign _zz_2738 = _zz_2739;
  assign _zz_2739 = ($signed(_zz_2740) >>> _zz_79);
  assign _zz_2740 = _zz_2741;
  assign _zz_2741 = ($signed(_zz_2743) - $signed(_zz_76));
  assign _zz_2742 = ({9'd0,data_mid_0_30_real} <<< 9);
  assign _zz_2743 = {{9{_zz_2742[26]}}, _zz_2742};
  assign _zz_2744 = fixTo_92_dout;
  assign _zz_2745 = _zz_2746[35 : 0];
  assign _zz_2746 = _zz_2747;
  assign _zz_2747 = ($signed(_zz_2748) >>> _zz_79);
  assign _zz_2748 = _zz_2749;
  assign _zz_2749 = ($signed(_zz_2751) - $signed(_zz_77));
  assign _zz_2750 = ({9'd0,data_mid_0_30_imag} <<< 9);
  assign _zz_2751 = {{9{_zz_2750[26]}}, _zz_2750};
  assign _zz_2752 = fixTo_93_dout;
  assign _zz_2753 = _zz_2754[35 : 0];
  assign _zz_2754 = _zz_2755;
  assign _zz_2755 = ($signed(_zz_2756) >>> _zz_80);
  assign _zz_2756 = _zz_2757;
  assign _zz_2757 = ($signed(_zz_2759) + $signed(_zz_76));
  assign _zz_2758 = ({9'd0,data_mid_0_30_real} <<< 9);
  assign _zz_2759 = {{9{_zz_2758[26]}}, _zz_2758};
  assign _zz_2760 = fixTo_94_dout;
  assign _zz_2761 = _zz_2762[35 : 0];
  assign _zz_2762 = _zz_2763;
  assign _zz_2763 = ($signed(_zz_2764) >>> _zz_80);
  assign _zz_2764 = _zz_2765;
  assign _zz_2765 = ($signed(_zz_2767) + $signed(_zz_77));
  assign _zz_2766 = ({9'd0,data_mid_0_30_imag} <<< 9);
  assign _zz_2767 = {{9{_zz_2766[26]}}, _zz_2766};
  assign _zz_2768 = fixTo_95_dout;
  assign _zz_2769 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2770 = ($signed(_zz_83) - $signed(_zz_2771));
  assign _zz_2771 = ($signed(_zz_2772) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2772 = ($signed(data_mid_0_33_real) + $signed(data_mid_0_33_imag));
  assign _zz_2773 = fixTo_96_dout;
  assign _zz_2774 = ($signed(_zz_83) + $signed(_zz_2775));
  assign _zz_2775 = ($signed(_zz_2776) * $signed(twiddle_factor_table_0_real));
  assign _zz_2776 = ($signed(data_mid_0_33_imag) - $signed(data_mid_0_33_real));
  assign _zz_2777 = fixTo_97_dout;
  assign _zz_2778 = _zz_2779[35 : 0];
  assign _zz_2779 = _zz_2780;
  assign _zz_2780 = ($signed(_zz_2781) >>> _zz_84);
  assign _zz_2781 = _zz_2782;
  assign _zz_2782 = ($signed(_zz_2784) - $signed(_zz_81));
  assign _zz_2783 = ({9'd0,data_mid_0_32_real} <<< 9);
  assign _zz_2784 = {{9{_zz_2783[26]}}, _zz_2783};
  assign _zz_2785 = fixTo_98_dout;
  assign _zz_2786 = _zz_2787[35 : 0];
  assign _zz_2787 = _zz_2788;
  assign _zz_2788 = ($signed(_zz_2789) >>> _zz_84);
  assign _zz_2789 = _zz_2790;
  assign _zz_2790 = ($signed(_zz_2792) - $signed(_zz_82));
  assign _zz_2791 = ({9'd0,data_mid_0_32_imag} <<< 9);
  assign _zz_2792 = {{9{_zz_2791[26]}}, _zz_2791};
  assign _zz_2793 = fixTo_99_dout;
  assign _zz_2794 = _zz_2795[35 : 0];
  assign _zz_2795 = _zz_2796;
  assign _zz_2796 = ($signed(_zz_2797) >>> _zz_85);
  assign _zz_2797 = _zz_2798;
  assign _zz_2798 = ($signed(_zz_2800) + $signed(_zz_81));
  assign _zz_2799 = ({9'd0,data_mid_0_32_real} <<< 9);
  assign _zz_2800 = {{9{_zz_2799[26]}}, _zz_2799};
  assign _zz_2801 = fixTo_100_dout;
  assign _zz_2802 = _zz_2803[35 : 0];
  assign _zz_2803 = _zz_2804;
  assign _zz_2804 = ($signed(_zz_2805) >>> _zz_85);
  assign _zz_2805 = _zz_2806;
  assign _zz_2806 = ($signed(_zz_2808) + $signed(_zz_82));
  assign _zz_2807 = ({9'd0,data_mid_0_32_imag} <<< 9);
  assign _zz_2808 = {{9{_zz_2807[26]}}, _zz_2807};
  assign _zz_2809 = fixTo_101_dout;
  assign _zz_2810 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2811 = ($signed(_zz_88) - $signed(_zz_2812));
  assign _zz_2812 = ($signed(_zz_2813) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2813 = ($signed(data_mid_0_35_real) + $signed(data_mid_0_35_imag));
  assign _zz_2814 = fixTo_102_dout;
  assign _zz_2815 = ($signed(_zz_88) + $signed(_zz_2816));
  assign _zz_2816 = ($signed(_zz_2817) * $signed(twiddle_factor_table_0_real));
  assign _zz_2817 = ($signed(data_mid_0_35_imag) - $signed(data_mid_0_35_real));
  assign _zz_2818 = fixTo_103_dout;
  assign _zz_2819 = _zz_2820[35 : 0];
  assign _zz_2820 = _zz_2821;
  assign _zz_2821 = ($signed(_zz_2822) >>> _zz_89);
  assign _zz_2822 = _zz_2823;
  assign _zz_2823 = ($signed(_zz_2825) - $signed(_zz_86));
  assign _zz_2824 = ({9'd0,data_mid_0_34_real} <<< 9);
  assign _zz_2825 = {{9{_zz_2824[26]}}, _zz_2824};
  assign _zz_2826 = fixTo_104_dout;
  assign _zz_2827 = _zz_2828[35 : 0];
  assign _zz_2828 = _zz_2829;
  assign _zz_2829 = ($signed(_zz_2830) >>> _zz_89);
  assign _zz_2830 = _zz_2831;
  assign _zz_2831 = ($signed(_zz_2833) - $signed(_zz_87));
  assign _zz_2832 = ({9'd0,data_mid_0_34_imag} <<< 9);
  assign _zz_2833 = {{9{_zz_2832[26]}}, _zz_2832};
  assign _zz_2834 = fixTo_105_dout;
  assign _zz_2835 = _zz_2836[35 : 0];
  assign _zz_2836 = _zz_2837;
  assign _zz_2837 = ($signed(_zz_2838) >>> _zz_90);
  assign _zz_2838 = _zz_2839;
  assign _zz_2839 = ($signed(_zz_2841) + $signed(_zz_86));
  assign _zz_2840 = ({9'd0,data_mid_0_34_real} <<< 9);
  assign _zz_2841 = {{9{_zz_2840[26]}}, _zz_2840};
  assign _zz_2842 = fixTo_106_dout;
  assign _zz_2843 = _zz_2844[35 : 0];
  assign _zz_2844 = _zz_2845;
  assign _zz_2845 = ($signed(_zz_2846) >>> _zz_90);
  assign _zz_2846 = _zz_2847;
  assign _zz_2847 = ($signed(_zz_2849) + $signed(_zz_87));
  assign _zz_2848 = ({9'd0,data_mid_0_34_imag} <<< 9);
  assign _zz_2849 = {{9{_zz_2848[26]}}, _zz_2848};
  assign _zz_2850 = fixTo_107_dout;
  assign _zz_2851 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2852 = ($signed(_zz_93) - $signed(_zz_2853));
  assign _zz_2853 = ($signed(_zz_2854) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2854 = ($signed(data_mid_0_37_real) + $signed(data_mid_0_37_imag));
  assign _zz_2855 = fixTo_108_dout;
  assign _zz_2856 = ($signed(_zz_93) + $signed(_zz_2857));
  assign _zz_2857 = ($signed(_zz_2858) * $signed(twiddle_factor_table_0_real));
  assign _zz_2858 = ($signed(data_mid_0_37_imag) - $signed(data_mid_0_37_real));
  assign _zz_2859 = fixTo_109_dout;
  assign _zz_2860 = _zz_2861[35 : 0];
  assign _zz_2861 = _zz_2862;
  assign _zz_2862 = ($signed(_zz_2863) >>> _zz_94);
  assign _zz_2863 = _zz_2864;
  assign _zz_2864 = ($signed(_zz_2866) - $signed(_zz_91));
  assign _zz_2865 = ({9'd0,data_mid_0_36_real} <<< 9);
  assign _zz_2866 = {{9{_zz_2865[26]}}, _zz_2865};
  assign _zz_2867 = fixTo_110_dout;
  assign _zz_2868 = _zz_2869[35 : 0];
  assign _zz_2869 = _zz_2870;
  assign _zz_2870 = ($signed(_zz_2871) >>> _zz_94);
  assign _zz_2871 = _zz_2872;
  assign _zz_2872 = ($signed(_zz_2874) - $signed(_zz_92));
  assign _zz_2873 = ({9'd0,data_mid_0_36_imag} <<< 9);
  assign _zz_2874 = {{9{_zz_2873[26]}}, _zz_2873};
  assign _zz_2875 = fixTo_111_dout;
  assign _zz_2876 = _zz_2877[35 : 0];
  assign _zz_2877 = _zz_2878;
  assign _zz_2878 = ($signed(_zz_2879) >>> _zz_95);
  assign _zz_2879 = _zz_2880;
  assign _zz_2880 = ($signed(_zz_2882) + $signed(_zz_91));
  assign _zz_2881 = ({9'd0,data_mid_0_36_real} <<< 9);
  assign _zz_2882 = {{9{_zz_2881[26]}}, _zz_2881};
  assign _zz_2883 = fixTo_112_dout;
  assign _zz_2884 = _zz_2885[35 : 0];
  assign _zz_2885 = _zz_2886;
  assign _zz_2886 = ($signed(_zz_2887) >>> _zz_95);
  assign _zz_2887 = _zz_2888;
  assign _zz_2888 = ($signed(_zz_2890) + $signed(_zz_92));
  assign _zz_2889 = ({9'd0,data_mid_0_36_imag} <<< 9);
  assign _zz_2890 = {{9{_zz_2889[26]}}, _zz_2889};
  assign _zz_2891 = fixTo_113_dout;
  assign _zz_2892 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2893 = ($signed(_zz_98) - $signed(_zz_2894));
  assign _zz_2894 = ($signed(_zz_2895) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2895 = ($signed(data_mid_0_39_real) + $signed(data_mid_0_39_imag));
  assign _zz_2896 = fixTo_114_dout;
  assign _zz_2897 = ($signed(_zz_98) + $signed(_zz_2898));
  assign _zz_2898 = ($signed(_zz_2899) * $signed(twiddle_factor_table_0_real));
  assign _zz_2899 = ($signed(data_mid_0_39_imag) - $signed(data_mid_0_39_real));
  assign _zz_2900 = fixTo_115_dout;
  assign _zz_2901 = _zz_2902[35 : 0];
  assign _zz_2902 = _zz_2903;
  assign _zz_2903 = ($signed(_zz_2904) >>> _zz_99);
  assign _zz_2904 = _zz_2905;
  assign _zz_2905 = ($signed(_zz_2907) - $signed(_zz_96));
  assign _zz_2906 = ({9'd0,data_mid_0_38_real} <<< 9);
  assign _zz_2907 = {{9{_zz_2906[26]}}, _zz_2906};
  assign _zz_2908 = fixTo_116_dout;
  assign _zz_2909 = _zz_2910[35 : 0];
  assign _zz_2910 = _zz_2911;
  assign _zz_2911 = ($signed(_zz_2912) >>> _zz_99);
  assign _zz_2912 = _zz_2913;
  assign _zz_2913 = ($signed(_zz_2915) - $signed(_zz_97));
  assign _zz_2914 = ({9'd0,data_mid_0_38_imag} <<< 9);
  assign _zz_2915 = {{9{_zz_2914[26]}}, _zz_2914};
  assign _zz_2916 = fixTo_117_dout;
  assign _zz_2917 = _zz_2918[35 : 0];
  assign _zz_2918 = _zz_2919;
  assign _zz_2919 = ($signed(_zz_2920) >>> _zz_100);
  assign _zz_2920 = _zz_2921;
  assign _zz_2921 = ($signed(_zz_2923) + $signed(_zz_96));
  assign _zz_2922 = ({9'd0,data_mid_0_38_real} <<< 9);
  assign _zz_2923 = {{9{_zz_2922[26]}}, _zz_2922};
  assign _zz_2924 = fixTo_118_dout;
  assign _zz_2925 = _zz_2926[35 : 0];
  assign _zz_2926 = _zz_2927;
  assign _zz_2927 = ($signed(_zz_2928) >>> _zz_100);
  assign _zz_2928 = _zz_2929;
  assign _zz_2929 = ($signed(_zz_2931) + $signed(_zz_97));
  assign _zz_2930 = ({9'd0,data_mid_0_38_imag} <<< 9);
  assign _zz_2931 = {{9{_zz_2930[26]}}, _zz_2930};
  assign _zz_2932 = fixTo_119_dout;
  assign _zz_2933 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2934 = ($signed(_zz_103) - $signed(_zz_2935));
  assign _zz_2935 = ($signed(_zz_2936) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2936 = ($signed(data_mid_0_41_real) + $signed(data_mid_0_41_imag));
  assign _zz_2937 = fixTo_120_dout;
  assign _zz_2938 = ($signed(_zz_103) + $signed(_zz_2939));
  assign _zz_2939 = ($signed(_zz_2940) * $signed(twiddle_factor_table_0_real));
  assign _zz_2940 = ($signed(data_mid_0_41_imag) - $signed(data_mid_0_41_real));
  assign _zz_2941 = fixTo_121_dout;
  assign _zz_2942 = _zz_2943[35 : 0];
  assign _zz_2943 = _zz_2944;
  assign _zz_2944 = ($signed(_zz_2945) >>> _zz_104);
  assign _zz_2945 = _zz_2946;
  assign _zz_2946 = ($signed(_zz_2948) - $signed(_zz_101));
  assign _zz_2947 = ({9'd0,data_mid_0_40_real} <<< 9);
  assign _zz_2948 = {{9{_zz_2947[26]}}, _zz_2947};
  assign _zz_2949 = fixTo_122_dout;
  assign _zz_2950 = _zz_2951[35 : 0];
  assign _zz_2951 = _zz_2952;
  assign _zz_2952 = ($signed(_zz_2953) >>> _zz_104);
  assign _zz_2953 = _zz_2954;
  assign _zz_2954 = ($signed(_zz_2956) - $signed(_zz_102));
  assign _zz_2955 = ({9'd0,data_mid_0_40_imag} <<< 9);
  assign _zz_2956 = {{9{_zz_2955[26]}}, _zz_2955};
  assign _zz_2957 = fixTo_123_dout;
  assign _zz_2958 = _zz_2959[35 : 0];
  assign _zz_2959 = _zz_2960;
  assign _zz_2960 = ($signed(_zz_2961) >>> _zz_105);
  assign _zz_2961 = _zz_2962;
  assign _zz_2962 = ($signed(_zz_2964) + $signed(_zz_101));
  assign _zz_2963 = ({9'd0,data_mid_0_40_real} <<< 9);
  assign _zz_2964 = {{9{_zz_2963[26]}}, _zz_2963};
  assign _zz_2965 = fixTo_124_dout;
  assign _zz_2966 = _zz_2967[35 : 0];
  assign _zz_2967 = _zz_2968;
  assign _zz_2968 = ($signed(_zz_2969) >>> _zz_105);
  assign _zz_2969 = _zz_2970;
  assign _zz_2970 = ($signed(_zz_2972) + $signed(_zz_102));
  assign _zz_2971 = ({9'd0,data_mid_0_40_imag} <<< 9);
  assign _zz_2972 = {{9{_zz_2971[26]}}, _zz_2971};
  assign _zz_2973 = fixTo_125_dout;
  assign _zz_2974 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_2975 = ($signed(_zz_108) - $signed(_zz_2976));
  assign _zz_2976 = ($signed(_zz_2977) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2977 = ($signed(data_mid_0_43_real) + $signed(data_mid_0_43_imag));
  assign _zz_2978 = fixTo_126_dout;
  assign _zz_2979 = ($signed(_zz_108) + $signed(_zz_2980));
  assign _zz_2980 = ($signed(_zz_2981) * $signed(twiddle_factor_table_0_real));
  assign _zz_2981 = ($signed(data_mid_0_43_imag) - $signed(data_mid_0_43_real));
  assign _zz_2982 = fixTo_127_dout;
  assign _zz_2983 = _zz_2984[35 : 0];
  assign _zz_2984 = _zz_2985;
  assign _zz_2985 = ($signed(_zz_2986) >>> _zz_109);
  assign _zz_2986 = _zz_2987;
  assign _zz_2987 = ($signed(_zz_2989) - $signed(_zz_106));
  assign _zz_2988 = ({9'd0,data_mid_0_42_real} <<< 9);
  assign _zz_2989 = {{9{_zz_2988[26]}}, _zz_2988};
  assign _zz_2990 = fixTo_128_dout;
  assign _zz_2991 = _zz_2992[35 : 0];
  assign _zz_2992 = _zz_2993;
  assign _zz_2993 = ($signed(_zz_2994) >>> _zz_109);
  assign _zz_2994 = _zz_2995;
  assign _zz_2995 = ($signed(_zz_2997) - $signed(_zz_107));
  assign _zz_2996 = ({9'd0,data_mid_0_42_imag} <<< 9);
  assign _zz_2997 = {{9{_zz_2996[26]}}, _zz_2996};
  assign _zz_2998 = fixTo_129_dout;
  assign _zz_2999 = _zz_3000[35 : 0];
  assign _zz_3000 = _zz_3001;
  assign _zz_3001 = ($signed(_zz_3002) >>> _zz_110);
  assign _zz_3002 = _zz_3003;
  assign _zz_3003 = ($signed(_zz_3005) + $signed(_zz_106));
  assign _zz_3004 = ({9'd0,data_mid_0_42_real} <<< 9);
  assign _zz_3005 = {{9{_zz_3004[26]}}, _zz_3004};
  assign _zz_3006 = fixTo_130_dout;
  assign _zz_3007 = _zz_3008[35 : 0];
  assign _zz_3008 = _zz_3009;
  assign _zz_3009 = ($signed(_zz_3010) >>> _zz_110);
  assign _zz_3010 = _zz_3011;
  assign _zz_3011 = ($signed(_zz_3013) + $signed(_zz_107));
  assign _zz_3012 = ({9'd0,data_mid_0_42_imag} <<< 9);
  assign _zz_3013 = {{9{_zz_3012[26]}}, _zz_3012};
  assign _zz_3014 = fixTo_131_dout;
  assign _zz_3015 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_3016 = ($signed(_zz_113) - $signed(_zz_3017));
  assign _zz_3017 = ($signed(_zz_3018) * $signed(twiddle_factor_table_0_imag));
  assign _zz_3018 = ($signed(data_mid_0_45_real) + $signed(data_mid_0_45_imag));
  assign _zz_3019 = fixTo_132_dout;
  assign _zz_3020 = ($signed(_zz_113) + $signed(_zz_3021));
  assign _zz_3021 = ($signed(_zz_3022) * $signed(twiddle_factor_table_0_real));
  assign _zz_3022 = ($signed(data_mid_0_45_imag) - $signed(data_mid_0_45_real));
  assign _zz_3023 = fixTo_133_dout;
  assign _zz_3024 = _zz_3025[35 : 0];
  assign _zz_3025 = _zz_3026;
  assign _zz_3026 = ($signed(_zz_3027) >>> _zz_114);
  assign _zz_3027 = _zz_3028;
  assign _zz_3028 = ($signed(_zz_3030) - $signed(_zz_111));
  assign _zz_3029 = ({9'd0,data_mid_0_44_real} <<< 9);
  assign _zz_3030 = {{9{_zz_3029[26]}}, _zz_3029};
  assign _zz_3031 = fixTo_134_dout;
  assign _zz_3032 = _zz_3033[35 : 0];
  assign _zz_3033 = _zz_3034;
  assign _zz_3034 = ($signed(_zz_3035) >>> _zz_114);
  assign _zz_3035 = _zz_3036;
  assign _zz_3036 = ($signed(_zz_3038) - $signed(_zz_112));
  assign _zz_3037 = ({9'd0,data_mid_0_44_imag} <<< 9);
  assign _zz_3038 = {{9{_zz_3037[26]}}, _zz_3037};
  assign _zz_3039 = fixTo_135_dout;
  assign _zz_3040 = _zz_3041[35 : 0];
  assign _zz_3041 = _zz_3042;
  assign _zz_3042 = ($signed(_zz_3043) >>> _zz_115);
  assign _zz_3043 = _zz_3044;
  assign _zz_3044 = ($signed(_zz_3046) + $signed(_zz_111));
  assign _zz_3045 = ({9'd0,data_mid_0_44_real} <<< 9);
  assign _zz_3046 = {{9{_zz_3045[26]}}, _zz_3045};
  assign _zz_3047 = fixTo_136_dout;
  assign _zz_3048 = _zz_3049[35 : 0];
  assign _zz_3049 = _zz_3050;
  assign _zz_3050 = ($signed(_zz_3051) >>> _zz_115);
  assign _zz_3051 = _zz_3052;
  assign _zz_3052 = ($signed(_zz_3054) + $signed(_zz_112));
  assign _zz_3053 = ({9'd0,data_mid_0_44_imag} <<< 9);
  assign _zz_3054 = {{9{_zz_3053[26]}}, _zz_3053};
  assign _zz_3055 = fixTo_137_dout;
  assign _zz_3056 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_3057 = ($signed(_zz_118) - $signed(_zz_3058));
  assign _zz_3058 = ($signed(_zz_3059) * $signed(twiddle_factor_table_0_imag));
  assign _zz_3059 = ($signed(data_mid_0_47_real) + $signed(data_mid_0_47_imag));
  assign _zz_3060 = fixTo_138_dout;
  assign _zz_3061 = ($signed(_zz_118) + $signed(_zz_3062));
  assign _zz_3062 = ($signed(_zz_3063) * $signed(twiddle_factor_table_0_real));
  assign _zz_3063 = ($signed(data_mid_0_47_imag) - $signed(data_mid_0_47_real));
  assign _zz_3064 = fixTo_139_dout;
  assign _zz_3065 = _zz_3066[35 : 0];
  assign _zz_3066 = _zz_3067;
  assign _zz_3067 = ($signed(_zz_3068) >>> _zz_119);
  assign _zz_3068 = _zz_3069;
  assign _zz_3069 = ($signed(_zz_3071) - $signed(_zz_116));
  assign _zz_3070 = ({9'd0,data_mid_0_46_real} <<< 9);
  assign _zz_3071 = {{9{_zz_3070[26]}}, _zz_3070};
  assign _zz_3072 = fixTo_140_dout;
  assign _zz_3073 = _zz_3074[35 : 0];
  assign _zz_3074 = _zz_3075;
  assign _zz_3075 = ($signed(_zz_3076) >>> _zz_119);
  assign _zz_3076 = _zz_3077;
  assign _zz_3077 = ($signed(_zz_3079) - $signed(_zz_117));
  assign _zz_3078 = ({9'd0,data_mid_0_46_imag} <<< 9);
  assign _zz_3079 = {{9{_zz_3078[26]}}, _zz_3078};
  assign _zz_3080 = fixTo_141_dout;
  assign _zz_3081 = _zz_3082[35 : 0];
  assign _zz_3082 = _zz_3083;
  assign _zz_3083 = ($signed(_zz_3084) >>> _zz_120);
  assign _zz_3084 = _zz_3085;
  assign _zz_3085 = ($signed(_zz_3087) + $signed(_zz_116));
  assign _zz_3086 = ({9'd0,data_mid_0_46_real} <<< 9);
  assign _zz_3087 = {{9{_zz_3086[26]}}, _zz_3086};
  assign _zz_3088 = fixTo_142_dout;
  assign _zz_3089 = _zz_3090[35 : 0];
  assign _zz_3090 = _zz_3091;
  assign _zz_3091 = ($signed(_zz_3092) >>> _zz_120);
  assign _zz_3092 = _zz_3093;
  assign _zz_3093 = ($signed(_zz_3095) + $signed(_zz_117));
  assign _zz_3094 = ({9'd0,data_mid_0_46_imag} <<< 9);
  assign _zz_3095 = {{9{_zz_3094[26]}}, _zz_3094};
  assign _zz_3096 = fixTo_143_dout;
  assign _zz_3097 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_3098 = ($signed(_zz_123) - $signed(_zz_3099));
  assign _zz_3099 = ($signed(_zz_3100) * $signed(twiddle_factor_table_0_imag));
  assign _zz_3100 = ($signed(data_mid_0_49_real) + $signed(data_mid_0_49_imag));
  assign _zz_3101 = fixTo_144_dout;
  assign _zz_3102 = ($signed(_zz_123) + $signed(_zz_3103));
  assign _zz_3103 = ($signed(_zz_3104) * $signed(twiddle_factor_table_0_real));
  assign _zz_3104 = ($signed(data_mid_0_49_imag) - $signed(data_mid_0_49_real));
  assign _zz_3105 = fixTo_145_dout;
  assign _zz_3106 = _zz_3107[35 : 0];
  assign _zz_3107 = _zz_3108;
  assign _zz_3108 = ($signed(_zz_3109) >>> _zz_124);
  assign _zz_3109 = _zz_3110;
  assign _zz_3110 = ($signed(_zz_3112) - $signed(_zz_121));
  assign _zz_3111 = ({9'd0,data_mid_0_48_real} <<< 9);
  assign _zz_3112 = {{9{_zz_3111[26]}}, _zz_3111};
  assign _zz_3113 = fixTo_146_dout;
  assign _zz_3114 = _zz_3115[35 : 0];
  assign _zz_3115 = _zz_3116;
  assign _zz_3116 = ($signed(_zz_3117) >>> _zz_124);
  assign _zz_3117 = _zz_3118;
  assign _zz_3118 = ($signed(_zz_3120) - $signed(_zz_122));
  assign _zz_3119 = ({9'd0,data_mid_0_48_imag} <<< 9);
  assign _zz_3120 = {{9{_zz_3119[26]}}, _zz_3119};
  assign _zz_3121 = fixTo_147_dout;
  assign _zz_3122 = _zz_3123[35 : 0];
  assign _zz_3123 = _zz_3124;
  assign _zz_3124 = ($signed(_zz_3125) >>> _zz_125);
  assign _zz_3125 = _zz_3126;
  assign _zz_3126 = ($signed(_zz_3128) + $signed(_zz_121));
  assign _zz_3127 = ({9'd0,data_mid_0_48_real} <<< 9);
  assign _zz_3128 = {{9{_zz_3127[26]}}, _zz_3127};
  assign _zz_3129 = fixTo_148_dout;
  assign _zz_3130 = _zz_3131[35 : 0];
  assign _zz_3131 = _zz_3132;
  assign _zz_3132 = ($signed(_zz_3133) >>> _zz_125);
  assign _zz_3133 = _zz_3134;
  assign _zz_3134 = ($signed(_zz_3136) + $signed(_zz_122));
  assign _zz_3135 = ({9'd0,data_mid_0_48_imag} <<< 9);
  assign _zz_3136 = {{9{_zz_3135[26]}}, _zz_3135};
  assign _zz_3137 = fixTo_149_dout;
  assign _zz_3138 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_3139 = ($signed(_zz_128) - $signed(_zz_3140));
  assign _zz_3140 = ($signed(_zz_3141) * $signed(twiddle_factor_table_0_imag));
  assign _zz_3141 = ($signed(data_mid_0_51_real) + $signed(data_mid_0_51_imag));
  assign _zz_3142 = fixTo_150_dout;
  assign _zz_3143 = ($signed(_zz_128) + $signed(_zz_3144));
  assign _zz_3144 = ($signed(_zz_3145) * $signed(twiddle_factor_table_0_real));
  assign _zz_3145 = ($signed(data_mid_0_51_imag) - $signed(data_mid_0_51_real));
  assign _zz_3146 = fixTo_151_dout;
  assign _zz_3147 = _zz_3148[35 : 0];
  assign _zz_3148 = _zz_3149;
  assign _zz_3149 = ($signed(_zz_3150) >>> _zz_129);
  assign _zz_3150 = _zz_3151;
  assign _zz_3151 = ($signed(_zz_3153) - $signed(_zz_126));
  assign _zz_3152 = ({9'd0,data_mid_0_50_real} <<< 9);
  assign _zz_3153 = {{9{_zz_3152[26]}}, _zz_3152};
  assign _zz_3154 = fixTo_152_dout;
  assign _zz_3155 = _zz_3156[35 : 0];
  assign _zz_3156 = _zz_3157;
  assign _zz_3157 = ($signed(_zz_3158) >>> _zz_129);
  assign _zz_3158 = _zz_3159;
  assign _zz_3159 = ($signed(_zz_3161) - $signed(_zz_127));
  assign _zz_3160 = ({9'd0,data_mid_0_50_imag} <<< 9);
  assign _zz_3161 = {{9{_zz_3160[26]}}, _zz_3160};
  assign _zz_3162 = fixTo_153_dout;
  assign _zz_3163 = _zz_3164[35 : 0];
  assign _zz_3164 = _zz_3165;
  assign _zz_3165 = ($signed(_zz_3166) >>> _zz_130);
  assign _zz_3166 = _zz_3167;
  assign _zz_3167 = ($signed(_zz_3169) + $signed(_zz_126));
  assign _zz_3168 = ({9'd0,data_mid_0_50_real} <<< 9);
  assign _zz_3169 = {{9{_zz_3168[26]}}, _zz_3168};
  assign _zz_3170 = fixTo_154_dout;
  assign _zz_3171 = _zz_3172[35 : 0];
  assign _zz_3172 = _zz_3173;
  assign _zz_3173 = ($signed(_zz_3174) >>> _zz_130);
  assign _zz_3174 = _zz_3175;
  assign _zz_3175 = ($signed(_zz_3177) + $signed(_zz_127));
  assign _zz_3176 = ({9'd0,data_mid_0_50_imag} <<< 9);
  assign _zz_3177 = {{9{_zz_3176[26]}}, _zz_3176};
  assign _zz_3178 = fixTo_155_dout;
  assign _zz_3179 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_3180 = ($signed(_zz_133) - $signed(_zz_3181));
  assign _zz_3181 = ($signed(_zz_3182) * $signed(twiddle_factor_table_0_imag));
  assign _zz_3182 = ($signed(data_mid_0_53_real) + $signed(data_mid_0_53_imag));
  assign _zz_3183 = fixTo_156_dout;
  assign _zz_3184 = ($signed(_zz_133) + $signed(_zz_3185));
  assign _zz_3185 = ($signed(_zz_3186) * $signed(twiddle_factor_table_0_real));
  assign _zz_3186 = ($signed(data_mid_0_53_imag) - $signed(data_mid_0_53_real));
  assign _zz_3187 = fixTo_157_dout;
  assign _zz_3188 = _zz_3189[35 : 0];
  assign _zz_3189 = _zz_3190;
  assign _zz_3190 = ($signed(_zz_3191) >>> _zz_134);
  assign _zz_3191 = _zz_3192;
  assign _zz_3192 = ($signed(_zz_3194) - $signed(_zz_131));
  assign _zz_3193 = ({9'd0,data_mid_0_52_real} <<< 9);
  assign _zz_3194 = {{9{_zz_3193[26]}}, _zz_3193};
  assign _zz_3195 = fixTo_158_dout;
  assign _zz_3196 = _zz_3197[35 : 0];
  assign _zz_3197 = _zz_3198;
  assign _zz_3198 = ($signed(_zz_3199) >>> _zz_134);
  assign _zz_3199 = _zz_3200;
  assign _zz_3200 = ($signed(_zz_3202) - $signed(_zz_132));
  assign _zz_3201 = ({9'd0,data_mid_0_52_imag} <<< 9);
  assign _zz_3202 = {{9{_zz_3201[26]}}, _zz_3201};
  assign _zz_3203 = fixTo_159_dout;
  assign _zz_3204 = _zz_3205[35 : 0];
  assign _zz_3205 = _zz_3206;
  assign _zz_3206 = ($signed(_zz_3207) >>> _zz_135);
  assign _zz_3207 = _zz_3208;
  assign _zz_3208 = ($signed(_zz_3210) + $signed(_zz_131));
  assign _zz_3209 = ({9'd0,data_mid_0_52_real} <<< 9);
  assign _zz_3210 = {{9{_zz_3209[26]}}, _zz_3209};
  assign _zz_3211 = fixTo_160_dout;
  assign _zz_3212 = _zz_3213[35 : 0];
  assign _zz_3213 = _zz_3214;
  assign _zz_3214 = ($signed(_zz_3215) >>> _zz_135);
  assign _zz_3215 = _zz_3216;
  assign _zz_3216 = ($signed(_zz_3218) + $signed(_zz_132));
  assign _zz_3217 = ({9'd0,data_mid_0_52_imag} <<< 9);
  assign _zz_3218 = {{9{_zz_3217[26]}}, _zz_3217};
  assign _zz_3219 = fixTo_161_dout;
  assign _zz_3220 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_3221 = ($signed(_zz_138) - $signed(_zz_3222));
  assign _zz_3222 = ($signed(_zz_3223) * $signed(twiddle_factor_table_0_imag));
  assign _zz_3223 = ($signed(data_mid_0_55_real) + $signed(data_mid_0_55_imag));
  assign _zz_3224 = fixTo_162_dout;
  assign _zz_3225 = ($signed(_zz_138) + $signed(_zz_3226));
  assign _zz_3226 = ($signed(_zz_3227) * $signed(twiddle_factor_table_0_real));
  assign _zz_3227 = ($signed(data_mid_0_55_imag) - $signed(data_mid_0_55_real));
  assign _zz_3228 = fixTo_163_dout;
  assign _zz_3229 = _zz_3230[35 : 0];
  assign _zz_3230 = _zz_3231;
  assign _zz_3231 = ($signed(_zz_3232) >>> _zz_139);
  assign _zz_3232 = _zz_3233;
  assign _zz_3233 = ($signed(_zz_3235) - $signed(_zz_136));
  assign _zz_3234 = ({9'd0,data_mid_0_54_real} <<< 9);
  assign _zz_3235 = {{9{_zz_3234[26]}}, _zz_3234};
  assign _zz_3236 = fixTo_164_dout;
  assign _zz_3237 = _zz_3238[35 : 0];
  assign _zz_3238 = _zz_3239;
  assign _zz_3239 = ($signed(_zz_3240) >>> _zz_139);
  assign _zz_3240 = _zz_3241;
  assign _zz_3241 = ($signed(_zz_3243) - $signed(_zz_137));
  assign _zz_3242 = ({9'd0,data_mid_0_54_imag} <<< 9);
  assign _zz_3243 = {{9{_zz_3242[26]}}, _zz_3242};
  assign _zz_3244 = fixTo_165_dout;
  assign _zz_3245 = _zz_3246[35 : 0];
  assign _zz_3246 = _zz_3247;
  assign _zz_3247 = ($signed(_zz_3248) >>> _zz_140);
  assign _zz_3248 = _zz_3249;
  assign _zz_3249 = ($signed(_zz_3251) + $signed(_zz_136));
  assign _zz_3250 = ({9'd0,data_mid_0_54_real} <<< 9);
  assign _zz_3251 = {{9{_zz_3250[26]}}, _zz_3250};
  assign _zz_3252 = fixTo_166_dout;
  assign _zz_3253 = _zz_3254[35 : 0];
  assign _zz_3254 = _zz_3255;
  assign _zz_3255 = ($signed(_zz_3256) >>> _zz_140);
  assign _zz_3256 = _zz_3257;
  assign _zz_3257 = ($signed(_zz_3259) + $signed(_zz_137));
  assign _zz_3258 = ({9'd0,data_mid_0_54_imag} <<< 9);
  assign _zz_3259 = {{9{_zz_3258[26]}}, _zz_3258};
  assign _zz_3260 = fixTo_167_dout;
  assign _zz_3261 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_3262 = ($signed(_zz_143) - $signed(_zz_3263));
  assign _zz_3263 = ($signed(_zz_3264) * $signed(twiddle_factor_table_0_imag));
  assign _zz_3264 = ($signed(data_mid_0_57_real) + $signed(data_mid_0_57_imag));
  assign _zz_3265 = fixTo_168_dout;
  assign _zz_3266 = ($signed(_zz_143) + $signed(_zz_3267));
  assign _zz_3267 = ($signed(_zz_3268) * $signed(twiddle_factor_table_0_real));
  assign _zz_3268 = ($signed(data_mid_0_57_imag) - $signed(data_mid_0_57_real));
  assign _zz_3269 = fixTo_169_dout;
  assign _zz_3270 = _zz_3271[35 : 0];
  assign _zz_3271 = _zz_3272;
  assign _zz_3272 = ($signed(_zz_3273) >>> _zz_144);
  assign _zz_3273 = _zz_3274;
  assign _zz_3274 = ($signed(_zz_3276) - $signed(_zz_141));
  assign _zz_3275 = ({9'd0,data_mid_0_56_real} <<< 9);
  assign _zz_3276 = {{9{_zz_3275[26]}}, _zz_3275};
  assign _zz_3277 = fixTo_170_dout;
  assign _zz_3278 = _zz_3279[35 : 0];
  assign _zz_3279 = _zz_3280;
  assign _zz_3280 = ($signed(_zz_3281) >>> _zz_144);
  assign _zz_3281 = _zz_3282;
  assign _zz_3282 = ($signed(_zz_3284) - $signed(_zz_142));
  assign _zz_3283 = ({9'd0,data_mid_0_56_imag} <<< 9);
  assign _zz_3284 = {{9{_zz_3283[26]}}, _zz_3283};
  assign _zz_3285 = fixTo_171_dout;
  assign _zz_3286 = _zz_3287[35 : 0];
  assign _zz_3287 = _zz_3288;
  assign _zz_3288 = ($signed(_zz_3289) >>> _zz_145);
  assign _zz_3289 = _zz_3290;
  assign _zz_3290 = ($signed(_zz_3292) + $signed(_zz_141));
  assign _zz_3291 = ({9'd0,data_mid_0_56_real} <<< 9);
  assign _zz_3292 = {{9{_zz_3291[26]}}, _zz_3291};
  assign _zz_3293 = fixTo_172_dout;
  assign _zz_3294 = _zz_3295[35 : 0];
  assign _zz_3295 = _zz_3296;
  assign _zz_3296 = ($signed(_zz_3297) >>> _zz_145);
  assign _zz_3297 = _zz_3298;
  assign _zz_3298 = ($signed(_zz_3300) + $signed(_zz_142));
  assign _zz_3299 = ({9'd0,data_mid_0_56_imag} <<< 9);
  assign _zz_3300 = {{9{_zz_3299[26]}}, _zz_3299};
  assign _zz_3301 = fixTo_173_dout;
  assign _zz_3302 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_3303 = ($signed(_zz_148) - $signed(_zz_3304));
  assign _zz_3304 = ($signed(_zz_3305) * $signed(twiddle_factor_table_0_imag));
  assign _zz_3305 = ($signed(data_mid_0_59_real) + $signed(data_mid_0_59_imag));
  assign _zz_3306 = fixTo_174_dout;
  assign _zz_3307 = ($signed(_zz_148) + $signed(_zz_3308));
  assign _zz_3308 = ($signed(_zz_3309) * $signed(twiddle_factor_table_0_real));
  assign _zz_3309 = ($signed(data_mid_0_59_imag) - $signed(data_mid_0_59_real));
  assign _zz_3310 = fixTo_175_dout;
  assign _zz_3311 = _zz_3312[35 : 0];
  assign _zz_3312 = _zz_3313;
  assign _zz_3313 = ($signed(_zz_3314) >>> _zz_149);
  assign _zz_3314 = _zz_3315;
  assign _zz_3315 = ($signed(_zz_3317) - $signed(_zz_146));
  assign _zz_3316 = ({9'd0,data_mid_0_58_real} <<< 9);
  assign _zz_3317 = {{9{_zz_3316[26]}}, _zz_3316};
  assign _zz_3318 = fixTo_176_dout;
  assign _zz_3319 = _zz_3320[35 : 0];
  assign _zz_3320 = _zz_3321;
  assign _zz_3321 = ($signed(_zz_3322) >>> _zz_149);
  assign _zz_3322 = _zz_3323;
  assign _zz_3323 = ($signed(_zz_3325) - $signed(_zz_147));
  assign _zz_3324 = ({9'd0,data_mid_0_58_imag} <<< 9);
  assign _zz_3325 = {{9{_zz_3324[26]}}, _zz_3324};
  assign _zz_3326 = fixTo_177_dout;
  assign _zz_3327 = _zz_3328[35 : 0];
  assign _zz_3328 = _zz_3329;
  assign _zz_3329 = ($signed(_zz_3330) >>> _zz_150);
  assign _zz_3330 = _zz_3331;
  assign _zz_3331 = ($signed(_zz_3333) + $signed(_zz_146));
  assign _zz_3332 = ({9'd0,data_mid_0_58_real} <<< 9);
  assign _zz_3333 = {{9{_zz_3332[26]}}, _zz_3332};
  assign _zz_3334 = fixTo_178_dout;
  assign _zz_3335 = _zz_3336[35 : 0];
  assign _zz_3336 = _zz_3337;
  assign _zz_3337 = ($signed(_zz_3338) >>> _zz_150);
  assign _zz_3338 = _zz_3339;
  assign _zz_3339 = ($signed(_zz_3341) + $signed(_zz_147));
  assign _zz_3340 = ({9'd0,data_mid_0_58_imag} <<< 9);
  assign _zz_3341 = {{9{_zz_3340[26]}}, _zz_3340};
  assign _zz_3342 = fixTo_179_dout;
  assign _zz_3343 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_3344 = ($signed(_zz_153) - $signed(_zz_3345));
  assign _zz_3345 = ($signed(_zz_3346) * $signed(twiddle_factor_table_0_imag));
  assign _zz_3346 = ($signed(data_mid_0_61_real) + $signed(data_mid_0_61_imag));
  assign _zz_3347 = fixTo_180_dout;
  assign _zz_3348 = ($signed(_zz_153) + $signed(_zz_3349));
  assign _zz_3349 = ($signed(_zz_3350) * $signed(twiddle_factor_table_0_real));
  assign _zz_3350 = ($signed(data_mid_0_61_imag) - $signed(data_mid_0_61_real));
  assign _zz_3351 = fixTo_181_dout;
  assign _zz_3352 = _zz_3353[35 : 0];
  assign _zz_3353 = _zz_3354;
  assign _zz_3354 = ($signed(_zz_3355) >>> _zz_154);
  assign _zz_3355 = _zz_3356;
  assign _zz_3356 = ($signed(_zz_3358) - $signed(_zz_151));
  assign _zz_3357 = ({9'd0,data_mid_0_60_real} <<< 9);
  assign _zz_3358 = {{9{_zz_3357[26]}}, _zz_3357};
  assign _zz_3359 = fixTo_182_dout;
  assign _zz_3360 = _zz_3361[35 : 0];
  assign _zz_3361 = _zz_3362;
  assign _zz_3362 = ($signed(_zz_3363) >>> _zz_154);
  assign _zz_3363 = _zz_3364;
  assign _zz_3364 = ($signed(_zz_3366) - $signed(_zz_152));
  assign _zz_3365 = ({9'd0,data_mid_0_60_imag} <<< 9);
  assign _zz_3366 = {{9{_zz_3365[26]}}, _zz_3365};
  assign _zz_3367 = fixTo_183_dout;
  assign _zz_3368 = _zz_3369[35 : 0];
  assign _zz_3369 = _zz_3370;
  assign _zz_3370 = ($signed(_zz_3371) >>> _zz_155);
  assign _zz_3371 = _zz_3372;
  assign _zz_3372 = ($signed(_zz_3374) + $signed(_zz_151));
  assign _zz_3373 = ({9'd0,data_mid_0_60_real} <<< 9);
  assign _zz_3374 = {{9{_zz_3373[26]}}, _zz_3373};
  assign _zz_3375 = fixTo_184_dout;
  assign _zz_3376 = _zz_3377[35 : 0];
  assign _zz_3377 = _zz_3378;
  assign _zz_3378 = ($signed(_zz_3379) >>> _zz_155);
  assign _zz_3379 = _zz_3380;
  assign _zz_3380 = ($signed(_zz_3382) + $signed(_zz_152));
  assign _zz_3381 = ({9'd0,data_mid_0_60_imag} <<< 9);
  assign _zz_3382 = {{9{_zz_3381[26]}}, _zz_3381};
  assign _zz_3383 = fixTo_185_dout;
  assign _zz_3384 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_3385 = ($signed(_zz_158) - $signed(_zz_3386));
  assign _zz_3386 = ($signed(_zz_3387) * $signed(twiddle_factor_table_0_imag));
  assign _zz_3387 = ($signed(data_mid_0_63_real) + $signed(data_mid_0_63_imag));
  assign _zz_3388 = fixTo_186_dout;
  assign _zz_3389 = ($signed(_zz_158) + $signed(_zz_3390));
  assign _zz_3390 = ($signed(_zz_3391) * $signed(twiddle_factor_table_0_real));
  assign _zz_3391 = ($signed(data_mid_0_63_imag) - $signed(data_mid_0_63_real));
  assign _zz_3392 = fixTo_187_dout;
  assign _zz_3393 = _zz_3394[35 : 0];
  assign _zz_3394 = _zz_3395;
  assign _zz_3395 = ($signed(_zz_3396) >>> _zz_159);
  assign _zz_3396 = _zz_3397;
  assign _zz_3397 = ($signed(_zz_3399) - $signed(_zz_156));
  assign _zz_3398 = ({9'd0,data_mid_0_62_real} <<< 9);
  assign _zz_3399 = {{9{_zz_3398[26]}}, _zz_3398};
  assign _zz_3400 = fixTo_188_dout;
  assign _zz_3401 = _zz_3402[35 : 0];
  assign _zz_3402 = _zz_3403;
  assign _zz_3403 = ($signed(_zz_3404) >>> _zz_159);
  assign _zz_3404 = _zz_3405;
  assign _zz_3405 = ($signed(_zz_3407) - $signed(_zz_157));
  assign _zz_3406 = ({9'd0,data_mid_0_62_imag} <<< 9);
  assign _zz_3407 = {{9{_zz_3406[26]}}, _zz_3406};
  assign _zz_3408 = fixTo_189_dout;
  assign _zz_3409 = _zz_3410[35 : 0];
  assign _zz_3410 = _zz_3411;
  assign _zz_3411 = ($signed(_zz_3412) >>> _zz_160);
  assign _zz_3412 = _zz_3413;
  assign _zz_3413 = ($signed(_zz_3415) + $signed(_zz_156));
  assign _zz_3414 = ({9'd0,data_mid_0_62_real} <<< 9);
  assign _zz_3415 = {{9{_zz_3414[26]}}, _zz_3414};
  assign _zz_3416 = fixTo_190_dout;
  assign _zz_3417 = _zz_3418[35 : 0];
  assign _zz_3418 = _zz_3419;
  assign _zz_3419 = ($signed(_zz_3420) >>> _zz_160);
  assign _zz_3420 = _zz_3421;
  assign _zz_3421 = ($signed(_zz_3423) + $signed(_zz_157));
  assign _zz_3422 = ({9'd0,data_mid_0_62_imag} <<< 9);
  assign _zz_3423 = {{9{_zz_3422[26]}}, _zz_3422};
  assign _zz_3424 = fixTo_191_dout;
  assign _zz_3425 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_3426 = ($signed(_zz_163) - $signed(_zz_3427));
  assign _zz_3427 = ($signed(_zz_3428) * $signed(twiddle_factor_table_1_imag));
  assign _zz_3428 = ($signed(data_mid_1_2_real) + $signed(data_mid_1_2_imag));
  assign _zz_3429 = fixTo_192_dout;
  assign _zz_3430 = ($signed(_zz_163) + $signed(_zz_3431));
  assign _zz_3431 = ($signed(_zz_3432) * $signed(twiddle_factor_table_1_real));
  assign _zz_3432 = ($signed(data_mid_1_2_imag) - $signed(data_mid_1_2_real));
  assign _zz_3433 = fixTo_193_dout;
  assign _zz_3434 = _zz_3435[35 : 0];
  assign _zz_3435 = _zz_3436;
  assign _zz_3436 = ($signed(_zz_3437) >>> _zz_164);
  assign _zz_3437 = _zz_3438;
  assign _zz_3438 = ($signed(_zz_3440) - $signed(_zz_161));
  assign _zz_3439 = ({9'd0,data_mid_1_0_real} <<< 9);
  assign _zz_3440 = {{9{_zz_3439[26]}}, _zz_3439};
  assign _zz_3441 = fixTo_194_dout;
  assign _zz_3442 = _zz_3443[35 : 0];
  assign _zz_3443 = _zz_3444;
  assign _zz_3444 = ($signed(_zz_3445) >>> _zz_164);
  assign _zz_3445 = _zz_3446;
  assign _zz_3446 = ($signed(_zz_3448) - $signed(_zz_162));
  assign _zz_3447 = ({9'd0,data_mid_1_0_imag} <<< 9);
  assign _zz_3448 = {{9{_zz_3447[26]}}, _zz_3447};
  assign _zz_3449 = fixTo_195_dout;
  assign _zz_3450 = _zz_3451[35 : 0];
  assign _zz_3451 = _zz_3452;
  assign _zz_3452 = ($signed(_zz_3453) >>> _zz_165);
  assign _zz_3453 = _zz_3454;
  assign _zz_3454 = ($signed(_zz_3456) + $signed(_zz_161));
  assign _zz_3455 = ({9'd0,data_mid_1_0_real} <<< 9);
  assign _zz_3456 = {{9{_zz_3455[26]}}, _zz_3455};
  assign _zz_3457 = fixTo_196_dout;
  assign _zz_3458 = _zz_3459[35 : 0];
  assign _zz_3459 = _zz_3460;
  assign _zz_3460 = ($signed(_zz_3461) >>> _zz_165);
  assign _zz_3461 = _zz_3462;
  assign _zz_3462 = ($signed(_zz_3464) + $signed(_zz_162));
  assign _zz_3463 = ({9'd0,data_mid_1_0_imag} <<< 9);
  assign _zz_3464 = {{9{_zz_3463[26]}}, _zz_3463};
  assign _zz_3465 = fixTo_197_dout;
  assign _zz_3466 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_3467 = ($signed(_zz_168) - $signed(_zz_3468));
  assign _zz_3468 = ($signed(_zz_3469) * $signed(twiddle_factor_table_2_imag));
  assign _zz_3469 = ($signed(data_mid_1_3_real) + $signed(data_mid_1_3_imag));
  assign _zz_3470 = fixTo_198_dout;
  assign _zz_3471 = ($signed(_zz_168) + $signed(_zz_3472));
  assign _zz_3472 = ($signed(_zz_3473) * $signed(twiddle_factor_table_2_real));
  assign _zz_3473 = ($signed(data_mid_1_3_imag) - $signed(data_mid_1_3_real));
  assign _zz_3474 = fixTo_199_dout;
  assign _zz_3475 = _zz_3476[35 : 0];
  assign _zz_3476 = _zz_3477;
  assign _zz_3477 = ($signed(_zz_3478) >>> _zz_169);
  assign _zz_3478 = _zz_3479;
  assign _zz_3479 = ($signed(_zz_3481) - $signed(_zz_166));
  assign _zz_3480 = ({9'd0,data_mid_1_1_real} <<< 9);
  assign _zz_3481 = {{9{_zz_3480[26]}}, _zz_3480};
  assign _zz_3482 = fixTo_200_dout;
  assign _zz_3483 = _zz_3484[35 : 0];
  assign _zz_3484 = _zz_3485;
  assign _zz_3485 = ($signed(_zz_3486) >>> _zz_169);
  assign _zz_3486 = _zz_3487;
  assign _zz_3487 = ($signed(_zz_3489) - $signed(_zz_167));
  assign _zz_3488 = ({9'd0,data_mid_1_1_imag} <<< 9);
  assign _zz_3489 = {{9{_zz_3488[26]}}, _zz_3488};
  assign _zz_3490 = fixTo_201_dout;
  assign _zz_3491 = _zz_3492[35 : 0];
  assign _zz_3492 = _zz_3493;
  assign _zz_3493 = ($signed(_zz_3494) >>> _zz_170);
  assign _zz_3494 = _zz_3495;
  assign _zz_3495 = ($signed(_zz_3497) + $signed(_zz_166));
  assign _zz_3496 = ({9'd0,data_mid_1_1_real} <<< 9);
  assign _zz_3497 = {{9{_zz_3496[26]}}, _zz_3496};
  assign _zz_3498 = fixTo_202_dout;
  assign _zz_3499 = _zz_3500[35 : 0];
  assign _zz_3500 = _zz_3501;
  assign _zz_3501 = ($signed(_zz_3502) >>> _zz_170);
  assign _zz_3502 = _zz_3503;
  assign _zz_3503 = ($signed(_zz_3505) + $signed(_zz_167));
  assign _zz_3504 = ({9'd0,data_mid_1_1_imag} <<< 9);
  assign _zz_3505 = {{9{_zz_3504[26]}}, _zz_3504};
  assign _zz_3506 = fixTo_203_dout;
  assign _zz_3507 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_3508 = ($signed(_zz_173) - $signed(_zz_3509));
  assign _zz_3509 = ($signed(_zz_3510) * $signed(twiddle_factor_table_1_imag));
  assign _zz_3510 = ($signed(data_mid_1_6_real) + $signed(data_mid_1_6_imag));
  assign _zz_3511 = fixTo_204_dout;
  assign _zz_3512 = ($signed(_zz_173) + $signed(_zz_3513));
  assign _zz_3513 = ($signed(_zz_3514) * $signed(twiddle_factor_table_1_real));
  assign _zz_3514 = ($signed(data_mid_1_6_imag) - $signed(data_mid_1_6_real));
  assign _zz_3515 = fixTo_205_dout;
  assign _zz_3516 = _zz_3517[35 : 0];
  assign _zz_3517 = _zz_3518;
  assign _zz_3518 = ($signed(_zz_3519) >>> _zz_174);
  assign _zz_3519 = _zz_3520;
  assign _zz_3520 = ($signed(_zz_3522) - $signed(_zz_171));
  assign _zz_3521 = ({9'd0,data_mid_1_4_real} <<< 9);
  assign _zz_3522 = {{9{_zz_3521[26]}}, _zz_3521};
  assign _zz_3523 = fixTo_206_dout;
  assign _zz_3524 = _zz_3525[35 : 0];
  assign _zz_3525 = _zz_3526;
  assign _zz_3526 = ($signed(_zz_3527) >>> _zz_174);
  assign _zz_3527 = _zz_3528;
  assign _zz_3528 = ($signed(_zz_3530) - $signed(_zz_172));
  assign _zz_3529 = ({9'd0,data_mid_1_4_imag} <<< 9);
  assign _zz_3530 = {{9{_zz_3529[26]}}, _zz_3529};
  assign _zz_3531 = fixTo_207_dout;
  assign _zz_3532 = _zz_3533[35 : 0];
  assign _zz_3533 = _zz_3534;
  assign _zz_3534 = ($signed(_zz_3535) >>> _zz_175);
  assign _zz_3535 = _zz_3536;
  assign _zz_3536 = ($signed(_zz_3538) + $signed(_zz_171));
  assign _zz_3537 = ({9'd0,data_mid_1_4_real} <<< 9);
  assign _zz_3538 = {{9{_zz_3537[26]}}, _zz_3537};
  assign _zz_3539 = fixTo_208_dout;
  assign _zz_3540 = _zz_3541[35 : 0];
  assign _zz_3541 = _zz_3542;
  assign _zz_3542 = ($signed(_zz_3543) >>> _zz_175);
  assign _zz_3543 = _zz_3544;
  assign _zz_3544 = ($signed(_zz_3546) + $signed(_zz_172));
  assign _zz_3545 = ({9'd0,data_mid_1_4_imag} <<< 9);
  assign _zz_3546 = {{9{_zz_3545[26]}}, _zz_3545};
  assign _zz_3547 = fixTo_209_dout;
  assign _zz_3548 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_3549 = ($signed(_zz_178) - $signed(_zz_3550));
  assign _zz_3550 = ($signed(_zz_3551) * $signed(twiddle_factor_table_2_imag));
  assign _zz_3551 = ($signed(data_mid_1_7_real) + $signed(data_mid_1_7_imag));
  assign _zz_3552 = fixTo_210_dout;
  assign _zz_3553 = ($signed(_zz_178) + $signed(_zz_3554));
  assign _zz_3554 = ($signed(_zz_3555) * $signed(twiddle_factor_table_2_real));
  assign _zz_3555 = ($signed(data_mid_1_7_imag) - $signed(data_mid_1_7_real));
  assign _zz_3556 = fixTo_211_dout;
  assign _zz_3557 = _zz_3558[35 : 0];
  assign _zz_3558 = _zz_3559;
  assign _zz_3559 = ($signed(_zz_3560) >>> _zz_179);
  assign _zz_3560 = _zz_3561;
  assign _zz_3561 = ($signed(_zz_3563) - $signed(_zz_176));
  assign _zz_3562 = ({9'd0,data_mid_1_5_real} <<< 9);
  assign _zz_3563 = {{9{_zz_3562[26]}}, _zz_3562};
  assign _zz_3564 = fixTo_212_dout;
  assign _zz_3565 = _zz_3566[35 : 0];
  assign _zz_3566 = _zz_3567;
  assign _zz_3567 = ($signed(_zz_3568) >>> _zz_179);
  assign _zz_3568 = _zz_3569;
  assign _zz_3569 = ($signed(_zz_3571) - $signed(_zz_177));
  assign _zz_3570 = ({9'd0,data_mid_1_5_imag} <<< 9);
  assign _zz_3571 = {{9{_zz_3570[26]}}, _zz_3570};
  assign _zz_3572 = fixTo_213_dout;
  assign _zz_3573 = _zz_3574[35 : 0];
  assign _zz_3574 = _zz_3575;
  assign _zz_3575 = ($signed(_zz_3576) >>> _zz_180);
  assign _zz_3576 = _zz_3577;
  assign _zz_3577 = ($signed(_zz_3579) + $signed(_zz_176));
  assign _zz_3578 = ({9'd0,data_mid_1_5_real} <<< 9);
  assign _zz_3579 = {{9{_zz_3578[26]}}, _zz_3578};
  assign _zz_3580 = fixTo_214_dout;
  assign _zz_3581 = _zz_3582[35 : 0];
  assign _zz_3582 = _zz_3583;
  assign _zz_3583 = ($signed(_zz_3584) >>> _zz_180);
  assign _zz_3584 = _zz_3585;
  assign _zz_3585 = ($signed(_zz_3587) + $signed(_zz_177));
  assign _zz_3586 = ({9'd0,data_mid_1_5_imag} <<< 9);
  assign _zz_3587 = {{9{_zz_3586[26]}}, _zz_3586};
  assign _zz_3588 = fixTo_215_dout;
  assign _zz_3589 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_3590 = ($signed(_zz_183) - $signed(_zz_3591));
  assign _zz_3591 = ($signed(_zz_3592) * $signed(twiddle_factor_table_1_imag));
  assign _zz_3592 = ($signed(data_mid_1_10_real) + $signed(data_mid_1_10_imag));
  assign _zz_3593 = fixTo_216_dout;
  assign _zz_3594 = ($signed(_zz_183) + $signed(_zz_3595));
  assign _zz_3595 = ($signed(_zz_3596) * $signed(twiddle_factor_table_1_real));
  assign _zz_3596 = ($signed(data_mid_1_10_imag) - $signed(data_mid_1_10_real));
  assign _zz_3597 = fixTo_217_dout;
  assign _zz_3598 = _zz_3599[35 : 0];
  assign _zz_3599 = _zz_3600;
  assign _zz_3600 = ($signed(_zz_3601) >>> _zz_184);
  assign _zz_3601 = _zz_3602;
  assign _zz_3602 = ($signed(_zz_3604) - $signed(_zz_181));
  assign _zz_3603 = ({9'd0,data_mid_1_8_real} <<< 9);
  assign _zz_3604 = {{9{_zz_3603[26]}}, _zz_3603};
  assign _zz_3605 = fixTo_218_dout;
  assign _zz_3606 = _zz_3607[35 : 0];
  assign _zz_3607 = _zz_3608;
  assign _zz_3608 = ($signed(_zz_3609) >>> _zz_184);
  assign _zz_3609 = _zz_3610;
  assign _zz_3610 = ($signed(_zz_3612) - $signed(_zz_182));
  assign _zz_3611 = ({9'd0,data_mid_1_8_imag} <<< 9);
  assign _zz_3612 = {{9{_zz_3611[26]}}, _zz_3611};
  assign _zz_3613 = fixTo_219_dout;
  assign _zz_3614 = _zz_3615[35 : 0];
  assign _zz_3615 = _zz_3616;
  assign _zz_3616 = ($signed(_zz_3617) >>> _zz_185);
  assign _zz_3617 = _zz_3618;
  assign _zz_3618 = ($signed(_zz_3620) + $signed(_zz_181));
  assign _zz_3619 = ({9'd0,data_mid_1_8_real} <<< 9);
  assign _zz_3620 = {{9{_zz_3619[26]}}, _zz_3619};
  assign _zz_3621 = fixTo_220_dout;
  assign _zz_3622 = _zz_3623[35 : 0];
  assign _zz_3623 = _zz_3624;
  assign _zz_3624 = ($signed(_zz_3625) >>> _zz_185);
  assign _zz_3625 = _zz_3626;
  assign _zz_3626 = ($signed(_zz_3628) + $signed(_zz_182));
  assign _zz_3627 = ({9'd0,data_mid_1_8_imag} <<< 9);
  assign _zz_3628 = {{9{_zz_3627[26]}}, _zz_3627};
  assign _zz_3629 = fixTo_221_dout;
  assign _zz_3630 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_3631 = ($signed(_zz_188) - $signed(_zz_3632));
  assign _zz_3632 = ($signed(_zz_3633) * $signed(twiddle_factor_table_2_imag));
  assign _zz_3633 = ($signed(data_mid_1_11_real) + $signed(data_mid_1_11_imag));
  assign _zz_3634 = fixTo_222_dout;
  assign _zz_3635 = ($signed(_zz_188) + $signed(_zz_3636));
  assign _zz_3636 = ($signed(_zz_3637) * $signed(twiddle_factor_table_2_real));
  assign _zz_3637 = ($signed(data_mid_1_11_imag) - $signed(data_mid_1_11_real));
  assign _zz_3638 = fixTo_223_dout;
  assign _zz_3639 = _zz_3640[35 : 0];
  assign _zz_3640 = _zz_3641;
  assign _zz_3641 = ($signed(_zz_3642) >>> _zz_189);
  assign _zz_3642 = _zz_3643;
  assign _zz_3643 = ($signed(_zz_3645) - $signed(_zz_186));
  assign _zz_3644 = ({9'd0,data_mid_1_9_real} <<< 9);
  assign _zz_3645 = {{9{_zz_3644[26]}}, _zz_3644};
  assign _zz_3646 = fixTo_224_dout;
  assign _zz_3647 = _zz_3648[35 : 0];
  assign _zz_3648 = _zz_3649;
  assign _zz_3649 = ($signed(_zz_3650) >>> _zz_189);
  assign _zz_3650 = _zz_3651;
  assign _zz_3651 = ($signed(_zz_3653) - $signed(_zz_187));
  assign _zz_3652 = ({9'd0,data_mid_1_9_imag} <<< 9);
  assign _zz_3653 = {{9{_zz_3652[26]}}, _zz_3652};
  assign _zz_3654 = fixTo_225_dout;
  assign _zz_3655 = _zz_3656[35 : 0];
  assign _zz_3656 = _zz_3657;
  assign _zz_3657 = ($signed(_zz_3658) >>> _zz_190);
  assign _zz_3658 = _zz_3659;
  assign _zz_3659 = ($signed(_zz_3661) + $signed(_zz_186));
  assign _zz_3660 = ({9'd0,data_mid_1_9_real} <<< 9);
  assign _zz_3661 = {{9{_zz_3660[26]}}, _zz_3660};
  assign _zz_3662 = fixTo_226_dout;
  assign _zz_3663 = _zz_3664[35 : 0];
  assign _zz_3664 = _zz_3665;
  assign _zz_3665 = ($signed(_zz_3666) >>> _zz_190);
  assign _zz_3666 = _zz_3667;
  assign _zz_3667 = ($signed(_zz_3669) + $signed(_zz_187));
  assign _zz_3668 = ({9'd0,data_mid_1_9_imag} <<< 9);
  assign _zz_3669 = {{9{_zz_3668[26]}}, _zz_3668};
  assign _zz_3670 = fixTo_227_dout;
  assign _zz_3671 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_3672 = ($signed(_zz_193) - $signed(_zz_3673));
  assign _zz_3673 = ($signed(_zz_3674) * $signed(twiddle_factor_table_1_imag));
  assign _zz_3674 = ($signed(data_mid_1_14_real) + $signed(data_mid_1_14_imag));
  assign _zz_3675 = fixTo_228_dout;
  assign _zz_3676 = ($signed(_zz_193) + $signed(_zz_3677));
  assign _zz_3677 = ($signed(_zz_3678) * $signed(twiddle_factor_table_1_real));
  assign _zz_3678 = ($signed(data_mid_1_14_imag) - $signed(data_mid_1_14_real));
  assign _zz_3679 = fixTo_229_dout;
  assign _zz_3680 = _zz_3681[35 : 0];
  assign _zz_3681 = _zz_3682;
  assign _zz_3682 = ($signed(_zz_3683) >>> _zz_194);
  assign _zz_3683 = _zz_3684;
  assign _zz_3684 = ($signed(_zz_3686) - $signed(_zz_191));
  assign _zz_3685 = ({9'd0,data_mid_1_12_real} <<< 9);
  assign _zz_3686 = {{9{_zz_3685[26]}}, _zz_3685};
  assign _zz_3687 = fixTo_230_dout;
  assign _zz_3688 = _zz_3689[35 : 0];
  assign _zz_3689 = _zz_3690;
  assign _zz_3690 = ($signed(_zz_3691) >>> _zz_194);
  assign _zz_3691 = _zz_3692;
  assign _zz_3692 = ($signed(_zz_3694) - $signed(_zz_192));
  assign _zz_3693 = ({9'd0,data_mid_1_12_imag} <<< 9);
  assign _zz_3694 = {{9{_zz_3693[26]}}, _zz_3693};
  assign _zz_3695 = fixTo_231_dout;
  assign _zz_3696 = _zz_3697[35 : 0];
  assign _zz_3697 = _zz_3698;
  assign _zz_3698 = ($signed(_zz_3699) >>> _zz_195);
  assign _zz_3699 = _zz_3700;
  assign _zz_3700 = ($signed(_zz_3702) + $signed(_zz_191));
  assign _zz_3701 = ({9'd0,data_mid_1_12_real} <<< 9);
  assign _zz_3702 = {{9{_zz_3701[26]}}, _zz_3701};
  assign _zz_3703 = fixTo_232_dout;
  assign _zz_3704 = _zz_3705[35 : 0];
  assign _zz_3705 = _zz_3706;
  assign _zz_3706 = ($signed(_zz_3707) >>> _zz_195);
  assign _zz_3707 = _zz_3708;
  assign _zz_3708 = ($signed(_zz_3710) + $signed(_zz_192));
  assign _zz_3709 = ({9'd0,data_mid_1_12_imag} <<< 9);
  assign _zz_3710 = {{9{_zz_3709[26]}}, _zz_3709};
  assign _zz_3711 = fixTo_233_dout;
  assign _zz_3712 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_3713 = ($signed(_zz_198) - $signed(_zz_3714));
  assign _zz_3714 = ($signed(_zz_3715) * $signed(twiddle_factor_table_2_imag));
  assign _zz_3715 = ($signed(data_mid_1_15_real) + $signed(data_mid_1_15_imag));
  assign _zz_3716 = fixTo_234_dout;
  assign _zz_3717 = ($signed(_zz_198) + $signed(_zz_3718));
  assign _zz_3718 = ($signed(_zz_3719) * $signed(twiddle_factor_table_2_real));
  assign _zz_3719 = ($signed(data_mid_1_15_imag) - $signed(data_mid_1_15_real));
  assign _zz_3720 = fixTo_235_dout;
  assign _zz_3721 = _zz_3722[35 : 0];
  assign _zz_3722 = _zz_3723;
  assign _zz_3723 = ($signed(_zz_3724) >>> _zz_199);
  assign _zz_3724 = _zz_3725;
  assign _zz_3725 = ($signed(_zz_3727) - $signed(_zz_196));
  assign _zz_3726 = ({9'd0,data_mid_1_13_real} <<< 9);
  assign _zz_3727 = {{9{_zz_3726[26]}}, _zz_3726};
  assign _zz_3728 = fixTo_236_dout;
  assign _zz_3729 = _zz_3730[35 : 0];
  assign _zz_3730 = _zz_3731;
  assign _zz_3731 = ($signed(_zz_3732) >>> _zz_199);
  assign _zz_3732 = _zz_3733;
  assign _zz_3733 = ($signed(_zz_3735) - $signed(_zz_197));
  assign _zz_3734 = ({9'd0,data_mid_1_13_imag} <<< 9);
  assign _zz_3735 = {{9{_zz_3734[26]}}, _zz_3734};
  assign _zz_3736 = fixTo_237_dout;
  assign _zz_3737 = _zz_3738[35 : 0];
  assign _zz_3738 = _zz_3739;
  assign _zz_3739 = ($signed(_zz_3740) >>> _zz_200);
  assign _zz_3740 = _zz_3741;
  assign _zz_3741 = ($signed(_zz_3743) + $signed(_zz_196));
  assign _zz_3742 = ({9'd0,data_mid_1_13_real} <<< 9);
  assign _zz_3743 = {{9{_zz_3742[26]}}, _zz_3742};
  assign _zz_3744 = fixTo_238_dout;
  assign _zz_3745 = _zz_3746[35 : 0];
  assign _zz_3746 = _zz_3747;
  assign _zz_3747 = ($signed(_zz_3748) >>> _zz_200);
  assign _zz_3748 = _zz_3749;
  assign _zz_3749 = ($signed(_zz_3751) + $signed(_zz_197));
  assign _zz_3750 = ({9'd0,data_mid_1_13_imag} <<< 9);
  assign _zz_3751 = {{9{_zz_3750[26]}}, _zz_3750};
  assign _zz_3752 = fixTo_239_dout;
  assign _zz_3753 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_3754 = ($signed(_zz_203) - $signed(_zz_3755));
  assign _zz_3755 = ($signed(_zz_3756) * $signed(twiddle_factor_table_1_imag));
  assign _zz_3756 = ($signed(data_mid_1_18_real) + $signed(data_mid_1_18_imag));
  assign _zz_3757 = fixTo_240_dout;
  assign _zz_3758 = ($signed(_zz_203) + $signed(_zz_3759));
  assign _zz_3759 = ($signed(_zz_3760) * $signed(twiddle_factor_table_1_real));
  assign _zz_3760 = ($signed(data_mid_1_18_imag) - $signed(data_mid_1_18_real));
  assign _zz_3761 = fixTo_241_dout;
  assign _zz_3762 = _zz_3763[35 : 0];
  assign _zz_3763 = _zz_3764;
  assign _zz_3764 = ($signed(_zz_3765) >>> _zz_204);
  assign _zz_3765 = _zz_3766;
  assign _zz_3766 = ($signed(_zz_3768) - $signed(_zz_201));
  assign _zz_3767 = ({9'd0,data_mid_1_16_real} <<< 9);
  assign _zz_3768 = {{9{_zz_3767[26]}}, _zz_3767};
  assign _zz_3769 = fixTo_242_dout;
  assign _zz_3770 = _zz_3771[35 : 0];
  assign _zz_3771 = _zz_3772;
  assign _zz_3772 = ($signed(_zz_3773) >>> _zz_204);
  assign _zz_3773 = _zz_3774;
  assign _zz_3774 = ($signed(_zz_3776) - $signed(_zz_202));
  assign _zz_3775 = ({9'd0,data_mid_1_16_imag} <<< 9);
  assign _zz_3776 = {{9{_zz_3775[26]}}, _zz_3775};
  assign _zz_3777 = fixTo_243_dout;
  assign _zz_3778 = _zz_3779[35 : 0];
  assign _zz_3779 = _zz_3780;
  assign _zz_3780 = ($signed(_zz_3781) >>> _zz_205);
  assign _zz_3781 = _zz_3782;
  assign _zz_3782 = ($signed(_zz_3784) + $signed(_zz_201));
  assign _zz_3783 = ({9'd0,data_mid_1_16_real} <<< 9);
  assign _zz_3784 = {{9{_zz_3783[26]}}, _zz_3783};
  assign _zz_3785 = fixTo_244_dout;
  assign _zz_3786 = _zz_3787[35 : 0];
  assign _zz_3787 = _zz_3788;
  assign _zz_3788 = ($signed(_zz_3789) >>> _zz_205);
  assign _zz_3789 = _zz_3790;
  assign _zz_3790 = ($signed(_zz_3792) + $signed(_zz_202));
  assign _zz_3791 = ({9'd0,data_mid_1_16_imag} <<< 9);
  assign _zz_3792 = {{9{_zz_3791[26]}}, _zz_3791};
  assign _zz_3793 = fixTo_245_dout;
  assign _zz_3794 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_3795 = ($signed(_zz_208) - $signed(_zz_3796));
  assign _zz_3796 = ($signed(_zz_3797) * $signed(twiddle_factor_table_2_imag));
  assign _zz_3797 = ($signed(data_mid_1_19_real) + $signed(data_mid_1_19_imag));
  assign _zz_3798 = fixTo_246_dout;
  assign _zz_3799 = ($signed(_zz_208) + $signed(_zz_3800));
  assign _zz_3800 = ($signed(_zz_3801) * $signed(twiddle_factor_table_2_real));
  assign _zz_3801 = ($signed(data_mid_1_19_imag) - $signed(data_mid_1_19_real));
  assign _zz_3802 = fixTo_247_dout;
  assign _zz_3803 = _zz_3804[35 : 0];
  assign _zz_3804 = _zz_3805;
  assign _zz_3805 = ($signed(_zz_3806) >>> _zz_209);
  assign _zz_3806 = _zz_3807;
  assign _zz_3807 = ($signed(_zz_3809) - $signed(_zz_206));
  assign _zz_3808 = ({9'd0,data_mid_1_17_real} <<< 9);
  assign _zz_3809 = {{9{_zz_3808[26]}}, _zz_3808};
  assign _zz_3810 = fixTo_248_dout;
  assign _zz_3811 = _zz_3812[35 : 0];
  assign _zz_3812 = _zz_3813;
  assign _zz_3813 = ($signed(_zz_3814) >>> _zz_209);
  assign _zz_3814 = _zz_3815;
  assign _zz_3815 = ($signed(_zz_3817) - $signed(_zz_207));
  assign _zz_3816 = ({9'd0,data_mid_1_17_imag} <<< 9);
  assign _zz_3817 = {{9{_zz_3816[26]}}, _zz_3816};
  assign _zz_3818 = fixTo_249_dout;
  assign _zz_3819 = _zz_3820[35 : 0];
  assign _zz_3820 = _zz_3821;
  assign _zz_3821 = ($signed(_zz_3822) >>> _zz_210);
  assign _zz_3822 = _zz_3823;
  assign _zz_3823 = ($signed(_zz_3825) + $signed(_zz_206));
  assign _zz_3824 = ({9'd0,data_mid_1_17_real} <<< 9);
  assign _zz_3825 = {{9{_zz_3824[26]}}, _zz_3824};
  assign _zz_3826 = fixTo_250_dout;
  assign _zz_3827 = _zz_3828[35 : 0];
  assign _zz_3828 = _zz_3829;
  assign _zz_3829 = ($signed(_zz_3830) >>> _zz_210);
  assign _zz_3830 = _zz_3831;
  assign _zz_3831 = ($signed(_zz_3833) + $signed(_zz_207));
  assign _zz_3832 = ({9'd0,data_mid_1_17_imag} <<< 9);
  assign _zz_3833 = {{9{_zz_3832[26]}}, _zz_3832};
  assign _zz_3834 = fixTo_251_dout;
  assign _zz_3835 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_3836 = ($signed(_zz_213) - $signed(_zz_3837));
  assign _zz_3837 = ($signed(_zz_3838) * $signed(twiddle_factor_table_1_imag));
  assign _zz_3838 = ($signed(data_mid_1_22_real) + $signed(data_mid_1_22_imag));
  assign _zz_3839 = fixTo_252_dout;
  assign _zz_3840 = ($signed(_zz_213) + $signed(_zz_3841));
  assign _zz_3841 = ($signed(_zz_3842) * $signed(twiddle_factor_table_1_real));
  assign _zz_3842 = ($signed(data_mid_1_22_imag) - $signed(data_mid_1_22_real));
  assign _zz_3843 = fixTo_253_dout;
  assign _zz_3844 = _zz_3845[35 : 0];
  assign _zz_3845 = _zz_3846;
  assign _zz_3846 = ($signed(_zz_3847) >>> _zz_214);
  assign _zz_3847 = _zz_3848;
  assign _zz_3848 = ($signed(_zz_3850) - $signed(_zz_211));
  assign _zz_3849 = ({9'd0,data_mid_1_20_real} <<< 9);
  assign _zz_3850 = {{9{_zz_3849[26]}}, _zz_3849};
  assign _zz_3851 = fixTo_254_dout;
  assign _zz_3852 = _zz_3853[35 : 0];
  assign _zz_3853 = _zz_3854;
  assign _zz_3854 = ($signed(_zz_3855) >>> _zz_214);
  assign _zz_3855 = _zz_3856;
  assign _zz_3856 = ($signed(_zz_3858) - $signed(_zz_212));
  assign _zz_3857 = ({9'd0,data_mid_1_20_imag} <<< 9);
  assign _zz_3858 = {{9{_zz_3857[26]}}, _zz_3857};
  assign _zz_3859 = fixTo_255_dout;
  assign _zz_3860 = _zz_3861[35 : 0];
  assign _zz_3861 = _zz_3862;
  assign _zz_3862 = ($signed(_zz_3863) >>> _zz_215);
  assign _zz_3863 = _zz_3864;
  assign _zz_3864 = ($signed(_zz_3866) + $signed(_zz_211));
  assign _zz_3865 = ({9'd0,data_mid_1_20_real} <<< 9);
  assign _zz_3866 = {{9{_zz_3865[26]}}, _zz_3865};
  assign _zz_3867 = fixTo_256_dout;
  assign _zz_3868 = _zz_3869[35 : 0];
  assign _zz_3869 = _zz_3870;
  assign _zz_3870 = ($signed(_zz_3871) >>> _zz_215);
  assign _zz_3871 = _zz_3872;
  assign _zz_3872 = ($signed(_zz_3874) + $signed(_zz_212));
  assign _zz_3873 = ({9'd0,data_mid_1_20_imag} <<< 9);
  assign _zz_3874 = {{9{_zz_3873[26]}}, _zz_3873};
  assign _zz_3875 = fixTo_257_dout;
  assign _zz_3876 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_3877 = ($signed(_zz_218) - $signed(_zz_3878));
  assign _zz_3878 = ($signed(_zz_3879) * $signed(twiddle_factor_table_2_imag));
  assign _zz_3879 = ($signed(data_mid_1_23_real) + $signed(data_mid_1_23_imag));
  assign _zz_3880 = fixTo_258_dout;
  assign _zz_3881 = ($signed(_zz_218) + $signed(_zz_3882));
  assign _zz_3882 = ($signed(_zz_3883) * $signed(twiddle_factor_table_2_real));
  assign _zz_3883 = ($signed(data_mid_1_23_imag) - $signed(data_mid_1_23_real));
  assign _zz_3884 = fixTo_259_dout;
  assign _zz_3885 = _zz_3886[35 : 0];
  assign _zz_3886 = _zz_3887;
  assign _zz_3887 = ($signed(_zz_3888) >>> _zz_219);
  assign _zz_3888 = _zz_3889;
  assign _zz_3889 = ($signed(_zz_3891) - $signed(_zz_216));
  assign _zz_3890 = ({9'd0,data_mid_1_21_real} <<< 9);
  assign _zz_3891 = {{9{_zz_3890[26]}}, _zz_3890};
  assign _zz_3892 = fixTo_260_dout;
  assign _zz_3893 = _zz_3894[35 : 0];
  assign _zz_3894 = _zz_3895;
  assign _zz_3895 = ($signed(_zz_3896) >>> _zz_219);
  assign _zz_3896 = _zz_3897;
  assign _zz_3897 = ($signed(_zz_3899) - $signed(_zz_217));
  assign _zz_3898 = ({9'd0,data_mid_1_21_imag} <<< 9);
  assign _zz_3899 = {{9{_zz_3898[26]}}, _zz_3898};
  assign _zz_3900 = fixTo_261_dout;
  assign _zz_3901 = _zz_3902[35 : 0];
  assign _zz_3902 = _zz_3903;
  assign _zz_3903 = ($signed(_zz_3904) >>> _zz_220);
  assign _zz_3904 = _zz_3905;
  assign _zz_3905 = ($signed(_zz_3907) + $signed(_zz_216));
  assign _zz_3906 = ({9'd0,data_mid_1_21_real} <<< 9);
  assign _zz_3907 = {{9{_zz_3906[26]}}, _zz_3906};
  assign _zz_3908 = fixTo_262_dout;
  assign _zz_3909 = _zz_3910[35 : 0];
  assign _zz_3910 = _zz_3911;
  assign _zz_3911 = ($signed(_zz_3912) >>> _zz_220);
  assign _zz_3912 = _zz_3913;
  assign _zz_3913 = ($signed(_zz_3915) + $signed(_zz_217));
  assign _zz_3914 = ({9'd0,data_mid_1_21_imag} <<< 9);
  assign _zz_3915 = {{9{_zz_3914[26]}}, _zz_3914};
  assign _zz_3916 = fixTo_263_dout;
  assign _zz_3917 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_3918 = ($signed(_zz_223) - $signed(_zz_3919));
  assign _zz_3919 = ($signed(_zz_3920) * $signed(twiddle_factor_table_1_imag));
  assign _zz_3920 = ($signed(data_mid_1_26_real) + $signed(data_mid_1_26_imag));
  assign _zz_3921 = fixTo_264_dout;
  assign _zz_3922 = ($signed(_zz_223) + $signed(_zz_3923));
  assign _zz_3923 = ($signed(_zz_3924) * $signed(twiddle_factor_table_1_real));
  assign _zz_3924 = ($signed(data_mid_1_26_imag) - $signed(data_mid_1_26_real));
  assign _zz_3925 = fixTo_265_dout;
  assign _zz_3926 = _zz_3927[35 : 0];
  assign _zz_3927 = _zz_3928;
  assign _zz_3928 = ($signed(_zz_3929) >>> _zz_224);
  assign _zz_3929 = _zz_3930;
  assign _zz_3930 = ($signed(_zz_3932) - $signed(_zz_221));
  assign _zz_3931 = ({9'd0,data_mid_1_24_real} <<< 9);
  assign _zz_3932 = {{9{_zz_3931[26]}}, _zz_3931};
  assign _zz_3933 = fixTo_266_dout;
  assign _zz_3934 = _zz_3935[35 : 0];
  assign _zz_3935 = _zz_3936;
  assign _zz_3936 = ($signed(_zz_3937) >>> _zz_224);
  assign _zz_3937 = _zz_3938;
  assign _zz_3938 = ($signed(_zz_3940) - $signed(_zz_222));
  assign _zz_3939 = ({9'd0,data_mid_1_24_imag} <<< 9);
  assign _zz_3940 = {{9{_zz_3939[26]}}, _zz_3939};
  assign _zz_3941 = fixTo_267_dout;
  assign _zz_3942 = _zz_3943[35 : 0];
  assign _zz_3943 = _zz_3944;
  assign _zz_3944 = ($signed(_zz_3945) >>> _zz_225);
  assign _zz_3945 = _zz_3946;
  assign _zz_3946 = ($signed(_zz_3948) + $signed(_zz_221));
  assign _zz_3947 = ({9'd0,data_mid_1_24_real} <<< 9);
  assign _zz_3948 = {{9{_zz_3947[26]}}, _zz_3947};
  assign _zz_3949 = fixTo_268_dout;
  assign _zz_3950 = _zz_3951[35 : 0];
  assign _zz_3951 = _zz_3952;
  assign _zz_3952 = ($signed(_zz_3953) >>> _zz_225);
  assign _zz_3953 = _zz_3954;
  assign _zz_3954 = ($signed(_zz_3956) + $signed(_zz_222));
  assign _zz_3955 = ({9'd0,data_mid_1_24_imag} <<< 9);
  assign _zz_3956 = {{9{_zz_3955[26]}}, _zz_3955};
  assign _zz_3957 = fixTo_269_dout;
  assign _zz_3958 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_3959 = ($signed(_zz_228) - $signed(_zz_3960));
  assign _zz_3960 = ($signed(_zz_3961) * $signed(twiddle_factor_table_2_imag));
  assign _zz_3961 = ($signed(data_mid_1_27_real) + $signed(data_mid_1_27_imag));
  assign _zz_3962 = fixTo_270_dout;
  assign _zz_3963 = ($signed(_zz_228) + $signed(_zz_3964));
  assign _zz_3964 = ($signed(_zz_3965) * $signed(twiddle_factor_table_2_real));
  assign _zz_3965 = ($signed(data_mid_1_27_imag) - $signed(data_mid_1_27_real));
  assign _zz_3966 = fixTo_271_dout;
  assign _zz_3967 = _zz_3968[35 : 0];
  assign _zz_3968 = _zz_3969;
  assign _zz_3969 = ($signed(_zz_3970) >>> _zz_229);
  assign _zz_3970 = _zz_3971;
  assign _zz_3971 = ($signed(_zz_3973) - $signed(_zz_226));
  assign _zz_3972 = ({9'd0,data_mid_1_25_real} <<< 9);
  assign _zz_3973 = {{9{_zz_3972[26]}}, _zz_3972};
  assign _zz_3974 = fixTo_272_dout;
  assign _zz_3975 = _zz_3976[35 : 0];
  assign _zz_3976 = _zz_3977;
  assign _zz_3977 = ($signed(_zz_3978) >>> _zz_229);
  assign _zz_3978 = _zz_3979;
  assign _zz_3979 = ($signed(_zz_3981) - $signed(_zz_227));
  assign _zz_3980 = ({9'd0,data_mid_1_25_imag} <<< 9);
  assign _zz_3981 = {{9{_zz_3980[26]}}, _zz_3980};
  assign _zz_3982 = fixTo_273_dout;
  assign _zz_3983 = _zz_3984[35 : 0];
  assign _zz_3984 = _zz_3985;
  assign _zz_3985 = ($signed(_zz_3986) >>> _zz_230);
  assign _zz_3986 = _zz_3987;
  assign _zz_3987 = ($signed(_zz_3989) + $signed(_zz_226));
  assign _zz_3988 = ({9'd0,data_mid_1_25_real} <<< 9);
  assign _zz_3989 = {{9{_zz_3988[26]}}, _zz_3988};
  assign _zz_3990 = fixTo_274_dout;
  assign _zz_3991 = _zz_3992[35 : 0];
  assign _zz_3992 = _zz_3993;
  assign _zz_3993 = ($signed(_zz_3994) >>> _zz_230);
  assign _zz_3994 = _zz_3995;
  assign _zz_3995 = ($signed(_zz_3997) + $signed(_zz_227));
  assign _zz_3996 = ({9'd0,data_mid_1_25_imag} <<< 9);
  assign _zz_3997 = {{9{_zz_3996[26]}}, _zz_3996};
  assign _zz_3998 = fixTo_275_dout;
  assign _zz_3999 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_4000 = ($signed(_zz_233) - $signed(_zz_4001));
  assign _zz_4001 = ($signed(_zz_4002) * $signed(twiddle_factor_table_1_imag));
  assign _zz_4002 = ($signed(data_mid_1_30_real) + $signed(data_mid_1_30_imag));
  assign _zz_4003 = fixTo_276_dout;
  assign _zz_4004 = ($signed(_zz_233) + $signed(_zz_4005));
  assign _zz_4005 = ($signed(_zz_4006) * $signed(twiddle_factor_table_1_real));
  assign _zz_4006 = ($signed(data_mid_1_30_imag) - $signed(data_mid_1_30_real));
  assign _zz_4007 = fixTo_277_dout;
  assign _zz_4008 = _zz_4009[35 : 0];
  assign _zz_4009 = _zz_4010;
  assign _zz_4010 = ($signed(_zz_4011) >>> _zz_234);
  assign _zz_4011 = _zz_4012;
  assign _zz_4012 = ($signed(_zz_4014) - $signed(_zz_231));
  assign _zz_4013 = ({9'd0,data_mid_1_28_real} <<< 9);
  assign _zz_4014 = {{9{_zz_4013[26]}}, _zz_4013};
  assign _zz_4015 = fixTo_278_dout;
  assign _zz_4016 = _zz_4017[35 : 0];
  assign _zz_4017 = _zz_4018;
  assign _zz_4018 = ($signed(_zz_4019) >>> _zz_234);
  assign _zz_4019 = _zz_4020;
  assign _zz_4020 = ($signed(_zz_4022) - $signed(_zz_232));
  assign _zz_4021 = ({9'd0,data_mid_1_28_imag} <<< 9);
  assign _zz_4022 = {{9{_zz_4021[26]}}, _zz_4021};
  assign _zz_4023 = fixTo_279_dout;
  assign _zz_4024 = _zz_4025[35 : 0];
  assign _zz_4025 = _zz_4026;
  assign _zz_4026 = ($signed(_zz_4027) >>> _zz_235);
  assign _zz_4027 = _zz_4028;
  assign _zz_4028 = ($signed(_zz_4030) + $signed(_zz_231));
  assign _zz_4029 = ({9'd0,data_mid_1_28_real} <<< 9);
  assign _zz_4030 = {{9{_zz_4029[26]}}, _zz_4029};
  assign _zz_4031 = fixTo_280_dout;
  assign _zz_4032 = _zz_4033[35 : 0];
  assign _zz_4033 = _zz_4034;
  assign _zz_4034 = ($signed(_zz_4035) >>> _zz_235);
  assign _zz_4035 = _zz_4036;
  assign _zz_4036 = ($signed(_zz_4038) + $signed(_zz_232));
  assign _zz_4037 = ({9'd0,data_mid_1_28_imag} <<< 9);
  assign _zz_4038 = {{9{_zz_4037[26]}}, _zz_4037};
  assign _zz_4039 = fixTo_281_dout;
  assign _zz_4040 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_4041 = ($signed(_zz_238) - $signed(_zz_4042));
  assign _zz_4042 = ($signed(_zz_4043) * $signed(twiddle_factor_table_2_imag));
  assign _zz_4043 = ($signed(data_mid_1_31_real) + $signed(data_mid_1_31_imag));
  assign _zz_4044 = fixTo_282_dout;
  assign _zz_4045 = ($signed(_zz_238) + $signed(_zz_4046));
  assign _zz_4046 = ($signed(_zz_4047) * $signed(twiddle_factor_table_2_real));
  assign _zz_4047 = ($signed(data_mid_1_31_imag) - $signed(data_mid_1_31_real));
  assign _zz_4048 = fixTo_283_dout;
  assign _zz_4049 = _zz_4050[35 : 0];
  assign _zz_4050 = _zz_4051;
  assign _zz_4051 = ($signed(_zz_4052) >>> _zz_239);
  assign _zz_4052 = _zz_4053;
  assign _zz_4053 = ($signed(_zz_4055) - $signed(_zz_236));
  assign _zz_4054 = ({9'd0,data_mid_1_29_real} <<< 9);
  assign _zz_4055 = {{9{_zz_4054[26]}}, _zz_4054};
  assign _zz_4056 = fixTo_284_dout;
  assign _zz_4057 = _zz_4058[35 : 0];
  assign _zz_4058 = _zz_4059;
  assign _zz_4059 = ($signed(_zz_4060) >>> _zz_239);
  assign _zz_4060 = _zz_4061;
  assign _zz_4061 = ($signed(_zz_4063) - $signed(_zz_237));
  assign _zz_4062 = ({9'd0,data_mid_1_29_imag} <<< 9);
  assign _zz_4063 = {{9{_zz_4062[26]}}, _zz_4062};
  assign _zz_4064 = fixTo_285_dout;
  assign _zz_4065 = _zz_4066[35 : 0];
  assign _zz_4066 = _zz_4067;
  assign _zz_4067 = ($signed(_zz_4068) >>> _zz_240);
  assign _zz_4068 = _zz_4069;
  assign _zz_4069 = ($signed(_zz_4071) + $signed(_zz_236));
  assign _zz_4070 = ({9'd0,data_mid_1_29_real} <<< 9);
  assign _zz_4071 = {{9{_zz_4070[26]}}, _zz_4070};
  assign _zz_4072 = fixTo_286_dout;
  assign _zz_4073 = _zz_4074[35 : 0];
  assign _zz_4074 = _zz_4075;
  assign _zz_4075 = ($signed(_zz_4076) >>> _zz_240);
  assign _zz_4076 = _zz_4077;
  assign _zz_4077 = ($signed(_zz_4079) + $signed(_zz_237));
  assign _zz_4078 = ({9'd0,data_mid_1_29_imag} <<< 9);
  assign _zz_4079 = {{9{_zz_4078[26]}}, _zz_4078};
  assign _zz_4080 = fixTo_287_dout;
  assign _zz_4081 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_4082 = ($signed(_zz_243) - $signed(_zz_4083));
  assign _zz_4083 = ($signed(_zz_4084) * $signed(twiddle_factor_table_1_imag));
  assign _zz_4084 = ($signed(data_mid_1_34_real) + $signed(data_mid_1_34_imag));
  assign _zz_4085 = fixTo_288_dout;
  assign _zz_4086 = ($signed(_zz_243) + $signed(_zz_4087));
  assign _zz_4087 = ($signed(_zz_4088) * $signed(twiddle_factor_table_1_real));
  assign _zz_4088 = ($signed(data_mid_1_34_imag) - $signed(data_mid_1_34_real));
  assign _zz_4089 = fixTo_289_dout;
  assign _zz_4090 = _zz_4091[35 : 0];
  assign _zz_4091 = _zz_4092;
  assign _zz_4092 = ($signed(_zz_4093) >>> _zz_244);
  assign _zz_4093 = _zz_4094;
  assign _zz_4094 = ($signed(_zz_4096) - $signed(_zz_241));
  assign _zz_4095 = ({9'd0,data_mid_1_32_real} <<< 9);
  assign _zz_4096 = {{9{_zz_4095[26]}}, _zz_4095};
  assign _zz_4097 = fixTo_290_dout;
  assign _zz_4098 = _zz_4099[35 : 0];
  assign _zz_4099 = _zz_4100;
  assign _zz_4100 = ($signed(_zz_4101) >>> _zz_244);
  assign _zz_4101 = _zz_4102;
  assign _zz_4102 = ($signed(_zz_4104) - $signed(_zz_242));
  assign _zz_4103 = ({9'd0,data_mid_1_32_imag} <<< 9);
  assign _zz_4104 = {{9{_zz_4103[26]}}, _zz_4103};
  assign _zz_4105 = fixTo_291_dout;
  assign _zz_4106 = _zz_4107[35 : 0];
  assign _zz_4107 = _zz_4108;
  assign _zz_4108 = ($signed(_zz_4109) >>> _zz_245);
  assign _zz_4109 = _zz_4110;
  assign _zz_4110 = ($signed(_zz_4112) + $signed(_zz_241));
  assign _zz_4111 = ({9'd0,data_mid_1_32_real} <<< 9);
  assign _zz_4112 = {{9{_zz_4111[26]}}, _zz_4111};
  assign _zz_4113 = fixTo_292_dout;
  assign _zz_4114 = _zz_4115[35 : 0];
  assign _zz_4115 = _zz_4116;
  assign _zz_4116 = ($signed(_zz_4117) >>> _zz_245);
  assign _zz_4117 = _zz_4118;
  assign _zz_4118 = ($signed(_zz_4120) + $signed(_zz_242));
  assign _zz_4119 = ({9'd0,data_mid_1_32_imag} <<< 9);
  assign _zz_4120 = {{9{_zz_4119[26]}}, _zz_4119};
  assign _zz_4121 = fixTo_293_dout;
  assign _zz_4122 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_4123 = ($signed(_zz_248) - $signed(_zz_4124));
  assign _zz_4124 = ($signed(_zz_4125) * $signed(twiddle_factor_table_2_imag));
  assign _zz_4125 = ($signed(data_mid_1_35_real) + $signed(data_mid_1_35_imag));
  assign _zz_4126 = fixTo_294_dout;
  assign _zz_4127 = ($signed(_zz_248) + $signed(_zz_4128));
  assign _zz_4128 = ($signed(_zz_4129) * $signed(twiddle_factor_table_2_real));
  assign _zz_4129 = ($signed(data_mid_1_35_imag) - $signed(data_mid_1_35_real));
  assign _zz_4130 = fixTo_295_dout;
  assign _zz_4131 = _zz_4132[35 : 0];
  assign _zz_4132 = _zz_4133;
  assign _zz_4133 = ($signed(_zz_4134) >>> _zz_249);
  assign _zz_4134 = _zz_4135;
  assign _zz_4135 = ($signed(_zz_4137) - $signed(_zz_246));
  assign _zz_4136 = ({9'd0,data_mid_1_33_real} <<< 9);
  assign _zz_4137 = {{9{_zz_4136[26]}}, _zz_4136};
  assign _zz_4138 = fixTo_296_dout;
  assign _zz_4139 = _zz_4140[35 : 0];
  assign _zz_4140 = _zz_4141;
  assign _zz_4141 = ($signed(_zz_4142) >>> _zz_249);
  assign _zz_4142 = _zz_4143;
  assign _zz_4143 = ($signed(_zz_4145) - $signed(_zz_247));
  assign _zz_4144 = ({9'd0,data_mid_1_33_imag} <<< 9);
  assign _zz_4145 = {{9{_zz_4144[26]}}, _zz_4144};
  assign _zz_4146 = fixTo_297_dout;
  assign _zz_4147 = _zz_4148[35 : 0];
  assign _zz_4148 = _zz_4149;
  assign _zz_4149 = ($signed(_zz_4150) >>> _zz_250);
  assign _zz_4150 = _zz_4151;
  assign _zz_4151 = ($signed(_zz_4153) + $signed(_zz_246));
  assign _zz_4152 = ({9'd0,data_mid_1_33_real} <<< 9);
  assign _zz_4153 = {{9{_zz_4152[26]}}, _zz_4152};
  assign _zz_4154 = fixTo_298_dout;
  assign _zz_4155 = _zz_4156[35 : 0];
  assign _zz_4156 = _zz_4157;
  assign _zz_4157 = ($signed(_zz_4158) >>> _zz_250);
  assign _zz_4158 = _zz_4159;
  assign _zz_4159 = ($signed(_zz_4161) + $signed(_zz_247));
  assign _zz_4160 = ({9'd0,data_mid_1_33_imag} <<< 9);
  assign _zz_4161 = {{9{_zz_4160[26]}}, _zz_4160};
  assign _zz_4162 = fixTo_299_dout;
  assign _zz_4163 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_4164 = ($signed(_zz_253) - $signed(_zz_4165));
  assign _zz_4165 = ($signed(_zz_4166) * $signed(twiddle_factor_table_1_imag));
  assign _zz_4166 = ($signed(data_mid_1_38_real) + $signed(data_mid_1_38_imag));
  assign _zz_4167 = fixTo_300_dout;
  assign _zz_4168 = ($signed(_zz_253) + $signed(_zz_4169));
  assign _zz_4169 = ($signed(_zz_4170) * $signed(twiddle_factor_table_1_real));
  assign _zz_4170 = ($signed(data_mid_1_38_imag) - $signed(data_mid_1_38_real));
  assign _zz_4171 = fixTo_301_dout;
  assign _zz_4172 = _zz_4173[35 : 0];
  assign _zz_4173 = _zz_4174;
  assign _zz_4174 = ($signed(_zz_4175) >>> _zz_254);
  assign _zz_4175 = _zz_4176;
  assign _zz_4176 = ($signed(_zz_4178) - $signed(_zz_251));
  assign _zz_4177 = ({9'd0,data_mid_1_36_real} <<< 9);
  assign _zz_4178 = {{9{_zz_4177[26]}}, _zz_4177};
  assign _zz_4179 = fixTo_302_dout;
  assign _zz_4180 = _zz_4181[35 : 0];
  assign _zz_4181 = _zz_4182;
  assign _zz_4182 = ($signed(_zz_4183) >>> _zz_254);
  assign _zz_4183 = _zz_4184;
  assign _zz_4184 = ($signed(_zz_4186) - $signed(_zz_252));
  assign _zz_4185 = ({9'd0,data_mid_1_36_imag} <<< 9);
  assign _zz_4186 = {{9{_zz_4185[26]}}, _zz_4185};
  assign _zz_4187 = fixTo_303_dout;
  assign _zz_4188 = _zz_4189[35 : 0];
  assign _zz_4189 = _zz_4190;
  assign _zz_4190 = ($signed(_zz_4191) >>> _zz_255);
  assign _zz_4191 = _zz_4192;
  assign _zz_4192 = ($signed(_zz_4194) + $signed(_zz_251));
  assign _zz_4193 = ({9'd0,data_mid_1_36_real} <<< 9);
  assign _zz_4194 = {{9{_zz_4193[26]}}, _zz_4193};
  assign _zz_4195 = fixTo_304_dout;
  assign _zz_4196 = _zz_4197[35 : 0];
  assign _zz_4197 = _zz_4198;
  assign _zz_4198 = ($signed(_zz_4199) >>> _zz_255);
  assign _zz_4199 = _zz_4200;
  assign _zz_4200 = ($signed(_zz_4202) + $signed(_zz_252));
  assign _zz_4201 = ({9'd0,data_mid_1_36_imag} <<< 9);
  assign _zz_4202 = {{9{_zz_4201[26]}}, _zz_4201};
  assign _zz_4203 = fixTo_305_dout;
  assign _zz_4204 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_4205 = ($signed(_zz_258) - $signed(_zz_4206));
  assign _zz_4206 = ($signed(_zz_4207) * $signed(twiddle_factor_table_2_imag));
  assign _zz_4207 = ($signed(data_mid_1_39_real) + $signed(data_mid_1_39_imag));
  assign _zz_4208 = fixTo_306_dout;
  assign _zz_4209 = ($signed(_zz_258) + $signed(_zz_4210));
  assign _zz_4210 = ($signed(_zz_4211) * $signed(twiddle_factor_table_2_real));
  assign _zz_4211 = ($signed(data_mid_1_39_imag) - $signed(data_mid_1_39_real));
  assign _zz_4212 = fixTo_307_dout;
  assign _zz_4213 = _zz_4214[35 : 0];
  assign _zz_4214 = _zz_4215;
  assign _zz_4215 = ($signed(_zz_4216) >>> _zz_259);
  assign _zz_4216 = _zz_4217;
  assign _zz_4217 = ($signed(_zz_4219) - $signed(_zz_256));
  assign _zz_4218 = ({9'd0,data_mid_1_37_real} <<< 9);
  assign _zz_4219 = {{9{_zz_4218[26]}}, _zz_4218};
  assign _zz_4220 = fixTo_308_dout;
  assign _zz_4221 = _zz_4222[35 : 0];
  assign _zz_4222 = _zz_4223;
  assign _zz_4223 = ($signed(_zz_4224) >>> _zz_259);
  assign _zz_4224 = _zz_4225;
  assign _zz_4225 = ($signed(_zz_4227) - $signed(_zz_257));
  assign _zz_4226 = ({9'd0,data_mid_1_37_imag} <<< 9);
  assign _zz_4227 = {{9{_zz_4226[26]}}, _zz_4226};
  assign _zz_4228 = fixTo_309_dout;
  assign _zz_4229 = _zz_4230[35 : 0];
  assign _zz_4230 = _zz_4231;
  assign _zz_4231 = ($signed(_zz_4232) >>> _zz_260);
  assign _zz_4232 = _zz_4233;
  assign _zz_4233 = ($signed(_zz_4235) + $signed(_zz_256));
  assign _zz_4234 = ({9'd0,data_mid_1_37_real} <<< 9);
  assign _zz_4235 = {{9{_zz_4234[26]}}, _zz_4234};
  assign _zz_4236 = fixTo_310_dout;
  assign _zz_4237 = _zz_4238[35 : 0];
  assign _zz_4238 = _zz_4239;
  assign _zz_4239 = ($signed(_zz_4240) >>> _zz_260);
  assign _zz_4240 = _zz_4241;
  assign _zz_4241 = ($signed(_zz_4243) + $signed(_zz_257));
  assign _zz_4242 = ({9'd0,data_mid_1_37_imag} <<< 9);
  assign _zz_4243 = {{9{_zz_4242[26]}}, _zz_4242};
  assign _zz_4244 = fixTo_311_dout;
  assign _zz_4245 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_4246 = ($signed(_zz_263) - $signed(_zz_4247));
  assign _zz_4247 = ($signed(_zz_4248) * $signed(twiddle_factor_table_1_imag));
  assign _zz_4248 = ($signed(data_mid_1_42_real) + $signed(data_mid_1_42_imag));
  assign _zz_4249 = fixTo_312_dout;
  assign _zz_4250 = ($signed(_zz_263) + $signed(_zz_4251));
  assign _zz_4251 = ($signed(_zz_4252) * $signed(twiddle_factor_table_1_real));
  assign _zz_4252 = ($signed(data_mid_1_42_imag) - $signed(data_mid_1_42_real));
  assign _zz_4253 = fixTo_313_dout;
  assign _zz_4254 = _zz_4255[35 : 0];
  assign _zz_4255 = _zz_4256;
  assign _zz_4256 = ($signed(_zz_4257) >>> _zz_264);
  assign _zz_4257 = _zz_4258;
  assign _zz_4258 = ($signed(_zz_4260) - $signed(_zz_261));
  assign _zz_4259 = ({9'd0,data_mid_1_40_real} <<< 9);
  assign _zz_4260 = {{9{_zz_4259[26]}}, _zz_4259};
  assign _zz_4261 = fixTo_314_dout;
  assign _zz_4262 = _zz_4263[35 : 0];
  assign _zz_4263 = _zz_4264;
  assign _zz_4264 = ($signed(_zz_4265) >>> _zz_264);
  assign _zz_4265 = _zz_4266;
  assign _zz_4266 = ($signed(_zz_4268) - $signed(_zz_262));
  assign _zz_4267 = ({9'd0,data_mid_1_40_imag} <<< 9);
  assign _zz_4268 = {{9{_zz_4267[26]}}, _zz_4267};
  assign _zz_4269 = fixTo_315_dout;
  assign _zz_4270 = _zz_4271[35 : 0];
  assign _zz_4271 = _zz_4272;
  assign _zz_4272 = ($signed(_zz_4273) >>> _zz_265);
  assign _zz_4273 = _zz_4274;
  assign _zz_4274 = ($signed(_zz_4276) + $signed(_zz_261));
  assign _zz_4275 = ({9'd0,data_mid_1_40_real} <<< 9);
  assign _zz_4276 = {{9{_zz_4275[26]}}, _zz_4275};
  assign _zz_4277 = fixTo_316_dout;
  assign _zz_4278 = _zz_4279[35 : 0];
  assign _zz_4279 = _zz_4280;
  assign _zz_4280 = ($signed(_zz_4281) >>> _zz_265);
  assign _zz_4281 = _zz_4282;
  assign _zz_4282 = ($signed(_zz_4284) + $signed(_zz_262));
  assign _zz_4283 = ({9'd0,data_mid_1_40_imag} <<< 9);
  assign _zz_4284 = {{9{_zz_4283[26]}}, _zz_4283};
  assign _zz_4285 = fixTo_317_dout;
  assign _zz_4286 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_4287 = ($signed(_zz_268) - $signed(_zz_4288));
  assign _zz_4288 = ($signed(_zz_4289) * $signed(twiddle_factor_table_2_imag));
  assign _zz_4289 = ($signed(data_mid_1_43_real) + $signed(data_mid_1_43_imag));
  assign _zz_4290 = fixTo_318_dout;
  assign _zz_4291 = ($signed(_zz_268) + $signed(_zz_4292));
  assign _zz_4292 = ($signed(_zz_4293) * $signed(twiddle_factor_table_2_real));
  assign _zz_4293 = ($signed(data_mid_1_43_imag) - $signed(data_mid_1_43_real));
  assign _zz_4294 = fixTo_319_dout;
  assign _zz_4295 = _zz_4296[35 : 0];
  assign _zz_4296 = _zz_4297;
  assign _zz_4297 = ($signed(_zz_4298) >>> _zz_269);
  assign _zz_4298 = _zz_4299;
  assign _zz_4299 = ($signed(_zz_4301) - $signed(_zz_266));
  assign _zz_4300 = ({9'd0,data_mid_1_41_real} <<< 9);
  assign _zz_4301 = {{9{_zz_4300[26]}}, _zz_4300};
  assign _zz_4302 = fixTo_320_dout;
  assign _zz_4303 = _zz_4304[35 : 0];
  assign _zz_4304 = _zz_4305;
  assign _zz_4305 = ($signed(_zz_4306) >>> _zz_269);
  assign _zz_4306 = _zz_4307;
  assign _zz_4307 = ($signed(_zz_4309) - $signed(_zz_267));
  assign _zz_4308 = ({9'd0,data_mid_1_41_imag} <<< 9);
  assign _zz_4309 = {{9{_zz_4308[26]}}, _zz_4308};
  assign _zz_4310 = fixTo_321_dout;
  assign _zz_4311 = _zz_4312[35 : 0];
  assign _zz_4312 = _zz_4313;
  assign _zz_4313 = ($signed(_zz_4314) >>> _zz_270);
  assign _zz_4314 = _zz_4315;
  assign _zz_4315 = ($signed(_zz_4317) + $signed(_zz_266));
  assign _zz_4316 = ({9'd0,data_mid_1_41_real} <<< 9);
  assign _zz_4317 = {{9{_zz_4316[26]}}, _zz_4316};
  assign _zz_4318 = fixTo_322_dout;
  assign _zz_4319 = _zz_4320[35 : 0];
  assign _zz_4320 = _zz_4321;
  assign _zz_4321 = ($signed(_zz_4322) >>> _zz_270);
  assign _zz_4322 = _zz_4323;
  assign _zz_4323 = ($signed(_zz_4325) + $signed(_zz_267));
  assign _zz_4324 = ({9'd0,data_mid_1_41_imag} <<< 9);
  assign _zz_4325 = {{9{_zz_4324[26]}}, _zz_4324};
  assign _zz_4326 = fixTo_323_dout;
  assign _zz_4327 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_4328 = ($signed(_zz_273) - $signed(_zz_4329));
  assign _zz_4329 = ($signed(_zz_4330) * $signed(twiddle_factor_table_1_imag));
  assign _zz_4330 = ($signed(data_mid_1_46_real) + $signed(data_mid_1_46_imag));
  assign _zz_4331 = fixTo_324_dout;
  assign _zz_4332 = ($signed(_zz_273) + $signed(_zz_4333));
  assign _zz_4333 = ($signed(_zz_4334) * $signed(twiddle_factor_table_1_real));
  assign _zz_4334 = ($signed(data_mid_1_46_imag) - $signed(data_mid_1_46_real));
  assign _zz_4335 = fixTo_325_dout;
  assign _zz_4336 = _zz_4337[35 : 0];
  assign _zz_4337 = _zz_4338;
  assign _zz_4338 = ($signed(_zz_4339) >>> _zz_274);
  assign _zz_4339 = _zz_4340;
  assign _zz_4340 = ($signed(_zz_4342) - $signed(_zz_271));
  assign _zz_4341 = ({9'd0,data_mid_1_44_real} <<< 9);
  assign _zz_4342 = {{9{_zz_4341[26]}}, _zz_4341};
  assign _zz_4343 = fixTo_326_dout;
  assign _zz_4344 = _zz_4345[35 : 0];
  assign _zz_4345 = _zz_4346;
  assign _zz_4346 = ($signed(_zz_4347) >>> _zz_274);
  assign _zz_4347 = _zz_4348;
  assign _zz_4348 = ($signed(_zz_4350) - $signed(_zz_272));
  assign _zz_4349 = ({9'd0,data_mid_1_44_imag} <<< 9);
  assign _zz_4350 = {{9{_zz_4349[26]}}, _zz_4349};
  assign _zz_4351 = fixTo_327_dout;
  assign _zz_4352 = _zz_4353[35 : 0];
  assign _zz_4353 = _zz_4354;
  assign _zz_4354 = ($signed(_zz_4355) >>> _zz_275);
  assign _zz_4355 = _zz_4356;
  assign _zz_4356 = ($signed(_zz_4358) + $signed(_zz_271));
  assign _zz_4357 = ({9'd0,data_mid_1_44_real} <<< 9);
  assign _zz_4358 = {{9{_zz_4357[26]}}, _zz_4357};
  assign _zz_4359 = fixTo_328_dout;
  assign _zz_4360 = _zz_4361[35 : 0];
  assign _zz_4361 = _zz_4362;
  assign _zz_4362 = ($signed(_zz_4363) >>> _zz_275);
  assign _zz_4363 = _zz_4364;
  assign _zz_4364 = ($signed(_zz_4366) + $signed(_zz_272));
  assign _zz_4365 = ({9'd0,data_mid_1_44_imag} <<< 9);
  assign _zz_4366 = {{9{_zz_4365[26]}}, _zz_4365};
  assign _zz_4367 = fixTo_329_dout;
  assign _zz_4368 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_4369 = ($signed(_zz_278) - $signed(_zz_4370));
  assign _zz_4370 = ($signed(_zz_4371) * $signed(twiddle_factor_table_2_imag));
  assign _zz_4371 = ($signed(data_mid_1_47_real) + $signed(data_mid_1_47_imag));
  assign _zz_4372 = fixTo_330_dout;
  assign _zz_4373 = ($signed(_zz_278) + $signed(_zz_4374));
  assign _zz_4374 = ($signed(_zz_4375) * $signed(twiddle_factor_table_2_real));
  assign _zz_4375 = ($signed(data_mid_1_47_imag) - $signed(data_mid_1_47_real));
  assign _zz_4376 = fixTo_331_dout;
  assign _zz_4377 = _zz_4378[35 : 0];
  assign _zz_4378 = _zz_4379;
  assign _zz_4379 = ($signed(_zz_4380) >>> _zz_279);
  assign _zz_4380 = _zz_4381;
  assign _zz_4381 = ($signed(_zz_4383) - $signed(_zz_276));
  assign _zz_4382 = ({9'd0,data_mid_1_45_real} <<< 9);
  assign _zz_4383 = {{9{_zz_4382[26]}}, _zz_4382};
  assign _zz_4384 = fixTo_332_dout;
  assign _zz_4385 = _zz_4386[35 : 0];
  assign _zz_4386 = _zz_4387;
  assign _zz_4387 = ($signed(_zz_4388) >>> _zz_279);
  assign _zz_4388 = _zz_4389;
  assign _zz_4389 = ($signed(_zz_4391) - $signed(_zz_277));
  assign _zz_4390 = ({9'd0,data_mid_1_45_imag} <<< 9);
  assign _zz_4391 = {{9{_zz_4390[26]}}, _zz_4390};
  assign _zz_4392 = fixTo_333_dout;
  assign _zz_4393 = _zz_4394[35 : 0];
  assign _zz_4394 = _zz_4395;
  assign _zz_4395 = ($signed(_zz_4396) >>> _zz_280);
  assign _zz_4396 = _zz_4397;
  assign _zz_4397 = ($signed(_zz_4399) + $signed(_zz_276));
  assign _zz_4398 = ({9'd0,data_mid_1_45_real} <<< 9);
  assign _zz_4399 = {{9{_zz_4398[26]}}, _zz_4398};
  assign _zz_4400 = fixTo_334_dout;
  assign _zz_4401 = _zz_4402[35 : 0];
  assign _zz_4402 = _zz_4403;
  assign _zz_4403 = ($signed(_zz_4404) >>> _zz_280);
  assign _zz_4404 = _zz_4405;
  assign _zz_4405 = ($signed(_zz_4407) + $signed(_zz_277));
  assign _zz_4406 = ({9'd0,data_mid_1_45_imag} <<< 9);
  assign _zz_4407 = {{9{_zz_4406[26]}}, _zz_4406};
  assign _zz_4408 = fixTo_335_dout;
  assign _zz_4409 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_4410 = ($signed(_zz_283) - $signed(_zz_4411));
  assign _zz_4411 = ($signed(_zz_4412) * $signed(twiddle_factor_table_1_imag));
  assign _zz_4412 = ($signed(data_mid_1_50_real) + $signed(data_mid_1_50_imag));
  assign _zz_4413 = fixTo_336_dout;
  assign _zz_4414 = ($signed(_zz_283) + $signed(_zz_4415));
  assign _zz_4415 = ($signed(_zz_4416) * $signed(twiddle_factor_table_1_real));
  assign _zz_4416 = ($signed(data_mid_1_50_imag) - $signed(data_mid_1_50_real));
  assign _zz_4417 = fixTo_337_dout;
  assign _zz_4418 = _zz_4419[35 : 0];
  assign _zz_4419 = _zz_4420;
  assign _zz_4420 = ($signed(_zz_4421) >>> _zz_284);
  assign _zz_4421 = _zz_4422;
  assign _zz_4422 = ($signed(_zz_4424) - $signed(_zz_281));
  assign _zz_4423 = ({9'd0,data_mid_1_48_real} <<< 9);
  assign _zz_4424 = {{9{_zz_4423[26]}}, _zz_4423};
  assign _zz_4425 = fixTo_338_dout;
  assign _zz_4426 = _zz_4427[35 : 0];
  assign _zz_4427 = _zz_4428;
  assign _zz_4428 = ($signed(_zz_4429) >>> _zz_284);
  assign _zz_4429 = _zz_4430;
  assign _zz_4430 = ($signed(_zz_4432) - $signed(_zz_282));
  assign _zz_4431 = ({9'd0,data_mid_1_48_imag} <<< 9);
  assign _zz_4432 = {{9{_zz_4431[26]}}, _zz_4431};
  assign _zz_4433 = fixTo_339_dout;
  assign _zz_4434 = _zz_4435[35 : 0];
  assign _zz_4435 = _zz_4436;
  assign _zz_4436 = ($signed(_zz_4437) >>> _zz_285);
  assign _zz_4437 = _zz_4438;
  assign _zz_4438 = ($signed(_zz_4440) + $signed(_zz_281));
  assign _zz_4439 = ({9'd0,data_mid_1_48_real} <<< 9);
  assign _zz_4440 = {{9{_zz_4439[26]}}, _zz_4439};
  assign _zz_4441 = fixTo_340_dout;
  assign _zz_4442 = _zz_4443[35 : 0];
  assign _zz_4443 = _zz_4444;
  assign _zz_4444 = ($signed(_zz_4445) >>> _zz_285);
  assign _zz_4445 = _zz_4446;
  assign _zz_4446 = ($signed(_zz_4448) + $signed(_zz_282));
  assign _zz_4447 = ({9'd0,data_mid_1_48_imag} <<< 9);
  assign _zz_4448 = {{9{_zz_4447[26]}}, _zz_4447};
  assign _zz_4449 = fixTo_341_dout;
  assign _zz_4450 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_4451 = ($signed(_zz_288) - $signed(_zz_4452));
  assign _zz_4452 = ($signed(_zz_4453) * $signed(twiddle_factor_table_2_imag));
  assign _zz_4453 = ($signed(data_mid_1_51_real) + $signed(data_mid_1_51_imag));
  assign _zz_4454 = fixTo_342_dout;
  assign _zz_4455 = ($signed(_zz_288) + $signed(_zz_4456));
  assign _zz_4456 = ($signed(_zz_4457) * $signed(twiddle_factor_table_2_real));
  assign _zz_4457 = ($signed(data_mid_1_51_imag) - $signed(data_mid_1_51_real));
  assign _zz_4458 = fixTo_343_dout;
  assign _zz_4459 = _zz_4460[35 : 0];
  assign _zz_4460 = _zz_4461;
  assign _zz_4461 = ($signed(_zz_4462) >>> _zz_289);
  assign _zz_4462 = _zz_4463;
  assign _zz_4463 = ($signed(_zz_4465) - $signed(_zz_286));
  assign _zz_4464 = ({9'd0,data_mid_1_49_real} <<< 9);
  assign _zz_4465 = {{9{_zz_4464[26]}}, _zz_4464};
  assign _zz_4466 = fixTo_344_dout;
  assign _zz_4467 = _zz_4468[35 : 0];
  assign _zz_4468 = _zz_4469;
  assign _zz_4469 = ($signed(_zz_4470) >>> _zz_289);
  assign _zz_4470 = _zz_4471;
  assign _zz_4471 = ($signed(_zz_4473) - $signed(_zz_287));
  assign _zz_4472 = ({9'd0,data_mid_1_49_imag} <<< 9);
  assign _zz_4473 = {{9{_zz_4472[26]}}, _zz_4472};
  assign _zz_4474 = fixTo_345_dout;
  assign _zz_4475 = _zz_4476[35 : 0];
  assign _zz_4476 = _zz_4477;
  assign _zz_4477 = ($signed(_zz_4478) >>> _zz_290);
  assign _zz_4478 = _zz_4479;
  assign _zz_4479 = ($signed(_zz_4481) + $signed(_zz_286));
  assign _zz_4480 = ({9'd0,data_mid_1_49_real} <<< 9);
  assign _zz_4481 = {{9{_zz_4480[26]}}, _zz_4480};
  assign _zz_4482 = fixTo_346_dout;
  assign _zz_4483 = _zz_4484[35 : 0];
  assign _zz_4484 = _zz_4485;
  assign _zz_4485 = ($signed(_zz_4486) >>> _zz_290);
  assign _zz_4486 = _zz_4487;
  assign _zz_4487 = ($signed(_zz_4489) + $signed(_zz_287));
  assign _zz_4488 = ({9'd0,data_mid_1_49_imag} <<< 9);
  assign _zz_4489 = {{9{_zz_4488[26]}}, _zz_4488};
  assign _zz_4490 = fixTo_347_dout;
  assign _zz_4491 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_4492 = ($signed(_zz_293) - $signed(_zz_4493));
  assign _zz_4493 = ($signed(_zz_4494) * $signed(twiddle_factor_table_1_imag));
  assign _zz_4494 = ($signed(data_mid_1_54_real) + $signed(data_mid_1_54_imag));
  assign _zz_4495 = fixTo_348_dout;
  assign _zz_4496 = ($signed(_zz_293) + $signed(_zz_4497));
  assign _zz_4497 = ($signed(_zz_4498) * $signed(twiddle_factor_table_1_real));
  assign _zz_4498 = ($signed(data_mid_1_54_imag) - $signed(data_mid_1_54_real));
  assign _zz_4499 = fixTo_349_dout;
  assign _zz_4500 = _zz_4501[35 : 0];
  assign _zz_4501 = _zz_4502;
  assign _zz_4502 = ($signed(_zz_4503) >>> _zz_294);
  assign _zz_4503 = _zz_4504;
  assign _zz_4504 = ($signed(_zz_4506) - $signed(_zz_291));
  assign _zz_4505 = ({9'd0,data_mid_1_52_real} <<< 9);
  assign _zz_4506 = {{9{_zz_4505[26]}}, _zz_4505};
  assign _zz_4507 = fixTo_350_dout;
  assign _zz_4508 = _zz_4509[35 : 0];
  assign _zz_4509 = _zz_4510;
  assign _zz_4510 = ($signed(_zz_4511) >>> _zz_294);
  assign _zz_4511 = _zz_4512;
  assign _zz_4512 = ($signed(_zz_4514) - $signed(_zz_292));
  assign _zz_4513 = ({9'd0,data_mid_1_52_imag} <<< 9);
  assign _zz_4514 = {{9{_zz_4513[26]}}, _zz_4513};
  assign _zz_4515 = fixTo_351_dout;
  assign _zz_4516 = _zz_4517[35 : 0];
  assign _zz_4517 = _zz_4518;
  assign _zz_4518 = ($signed(_zz_4519) >>> _zz_295);
  assign _zz_4519 = _zz_4520;
  assign _zz_4520 = ($signed(_zz_4522) + $signed(_zz_291));
  assign _zz_4521 = ({9'd0,data_mid_1_52_real} <<< 9);
  assign _zz_4522 = {{9{_zz_4521[26]}}, _zz_4521};
  assign _zz_4523 = fixTo_352_dout;
  assign _zz_4524 = _zz_4525[35 : 0];
  assign _zz_4525 = _zz_4526;
  assign _zz_4526 = ($signed(_zz_4527) >>> _zz_295);
  assign _zz_4527 = _zz_4528;
  assign _zz_4528 = ($signed(_zz_4530) + $signed(_zz_292));
  assign _zz_4529 = ({9'd0,data_mid_1_52_imag} <<< 9);
  assign _zz_4530 = {{9{_zz_4529[26]}}, _zz_4529};
  assign _zz_4531 = fixTo_353_dout;
  assign _zz_4532 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_4533 = ($signed(_zz_298) - $signed(_zz_4534));
  assign _zz_4534 = ($signed(_zz_4535) * $signed(twiddle_factor_table_2_imag));
  assign _zz_4535 = ($signed(data_mid_1_55_real) + $signed(data_mid_1_55_imag));
  assign _zz_4536 = fixTo_354_dout;
  assign _zz_4537 = ($signed(_zz_298) + $signed(_zz_4538));
  assign _zz_4538 = ($signed(_zz_4539) * $signed(twiddle_factor_table_2_real));
  assign _zz_4539 = ($signed(data_mid_1_55_imag) - $signed(data_mid_1_55_real));
  assign _zz_4540 = fixTo_355_dout;
  assign _zz_4541 = _zz_4542[35 : 0];
  assign _zz_4542 = _zz_4543;
  assign _zz_4543 = ($signed(_zz_4544) >>> _zz_299);
  assign _zz_4544 = _zz_4545;
  assign _zz_4545 = ($signed(_zz_4547) - $signed(_zz_296));
  assign _zz_4546 = ({9'd0,data_mid_1_53_real} <<< 9);
  assign _zz_4547 = {{9{_zz_4546[26]}}, _zz_4546};
  assign _zz_4548 = fixTo_356_dout;
  assign _zz_4549 = _zz_4550[35 : 0];
  assign _zz_4550 = _zz_4551;
  assign _zz_4551 = ($signed(_zz_4552) >>> _zz_299);
  assign _zz_4552 = _zz_4553;
  assign _zz_4553 = ($signed(_zz_4555) - $signed(_zz_297));
  assign _zz_4554 = ({9'd0,data_mid_1_53_imag} <<< 9);
  assign _zz_4555 = {{9{_zz_4554[26]}}, _zz_4554};
  assign _zz_4556 = fixTo_357_dout;
  assign _zz_4557 = _zz_4558[35 : 0];
  assign _zz_4558 = _zz_4559;
  assign _zz_4559 = ($signed(_zz_4560) >>> _zz_300);
  assign _zz_4560 = _zz_4561;
  assign _zz_4561 = ($signed(_zz_4563) + $signed(_zz_296));
  assign _zz_4562 = ({9'd0,data_mid_1_53_real} <<< 9);
  assign _zz_4563 = {{9{_zz_4562[26]}}, _zz_4562};
  assign _zz_4564 = fixTo_358_dout;
  assign _zz_4565 = _zz_4566[35 : 0];
  assign _zz_4566 = _zz_4567;
  assign _zz_4567 = ($signed(_zz_4568) >>> _zz_300);
  assign _zz_4568 = _zz_4569;
  assign _zz_4569 = ($signed(_zz_4571) + $signed(_zz_297));
  assign _zz_4570 = ({9'd0,data_mid_1_53_imag} <<< 9);
  assign _zz_4571 = {{9{_zz_4570[26]}}, _zz_4570};
  assign _zz_4572 = fixTo_359_dout;
  assign _zz_4573 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_4574 = ($signed(_zz_303) - $signed(_zz_4575));
  assign _zz_4575 = ($signed(_zz_4576) * $signed(twiddle_factor_table_1_imag));
  assign _zz_4576 = ($signed(data_mid_1_58_real) + $signed(data_mid_1_58_imag));
  assign _zz_4577 = fixTo_360_dout;
  assign _zz_4578 = ($signed(_zz_303) + $signed(_zz_4579));
  assign _zz_4579 = ($signed(_zz_4580) * $signed(twiddle_factor_table_1_real));
  assign _zz_4580 = ($signed(data_mid_1_58_imag) - $signed(data_mid_1_58_real));
  assign _zz_4581 = fixTo_361_dout;
  assign _zz_4582 = _zz_4583[35 : 0];
  assign _zz_4583 = _zz_4584;
  assign _zz_4584 = ($signed(_zz_4585) >>> _zz_304);
  assign _zz_4585 = _zz_4586;
  assign _zz_4586 = ($signed(_zz_4588) - $signed(_zz_301));
  assign _zz_4587 = ({9'd0,data_mid_1_56_real} <<< 9);
  assign _zz_4588 = {{9{_zz_4587[26]}}, _zz_4587};
  assign _zz_4589 = fixTo_362_dout;
  assign _zz_4590 = _zz_4591[35 : 0];
  assign _zz_4591 = _zz_4592;
  assign _zz_4592 = ($signed(_zz_4593) >>> _zz_304);
  assign _zz_4593 = _zz_4594;
  assign _zz_4594 = ($signed(_zz_4596) - $signed(_zz_302));
  assign _zz_4595 = ({9'd0,data_mid_1_56_imag} <<< 9);
  assign _zz_4596 = {{9{_zz_4595[26]}}, _zz_4595};
  assign _zz_4597 = fixTo_363_dout;
  assign _zz_4598 = _zz_4599[35 : 0];
  assign _zz_4599 = _zz_4600;
  assign _zz_4600 = ($signed(_zz_4601) >>> _zz_305);
  assign _zz_4601 = _zz_4602;
  assign _zz_4602 = ($signed(_zz_4604) + $signed(_zz_301));
  assign _zz_4603 = ({9'd0,data_mid_1_56_real} <<< 9);
  assign _zz_4604 = {{9{_zz_4603[26]}}, _zz_4603};
  assign _zz_4605 = fixTo_364_dout;
  assign _zz_4606 = _zz_4607[35 : 0];
  assign _zz_4607 = _zz_4608;
  assign _zz_4608 = ($signed(_zz_4609) >>> _zz_305);
  assign _zz_4609 = _zz_4610;
  assign _zz_4610 = ($signed(_zz_4612) + $signed(_zz_302));
  assign _zz_4611 = ({9'd0,data_mid_1_56_imag} <<< 9);
  assign _zz_4612 = {{9{_zz_4611[26]}}, _zz_4611};
  assign _zz_4613 = fixTo_365_dout;
  assign _zz_4614 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_4615 = ($signed(_zz_308) - $signed(_zz_4616));
  assign _zz_4616 = ($signed(_zz_4617) * $signed(twiddle_factor_table_2_imag));
  assign _zz_4617 = ($signed(data_mid_1_59_real) + $signed(data_mid_1_59_imag));
  assign _zz_4618 = fixTo_366_dout;
  assign _zz_4619 = ($signed(_zz_308) + $signed(_zz_4620));
  assign _zz_4620 = ($signed(_zz_4621) * $signed(twiddle_factor_table_2_real));
  assign _zz_4621 = ($signed(data_mid_1_59_imag) - $signed(data_mid_1_59_real));
  assign _zz_4622 = fixTo_367_dout;
  assign _zz_4623 = _zz_4624[35 : 0];
  assign _zz_4624 = _zz_4625;
  assign _zz_4625 = ($signed(_zz_4626) >>> _zz_309);
  assign _zz_4626 = _zz_4627;
  assign _zz_4627 = ($signed(_zz_4629) - $signed(_zz_306));
  assign _zz_4628 = ({9'd0,data_mid_1_57_real} <<< 9);
  assign _zz_4629 = {{9{_zz_4628[26]}}, _zz_4628};
  assign _zz_4630 = fixTo_368_dout;
  assign _zz_4631 = _zz_4632[35 : 0];
  assign _zz_4632 = _zz_4633;
  assign _zz_4633 = ($signed(_zz_4634) >>> _zz_309);
  assign _zz_4634 = _zz_4635;
  assign _zz_4635 = ($signed(_zz_4637) - $signed(_zz_307));
  assign _zz_4636 = ({9'd0,data_mid_1_57_imag} <<< 9);
  assign _zz_4637 = {{9{_zz_4636[26]}}, _zz_4636};
  assign _zz_4638 = fixTo_369_dout;
  assign _zz_4639 = _zz_4640[35 : 0];
  assign _zz_4640 = _zz_4641;
  assign _zz_4641 = ($signed(_zz_4642) >>> _zz_310);
  assign _zz_4642 = _zz_4643;
  assign _zz_4643 = ($signed(_zz_4645) + $signed(_zz_306));
  assign _zz_4644 = ({9'd0,data_mid_1_57_real} <<< 9);
  assign _zz_4645 = {{9{_zz_4644[26]}}, _zz_4644};
  assign _zz_4646 = fixTo_370_dout;
  assign _zz_4647 = _zz_4648[35 : 0];
  assign _zz_4648 = _zz_4649;
  assign _zz_4649 = ($signed(_zz_4650) >>> _zz_310);
  assign _zz_4650 = _zz_4651;
  assign _zz_4651 = ($signed(_zz_4653) + $signed(_zz_307));
  assign _zz_4652 = ({9'd0,data_mid_1_57_imag} <<< 9);
  assign _zz_4653 = {{9{_zz_4652[26]}}, _zz_4652};
  assign _zz_4654 = fixTo_371_dout;
  assign _zz_4655 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_4656 = ($signed(_zz_313) - $signed(_zz_4657));
  assign _zz_4657 = ($signed(_zz_4658) * $signed(twiddle_factor_table_1_imag));
  assign _zz_4658 = ($signed(data_mid_1_62_real) + $signed(data_mid_1_62_imag));
  assign _zz_4659 = fixTo_372_dout;
  assign _zz_4660 = ($signed(_zz_313) + $signed(_zz_4661));
  assign _zz_4661 = ($signed(_zz_4662) * $signed(twiddle_factor_table_1_real));
  assign _zz_4662 = ($signed(data_mid_1_62_imag) - $signed(data_mid_1_62_real));
  assign _zz_4663 = fixTo_373_dout;
  assign _zz_4664 = _zz_4665[35 : 0];
  assign _zz_4665 = _zz_4666;
  assign _zz_4666 = ($signed(_zz_4667) >>> _zz_314);
  assign _zz_4667 = _zz_4668;
  assign _zz_4668 = ($signed(_zz_4670) - $signed(_zz_311));
  assign _zz_4669 = ({9'd0,data_mid_1_60_real} <<< 9);
  assign _zz_4670 = {{9{_zz_4669[26]}}, _zz_4669};
  assign _zz_4671 = fixTo_374_dout;
  assign _zz_4672 = _zz_4673[35 : 0];
  assign _zz_4673 = _zz_4674;
  assign _zz_4674 = ($signed(_zz_4675) >>> _zz_314);
  assign _zz_4675 = _zz_4676;
  assign _zz_4676 = ($signed(_zz_4678) - $signed(_zz_312));
  assign _zz_4677 = ({9'd0,data_mid_1_60_imag} <<< 9);
  assign _zz_4678 = {{9{_zz_4677[26]}}, _zz_4677};
  assign _zz_4679 = fixTo_375_dout;
  assign _zz_4680 = _zz_4681[35 : 0];
  assign _zz_4681 = _zz_4682;
  assign _zz_4682 = ($signed(_zz_4683) >>> _zz_315);
  assign _zz_4683 = _zz_4684;
  assign _zz_4684 = ($signed(_zz_4686) + $signed(_zz_311));
  assign _zz_4685 = ({9'd0,data_mid_1_60_real} <<< 9);
  assign _zz_4686 = {{9{_zz_4685[26]}}, _zz_4685};
  assign _zz_4687 = fixTo_376_dout;
  assign _zz_4688 = _zz_4689[35 : 0];
  assign _zz_4689 = _zz_4690;
  assign _zz_4690 = ($signed(_zz_4691) >>> _zz_315);
  assign _zz_4691 = _zz_4692;
  assign _zz_4692 = ($signed(_zz_4694) + $signed(_zz_312));
  assign _zz_4693 = ({9'd0,data_mid_1_60_imag} <<< 9);
  assign _zz_4694 = {{9{_zz_4693[26]}}, _zz_4693};
  assign _zz_4695 = fixTo_377_dout;
  assign _zz_4696 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_4697 = ($signed(_zz_318) - $signed(_zz_4698));
  assign _zz_4698 = ($signed(_zz_4699) * $signed(twiddle_factor_table_2_imag));
  assign _zz_4699 = ($signed(data_mid_1_63_real) + $signed(data_mid_1_63_imag));
  assign _zz_4700 = fixTo_378_dout;
  assign _zz_4701 = ($signed(_zz_318) + $signed(_zz_4702));
  assign _zz_4702 = ($signed(_zz_4703) * $signed(twiddle_factor_table_2_real));
  assign _zz_4703 = ($signed(data_mid_1_63_imag) - $signed(data_mid_1_63_real));
  assign _zz_4704 = fixTo_379_dout;
  assign _zz_4705 = _zz_4706[35 : 0];
  assign _zz_4706 = _zz_4707;
  assign _zz_4707 = ($signed(_zz_4708) >>> _zz_319);
  assign _zz_4708 = _zz_4709;
  assign _zz_4709 = ($signed(_zz_4711) - $signed(_zz_316));
  assign _zz_4710 = ({9'd0,data_mid_1_61_real} <<< 9);
  assign _zz_4711 = {{9{_zz_4710[26]}}, _zz_4710};
  assign _zz_4712 = fixTo_380_dout;
  assign _zz_4713 = _zz_4714[35 : 0];
  assign _zz_4714 = _zz_4715;
  assign _zz_4715 = ($signed(_zz_4716) >>> _zz_319);
  assign _zz_4716 = _zz_4717;
  assign _zz_4717 = ($signed(_zz_4719) - $signed(_zz_317));
  assign _zz_4718 = ({9'd0,data_mid_1_61_imag} <<< 9);
  assign _zz_4719 = {{9{_zz_4718[26]}}, _zz_4718};
  assign _zz_4720 = fixTo_381_dout;
  assign _zz_4721 = _zz_4722[35 : 0];
  assign _zz_4722 = _zz_4723;
  assign _zz_4723 = ($signed(_zz_4724) >>> _zz_320);
  assign _zz_4724 = _zz_4725;
  assign _zz_4725 = ($signed(_zz_4727) + $signed(_zz_316));
  assign _zz_4726 = ({9'd0,data_mid_1_61_real} <<< 9);
  assign _zz_4727 = {{9{_zz_4726[26]}}, _zz_4726};
  assign _zz_4728 = fixTo_382_dout;
  assign _zz_4729 = _zz_4730[35 : 0];
  assign _zz_4730 = _zz_4731;
  assign _zz_4731 = ($signed(_zz_4732) >>> _zz_320);
  assign _zz_4732 = _zz_4733;
  assign _zz_4733 = ($signed(_zz_4735) + $signed(_zz_317));
  assign _zz_4734 = ({9'd0,data_mid_1_61_imag} <<< 9);
  assign _zz_4735 = {{9{_zz_4734[26]}}, _zz_4734};
  assign _zz_4736 = fixTo_383_dout;
  assign _zz_4737 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_4738 = ($signed(_zz_323) - $signed(_zz_4739));
  assign _zz_4739 = ($signed(_zz_4740) * $signed(twiddle_factor_table_3_imag));
  assign _zz_4740 = ($signed(data_mid_2_4_real) + $signed(data_mid_2_4_imag));
  assign _zz_4741 = fixTo_384_dout;
  assign _zz_4742 = ($signed(_zz_323) + $signed(_zz_4743));
  assign _zz_4743 = ($signed(_zz_4744) * $signed(twiddle_factor_table_3_real));
  assign _zz_4744 = ($signed(data_mid_2_4_imag) - $signed(data_mid_2_4_real));
  assign _zz_4745 = fixTo_385_dout;
  assign _zz_4746 = _zz_4747[35 : 0];
  assign _zz_4747 = _zz_4748;
  assign _zz_4748 = ($signed(_zz_4749) >>> _zz_324);
  assign _zz_4749 = _zz_4750;
  assign _zz_4750 = ($signed(_zz_4752) - $signed(_zz_321));
  assign _zz_4751 = ({9'd0,data_mid_2_0_real} <<< 9);
  assign _zz_4752 = {{9{_zz_4751[26]}}, _zz_4751};
  assign _zz_4753 = fixTo_386_dout;
  assign _zz_4754 = _zz_4755[35 : 0];
  assign _zz_4755 = _zz_4756;
  assign _zz_4756 = ($signed(_zz_4757) >>> _zz_324);
  assign _zz_4757 = _zz_4758;
  assign _zz_4758 = ($signed(_zz_4760) - $signed(_zz_322));
  assign _zz_4759 = ({9'd0,data_mid_2_0_imag} <<< 9);
  assign _zz_4760 = {{9{_zz_4759[26]}}, _zz_4759};
  assign _zz_4761 = fixTo_387_dout;
  assign _zz_4762 = _zz_4763[35 : 0];
  assign _zz_4763 = _zz_4764;
  assign _zz_4764 = ($signed(_zz_4765) >>> _zz_325);
  assign _zz_4765 = _zz_4766;
  assign _zz_4766 = ($signed(_zz_4768) + $signed(_zz_321));
  assign _zz_4767 = ({9'd0,data_mid_2_0_real} <<< 9);
  assign _zz_4768 = {{9{_zz_4767[26]}}, _zz_4767};
  assign _zz_4769 = fixTo_388_dout;
  assign _zz_4770 = _zz_4771[35 : 0];
  assign _zz_4771 = _zz_4772;
  assign _zz_4772 = ($signed(_zz_4773) >>> _zz_325);
  assign _zz_4773 = _zz_4774;
  assign _zz_4774 = ($signed(_zz_4776) + $signed(_zz_322));
  assign _zz_4775 = ({9'd0,data_mid_2_0_imag} <<< 9);
  assign _zz_4776 = {{9{_zz_4775[26]}}, _zz_4775};
  assign _zz_4777 = fixTo_389_dout;
  assign _zz_4778 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_4779 = ($signed(_zz_328) - $signed(_zz_4780));
  assign _zz_4780 = ($signed(_zz_4781) * $signed(twiddle_factor_table_4_imag));
  assign _zz_4781 = ($signed(data_mid_2_5_real) + $signed(data_mid_2_5_imag));
  assign _zz_4782 = fixTo_390_dout;
  assign _zz_4783 = ($signed(_zz_328) + $signed(_zz_4784));
  assign _zz_4784 = ($signed(_zz_4785) * $signed(twiddle_factor_table_4_real));
  assign _zz_4785 = ($signed(data_mid_2_5_imag) - $signed(data_mid_2_5_real));
  assign _zz_4786 = fixTo_391_dout;
  assign _zz_4787 = _zz_4788[35 : 0];
  assign _zz_4788 = _zz_4789;
  assign _zz_4789 = ($signed(_zz_4790) >>> _zz_329);
  assign _zz_4790 = _zz_4791;
  assign _zz_4791 = ($signed(_zz_4793) - $signed(_zz_326));
  assign _zz_4792 = ({9'd0,data_mid_2_1_real} <<< 9);
  assign _zz_4793 = {{9{_zz_4792[26]}}, _zz_4792};
  assign _zz_4794 = fixTo_392_dout;
  assign _zz_4795 = _zz_4796[35 : 0];
  assign _zz_4796 = _zz_4797;
  assign _zz_4797 = ($signed(_zz_4798) >>> _zz_329);
  assign _zz_4798 = _zz_4799;
  assign _zz_4799 = ($signed(_zz_4801) - $signed(_zz_327));
  assign _zz_4800 = ({9'd0,data_mid_2_1_imag} <<< 9);
  assign _zz_4801 = {{9{_zz_4800[26]}}, _zz_4800};
  assign _zz_4802 = fixTo_393_dout;
  assign _zz_4803 = _zz_4804[35 : 0];
  assign _zz_4804 = _zz_4805;
  assign _zz_4805 = ($signed(_zz_4806) >>> _zz_330);
  assign _zz_4806 = _zz_4807;
  assign _zz_4807 = ($signed(_zz_4809) + $signed(_zz_326));
  assign _zz_4808 = ({9'd0,data_mid_2_1_real} <<< 9);
  assign _zz_4809 = {{9{_zz_4808[26]}}, _zz_4808};
  assign _zz_4810 = fixTo_394_dout;
  assign _zz_4811 = _zz_4812[35 : 0];
  assign _zz_4812 = _zz_4813;
  assign _zz_4813 = ($signed(_zz_4814) >>> _zz_330);
  assign _zz_4814 = _zz_4815;
  assign _zz_4815 = ($signed(_zz_4817) + $signed(_zz_327));
  assign _zz_4816 = ({9'd0,data_mid_2_1_imag} <<< 9);
  assign _zz_4817 = {{9{_zz_4816[26]}}, _zz_4816};
  assign _zz_4818 = fixTo_395_dout;
  assign _zz_4819 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_4820 = ($signed(_zz_333) - $signed(_zz_4821));
  assign _zz_4821 = ($signed(_zz_4822) * $signed(twiddle_factor_table_5_imag));
  assign _zz_4822 = ($signed(data_mid_2_6_real) + $signed(data_mid_2_6_imag));
  assign _zz_4823 = fixTo_396_dout;
  assign _zz_4824 = ($signed(_zz_333) + $signed(_zz_4825));
  assign _zz_4825 = ($signed(_zz_4826) * $signed(twiddle_factor_table_5_real));
  assign _zz_4826 = ($signed(data_mid_2_6_imag) - $signed(data_mid_2_6_real));
  assign _zz_4827 = fixTo_397_dout;
  assign _zz_4828 = _zz_4829[35 : 0];
  assign _zz_4829 = _zz_4830;
  assign _zz_4830 = ($signed(_zz_4831) >>> _zz_334);
  assign _zz_4831 = _zz_4832;
  assign _zz_4832 = ($signed(_zz_4834) - $signed(_zz_331));
  assign _zz_4833 = ({9'd0,data_mid_2_2_real} <<< 9);
  assign _zz_4834 = {{9{_zz_4833[26]}}, _zz_4833};
  assign _zz_4835 = fixTo_398_dout;
  assign _zz_4836 = _zz_4837[35 : 0];
  assign _zz_4837 = _zz_4838;
  assign _zz_4838 = ($signed(_zz_4839) >>> _zz_334);
  assign _zz_4839 = _zz_4840;
  assign _zz_4840 = ($signed(_zz_4842) - $signed(_zz_332));
  assign _zz_4841 = ({9'd0,data_mid_2_2_imag} <<< 9);
  assign _zz_4842 = {{9{_zz_4841[26]}}, _zz_4841};
  assign _zz_4843 = fixTo_399_dout;
  assign _zz_4844 = _zz_4845[35 : 0];
  assign _zz_4845 = _zz_4846;
  assign _zz_4846 = ($signed(_zz_4847) >>> _zz_335);
  assign _zz_4847 = _zz_4848;
  assign _zz_4848 = ($signed(_zz_4850) + $signed(_zz_331));
  assign _zz_4849 = ({9'd0,data_mid_2_2_real} <<< 9);
  assign _zz_4850 = {{9{_zz_4849[26]}}, _zz_4849};
  assign _zz_4851 = fixTo_400_dout;
  assign _zz_4852 = _zz_4853[35 : 0];
  assign _zz_4853 = _zz_4854;
  assign _zz_4854 = ($signed(_zz_4855) >>> _zz_335);
  assign _zz_4855 = _zz_4856;
  assign _zz_4856 = ($signed(_zz_4858) + $signed(_zz_332));
  assign _zz_4857 = ({9'd0,data_mid_2_2_imag} <<< 9);
  assign _zz_4858 = {{9{_zz_4857[26]}}, _zz_4857};
  assign _zz_4859 = fixTo_401_dout;
  assign _zz_4860 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_4861 = ($signed(_zz_338) - $signed(_zz_4862));
  assign _zz_4862 = ($signed(_zz_4863) * $signed(twiddle_factor_table_6_imag));
  assign _zz_4863 = ($signed(data_mid_2_7_real) + $signed(data_mid_2_7_imag));
  assign _zz_4864 = fixTo_402_dout;
  assign _zz_4865 = ($signed(_zz_338) + $signed(_zz_4866));
  assign _zz_4866 = ($signed(_zz_4867) * $signed(twiddle_factor_table_6_real));
  assign _zz_4867 = ($signed(data_mid_2_7_imag) - $signed(data_mid_2_7_real));
  assign _zz_4868 = fixTo_403_dout;
  assign _zz_4869 = _zz_4870[35 : 0];
  assign _zz_4870 = _zz_4871;
  assign _zz_4871 = ($signed(_zz_4872) >>> _zz_339);
  assign _zz_4872 = _zz_4873;
  assign _zz_4873 = ($signed(_zz_4875) - $signed(_zz_336));
  assign _zz_4874 = ({9'd0,data_mid_2_3_real} <<< 9);
  assign _zz_4875 = {{9{_zz_4874[26]}}, _zz_4874};
  assign _zz_4876 = fixTo_404_dout;
  assign _zz_4877 = _zz_4878[35 : 0];
  assign _zz_4878 = _zz_4879;
  assign _zz_4879 = ($signed(_zz_4880) >>> _zz_339);
  assign _zz_4880 = _zz_4881;
  assign _zz_4881 = ($signed(_zz_4883) - $signed(_zz_337));
  assign _zz_4882 = ({9'd0,data_mid_2_3_imag} <<< 9);
  assign _zz_4883 = {{9{_zz_4882[26]}}, _zz_4882};
  assign _zz_4884 = fixTo_405_dout;
  assign _zz_4885 = _zz_4886[35 : 0];
  assign _zz_4886 = _zz_4887;
  assign _zz_4887 = ($signed(_zz_4888) >>> _zz_340);
  assign _zz_4888 = _zz_4889;
  assign _zz_4889 = ($signed(_zz_4891) + $signed(_zz_336));
  assign _zz_4890 = ({9'd0,data_mid_2_3_real} <<< 9);
  assign _zz_4891 = {{9{_zz_4890[26]}}, _zz_4890};
  assign _zz_4892 = fixTo_406_dout;
  assign _zz_4893 = _zz_4894[35 : 0];
  assign _zz_4894 = _zz_4895;
  assign _zz_4895 = ($signed(_zz_4896) >>> _zz_340);
  assign _zz_4896 = _zz_4897;
  assign _zz_4897 = ($signed(_zz_4899) + $signed(_zz_337));
  assign _zz_4898 = ({9'd0,data_mid_2_3_imag} <<< 9);
  assign _zz_4899 = {{9{_zz_4898[26]}}, _zz_4898};
  assign _zz_4900 = fixTo_407_dout;
  assign _zz_4901 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_4902 = ($signed(_zz_343) - $signed(_zz_4903));
  assign _zz_4903 = ($signed(_zz_4904) * $signed(twiddle_factor_table_3_imag));
  assign _zz_4904 = ($signed(data_mid_2_12_real) + $signed(data_mid_2_12_imag));
  assign _zz_4905 = fixTo_408_dout;
  assign _zz_4906 = ($signed(_zz_343) + $signed(_zz_4907));
  assign _zz_4907 = ($signed(_zz_4908) * $signed(twiddle_factor_table_3_real));
  assign _zz_4908 = ($signed(data_mid_2_12_imag) - $signed(data_mid_2_12_real));
  assign _zz_4909 = fixTo_409_dout;
  assign _zz_4910 = _zz_4911[35 : 0];
  assign _zz_4911 = _zz_4912;
  assign _zz_4912 = ($signed(_zz_4913) >>> _zz_344);
  assign _zz_4913 = _zz_4914;
  assign _zz_4914 = ($signed(_zz_4916) - $signed(_zz_341));
  assign _zz_4915 = ({9'd0,data_mid_2_8_real} <<< 9);
  assign _zz_4916 = {{9{_zz_4915[26]}}, _zz_4915};
  assign _zz_4917 = fixTo_410_dout;
  assign _zz_4918 = _zz_4919[35 : 0];
  assign _zz_4919 = _zz_4920;
  assign _zz_4920 = ($signed(_zz_4921) >>> _zz_344);
  assign _zz_4921 = _zz_4922;
  assign _zz_4922 = ($signed(_zz_4924) - $signed(_zz_342));
  assign _zz_4923 = ({9'd0,data_mid_2_8_imag} <<< 9);
  assign _zz_4924 = {{9{_zz_4923[26]}}, _zz_4923};
  assign _zz_4925 = fixTo_411_dout;
  assign _zz_4926 = _zz_4927[35 : 0];
  assign _zz_4927 = _zz_4928;
  assign _zz_4928 = ($signed(_zz_4929) >>> _zz_345);
  assign _zz_4929 = _zz_4930;
  assign _zz_4930 = ($signed(_zz_4932) + $signed(_zz_341));
  assign _zz_4931 = ({9'd0,data_mid_2_8_real} <<< 9);
  assign _zz_4932 = {{9{_zz_4931[26]}}, _zz_4931};
  assign _zz_4933 = fixTo_412_dout;
  assign _zz_4934 = _zz_4935[35 : 0];
  assign _zz_4935 = _zz_4936;
  assign _zz_4936 = ($signed(_zz_4937) >>> _zz_345);
  assign _zz_4937 = _zz_4938;
  assign _zz_4938 = ($signed(_zz_4940) + $signed(_zz_342));
  assign _zz_4939 = ({9'd0,data_mid_2_8_imag} <<< 9);
  assign _zz_4940 = {{9{_zz_4939[26]}}, _zz_4939};
  assign _zz_4941 = fixTo_413_dout;
  assign _zz_4942 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_4943 = ($signed(_zz_348) - $signed(_zz_4944));
  assign _zz_4944 = ($signed(_zz_4945) * $signed(twiddle_factor_table_4_imag));
  assign _zz_4945 = ($signed(data_mid_2_13_real) + $signed(data_mid_2_13_imag));
  assign _zz_4946 = fixTo_414_dout;
  assign _zz_4947 = ($signed(_zz_348) + $signed(_zz_4948));
  assign _zz_4948 = ($signed(_zz_4949) * $signed(twiddle_factor_table_4_real));
  assign _zz_4949 = ($signed(data_mid_2_13_imag) - $signed(data_mid_2_13_real));
  assign _zz_4950 = fixTo_415_dout;
  assign _zz_4951 = _zz_4952[35 : 0];
  assign _zz_4952 = _zz_4953;
  assign _zz_4953 = ($signed(_zz_4954) >>> _zz_349);
  assign _zz_4954 = _zz_4955;
  assign _zz_4955 = ($signed(_zz_4957) - $signed(_zz_346));
  assign _zz_4956 = ({9'd0,data_mid_2_9_real} <<< 9);
  assign _zz_4957 = {{9{_zz_4956[26]}}, _zz_4956};
  assign _zz_4958 = fixTo_416_dout;
  assign _zz_4959 = _zz_4960[35 : 0];
  assign _zz_4960 = _zz_4961;
  assign _zz_4961 = ($signed(_zz_4962) >>> _zz_349);
  assign _zz_4962 = _zz_4963;
  assign _zz_4963 = ($signed(_zz_4965) - $signed(_zz_347));
  assign _zz_4964 = ({9'd0,data_mid_2_9_imag} <<< 9);
  assign _zz_4965 = {{9{_zz_4964[26]}}, _zz_4964};
  assign _zz_4966 = fixTo_417_dout;
  assign _zz_4967 = _zz_4968[35 : 0];
  assign _zz_4968 = _zz_4969;
  assign _zz_4969 = ($signed(_zz_4970) >>> _zz_350);
  assign _zz_4970 = _zz_4971;
  assign _zz_4971 = ($signed(_zz_4973) + $signed(_zz_346));
  assign _zz_4972 = ({9'd0,data_mid_2_9_real} <<< 9);
  assign _zz_4973 = {{9{_zz_4972[26]}}, _zz_4972};
  assign _zz_4974 = fixTo_418_dout;
  assign _zz_4975 = _zz_4976[35 : 0];
  assign _zz_4976 = _zz_4977;
  assign _zz_4977 = ($signed(_zz_4978) >>> _zz_350);
  assign _zz_4978 = _zz_4979;
  assign _zz_4979 = ($signed(_zz_4981) + $signed(_zz_347));
  assign _zz_4980 = ({9'd0,data_mid_2_9_imag} <<< 9);
  assign _zz_4981 = {{9{_zz_4980[26]}}, _zz_4980};
  assign _zz_4982 = fixTo_419_dout;
  assign _zz_4983 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_4984 = ($signed(_zz_353) - $signed(_zz_4985));
  assign _zz_4985 = ($signed(_zz_4986) * $signed(twiddle_factor_table_5_imag));
  assign _zz_4986 = ($signed(data_mid_2_14_real) + $signed(data_mid_2_14_imag));
  assign _zz_4987 = fixTo_420_dout;
  assign _zz_4988 = ($signed(_zz_353) + $signed(_zz_4989));
  assign _zz_4989 = ($signed(_zz_4990) * $signed(twiddle_factor_table_5_real));
  assign _zz_4990 = ($signed(data_mid_2_14_imag) - $signed(data_mid_2_14_real));
  assign _zz_4991 = fixTo_421_dout;
  assign _zz_4992 = _zz_4993[35 : 0];
  assign _zz_4993 = _zz_4994;
  assign _zz_4994 = ($signed(_zz_4995) >>> _zz_354);
  assign _zz_4995 = _zz_4996;
  assign _zz_4996 = ($signed(_zz_4998) - $signed(_zz_351));
  assign _zz_4997 = ({9'd0,data_mid_2_10_real} <<< 9);
  assign _zz_4998 = {{9{_zz_4997[26]}}, _zz_4997};
  assign _zz_4999 = fixTo_422_dout;
  assign _zz_5000 = _zz_5001[35 : 0];
  assign _zz_5001 = _zz_5002;
  assign _zz_5002 = ($signed(_zz_5003) >>> _zz_354);
  assign _zz_5003 = _zz_5004;
  assign _zz_5004 = ($signed(_zz_5006) - $signed(_zz_352));
  assign _zz_5005 = ({9'd0,data_mid_2_10_imag} <<< 9);
  assign _zz_5006 = {{9{_zz_5005[26]}}, _zz_5005};
  assign _zz_5007 = fixTo_423_dout;
  assign _zz_5008 = _zz_5009[35 : 0];
  assign _zz_5009 = _zz_5010;
  assign _zz_5010 = ($signed(_zz_5011) >>> _zz_355);
  assign _zz_5011 = _zz_5012;
  assign _zz_5012 = ($signed(_zz_5014) + $signed(_zz_351));
  assign _zz_5013 = ({9'd0,data_mid_2_10_real} <<< 9);
  assign _zz_5014 = {{9{_zz_5013[26]}}, _zz_5013};
  assign _zz_5015 = fixTo_424_dout;
  assign _zz_5016 = _zz_5017[35 : 0];
  assign _zz_5017 = _zz_5018;
  assign _zz_5018 = ($signed(_zz_5019) >>> _zz_355);
  assign _zz_5019 = _zz_5020;
  assign _zz_5020 = ($signed(_zz_5022) + $signed(_zz_352));
  assign _zz_5021 = ({9'd0,data_mid_2_10_imag} <<< 9);
  assign _zz_5022 = {{9{_zz_5021[26]}}, _zz_5021};
  assign _zz_5023 = fixTo_425_dout;
  assign _zz_5024 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_5025 = ($signed(_zz_358) - $signed(_zz_5026));
  assign _zz_5026 = ($signed(_zz_5027) * $signed(twiddle_factor_table_6_imag));
  assign _zz_5027 = ($signed(data_mid_2_15_real) + $signed(data_mid_2_15_imag));
  assign _zz_5028 = fixTo_426_dout;
  assign _zz_5029 = ($signed(_zz_358) + $signed(_zz_5030));
  assign _zz_5030 = ($signed(_zz_5031) * $signed(twiddle_factor_table_6_real));
  assign _zz_5031 = ($signed(data_mid_2_15_imag) - $signed(data_mid_2_15_real));
  assign _zz_5032 = fixTo_427_dout;
  assign _zz_5033 = _zz_5034[35 : 0];
  assign _zz_5034 = _zz_5035;
  assign _zz_5035 = ($signed(_zz_5036) >>> _zz_359);
  assign _zz_5036 = _zz_5037;
  assign _zz_5037 = ($signed(_zz_5039) - $signed(_zz_356));
  assign _zz_5038 = ({9'd0,data_mid_2_11_real} <<< 9);
  assign _zz_5039 = {{9{_zz_5038[26]}}, _zz_5038};
  assign _zz_5040 = fixTo_428_dout;
  assign _zz_5041 = _zz_5042[35 : 0];
  assign _zz_5042 = _zz_5043;
  assign _zz_5043 = ($signed(_zz_5044) >>> _zz_359);
  assign _zz_5044 = _zz_5045;
  assign _zz_5045 = ($signed(_zz_5047) - $signed(_zz_357));
  assign _zz_5046 = ({9'd0,data_mid_2_11_imag} <<< 9);
  assign _zz_5047 = {{9{_zz_5046[26]}}, _zz_5046};
  assign _zz_5048 = fixTo_429_dout;
  assign _zz_5049 = _zz_5050[35 : 0];
  assign _zz_5050 = _zz_5051;
  assign _zz_5051 = ($signed(_zz_5052) >>> _zz_360);
  assign _zz_5052 = _zz_5053;
  assign _zz_5053 = ($signed(_zz_5055) + $signed(_zz_356));
  assign _zz_5054 = ({9'd0,data_mid_2_11_real} <<< 9);
  assign _zz_5055 = {{9{_zz_5054[26]}}, _zz_5054};
  assign _zz_5056 = fixTo_430_dout;
  assign _zz_5057 = _zz_5058[35 : 0];
  assign _zz_5058 = _zz_5059;
  assign _zz_5059 = ($signed(_zz_5060) >>> _zz_360);
  assign _zz_5060 = _zz_5061;
  assign _zz_5061 = ($signed(_zz_5063) + $signed(_zz_357));
  assign _zz_5062 = ({9'd0,data_mid_2_11_imag} <<< 9);
  assign _zz_5063 = {{9{_zz_5062[26]}}, _zz_5062};
  assign _zz_5064 = fixTo_431_dout;
  assign _zz_5065 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_5066 = ($signed(_zz_363) - $signed(_zz_5067));
  assign _zz_5067 = ($signed(_zz_5068) * $signed(twiddle_factor_table_3_imag));
  assign _zz_5068 = ($signed(data_mid_2_20_real) + $signed(data_mid_2_20_imag));
  assign _zz_5069 = fixTo_432_dout;
  assign _zz_5070 = ($signed(_zz_363) + $signed(_zz_5071));
  assign _zz_5071 = ($signed(_zz_5072) * $signed(twiddle_factor_table_3_real));
  assign _zz_5072 = ($signed(data_mid_2_20_imag) - $signed(data_mid_2_20_real));
  assign _zz_5073 = fixTo_433_dout;
  assign _zz_5074 = _zz_5075[35 : 0];
  assign _zz_5075 = _zz_5076;
  assign _zz_5076 = ($signed(_zz_5077) >>> _zz_364);
  assign _zz_5077 = _zz_5078;
  assign _zz_5078 = ($signed(_zz_5080) - $signed(_zz_361));
  assign _zz_5079 = ({9'd0,data_mid_2_16_real} <<< 9);
  assign _zz_5080 = {{9{_zz_5079[26]}}, _zz_5079};
  assign _zz_5081 = fixTo_434_dout;
  assign _zz_5082 = _zz_5083[35 : 0];
  assign _zz_5083 = _zz_5084;
  assign _zz_5084 = ($signed(_zz_5085) >>> _zz_364);
  assign _zz_5085 = _zz_5086;
  assign _zz_5086 = ($signed(_zz_5088) - $signed(_zz_362));
  assign _zz_5087 = ({9'd0,data_mid_2_16_imag} <<< 9);
  assign _zz_5088 = {{9{_zz_5087[26]}}, _zz_5087};
  assign _zz_5089 = fixTo_435_dout;
  assign _zz_5090 = _zz_5091[35 : 0];
  assign _zz_5091 = _zz_5092;
  assign _zz_5092 = ($signed(_zz_5093) >>> _zz_365);
  assign _zz_5093 = _zz_5094;
  assign _zz_5094 = ($signed(_zz_5096) + $signed(_zz_361));
  assign _zz_5095 = ({9'd0,data_mid_2_16_real} <<< 9);
  assign _zz_5096 = {{9{_zz_5095[26]}}, _zz_5095};
  assign _zz_5097 = fixTo_436_dout;
  assign _zz_5098 = _zz_5099[35 : 0];
  assign _zz_5099 = _zz_5100;
  assign _zz_5100 = ($signed(_zz_5101) >>> _zz_365);
  assign _zz_5101 = _zz_5102;
  assign _zz_5102 = ($signed(_zz_5104) + $signed(_zz_362));
  assign _zz_5103 = ({9'd0,data_mid_2_16_imag} <<< 9);
  assign _zz_5104 = {{9{_zz_5103[26]}}, _zz_5103};
  assign _zz_5105 = fixTo_437_dout;
  assign _zz_5106 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_5107 = ($signed(_zz_368) - $signed(_zz_5108));
  assign _zz_5108 = ($signed(_zz_5109) * $signed(twiddle_factor_table_4_imag));
  assign _zz_5109 = ($signed(data_mid_2_21_real) + $signed(data_mid_2_21_imag));
  assign _zz_5110 = fixTo_438_dout;
  assign _zz_5111 = ($signed(_zz_368) + $signed(_zz_5112));
  assign _zz_5112 = ($signed(_zz_5113) * $signed(twiddle_factor_table_4_real));
  assign _zz_5113 = ($signed(data_mid_2_21_imag) - $signed(data_mid_2_21_real));
  assign _zz_5114 = fixTo_439_dout;
  assign _zz_5115 = _zz_5116[35 : 0];
  assign _zz_5116 = _zz_5117;
  assign _zz_5117 = ($signed(_zz_5118) >>> _zz_369);
  assign _zz_5118 = _zz_5119;
  assign _zz_5119 = ($signed(_zz_5121) - $signed(_zz_366));
  assign _zz_5120 = ({9'd0,data_mid_2_17_real} <<< 9);
  assign _zz_5121 = {{9{_zz_5120[26]}}, _zz_5120};
  assign _zz_5122 = fixTo_440_dout;
  assign _zz_5123 = _zz_5124[35 : 0];
  assign _zz_5124 = _zz_5125;
  assign _zz_5125 = ($signed(_zz_5126) >>> _zz_369);
  assign _zz_5126 = _zz_5127;
  assign _zz_5127 = ($signed(_zz_5129) - $signed(_zz_367));
  assign _zz_5128 = ({9'd0,data_mid_2_17_imag} <<< 9);
  assign _zz_5129 = {{9{_zz_5128[26]}}, _zz_5128};
  assign _zz_5130 = fixTo_441_dout;
  assign _zz_5131 = _zz_5132[35 : 0];
  assign _zz_5132 = _zz_5133;
  assign _zz_5133 = ($signed(_zz_5134) >>> _zz_370);
  assign _zz_5134 = _zz_5135;
  assign _zz_5135 = ($signed(_zz_5137) + $signed(_zz_366));
  assign _zz_5136 = ({9'd0,data_mid_2_17_real} <<< 9);
  assign _zz_5137 = {{9{_zz_5136[26]}}, _zz_5136};
  assign _zz_5138 = fixTo_442_dout;
  assign _zz_5139 = _zz_5140[35 : 0];
  assign _zz_5140 = _zz_5141;
  assign _zz_5141 = ($signed(_zz_5142) >>> _zz_370);
  assign _zz_5142 = _zz_5143;
  assign _zz_5143 = ($signed(_zz_5145) + $signed(_zz_367));
  assign _zz_5144 = ({9'd0,data_mid_2_17_imag} <<< 9);
  assign _zz_5145 = {{9{_zz_5144[26]}}, _zz_5144};
  assign _zz_5146 = fixTo_443_dout;
  assign _zz_5147 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_5148 = ($signed(_zz_373) - $signed(_zz_5149));
  assign _zz_5149 = ($signed(_zz_5150) * $signed(twiddle_factor_table_5_imag));
  assign _zz_5150 = ($signed(data_mid_2_22_real) + $signed(data_mid_2_22_imag));
  assign _zz_5151 = fixTo_444_dout;
  assign _zz_5152 = ($signed(_zz_373) + $signed(_zz_5153));
  assign _zz_5153 = ($signed(_zz_5154) * $signed(twiddle_factor_table_5_real));
  assign _zz_5154 = ($signed(data_mid_2_22_imag) - $signed(data_mid_2_22_real));
  assign _zz_5155 = fixTo_445_dout;
  assign _zz_5156 = _zz_5157[35 : 0];
  assign _zz_5157 = _zz_5158;
  assign _zz_5158 = ($signed(_zz_5159) >>> _zz_374);
  assign _zz_5159 = _zz_5160;
  assign _zz_5160 = ($signed(_zz_5162) - $signed(_zz_371));
  assign _zz_5161 = ({9'd0,data_mid_2_18_real} <<< 9);
  assign _zz_5162 = {{9{_zz_5161[26]}}, _zz_5161};
  assign _zz_5163 = fixTo_446_dout;
  assign _zz_5164 = _zz_5165[35 : 0];
  assign _zz_5165 = _zz_5166;
  assign _zz_5166 = ($signed(_zz_5167) >>> _zz_374);
  assign _zz_5167 = _zz_5168;
  assign _zz_5168 = ($signed(_zz_5170) - $signed(_zz_372));
  assign _zz_5169 = ({9'd0,data_mid_2_18_imag} <<< 9);
  assign _zz_5170 = {{9{_zz_5169[26]}}, _zz_5169};
  assign _zz_5171 = fixTo_447_dout;
  assign _zz_5172 = _zz_5173[35 : 0];
  assign _zz_5173 = _zz_5174;
  assign _zz_5174 = ($signed(_zz_5175) >>> _zz_375);
  assign _zz_5175 = _zz_5176;
  assign _zz_5176 = ($signed(_zz_5178) + $signed(_zz_371));
  assign _zz_5177 = ({9'd0,data_mid_2_18_real} <<< 9);
  assign _zz_5178 = {{9{_zz_5177[26]}}, _zz_5177};
  assign _zz_5179 = fixTo_448_dout;
  assign _zz_5180 = _zz_5181[35 : 0];
  assign _zz_5181 = _zz_5182;
  assign _zz_5182 = ($signed(_zz_5183) >>> _zz_375);
  assign _zz_5183 = _zz_5184;
  assign _zz_5184 = ($signed(_zz_5186) + $signed(_zz_372));
  assign _zz_5185 = ({9'd0,data_mid_2_18_imag} <<< 9);
  assign _zz_5186 = {{9{_zz_5185[26]}}, _zz_5185};
  assign _zz_5187 = fixTo_449_dout;
  assign _zz_5188 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_5189 = ($signed(_zz_378) - $signed(_zz_5190));
  assign _zz_5190 = ($signed(_zz_5191) * $signed(twiddle_factor_table_6_imag));
  assign _zz_5191 = ($signed(data_mid_2_23_real) + $signed(data_mid_2_23_imag));
  assign _zz_5192 = fixTo_450_dout;
  assign _zz_5193 = ($signed(_zz_378) + $signed(_zz_5194));
  assign _zz_5194 = ($signed(_zz_5195) * $signed(twiddle_factor_table_6_real));
  assign _zz_5195 = ($signed(data_mid_2_23_imag) - $signed(data_mid_2_23_real));
  assign _zz_5196 = fixTo_451_dout;
  assign _zz_5197 = _zz_5198[35 : 0];
  assign _zz_5198 = _zz_5199;
  assign _zz_5199 = ($signed(_zz_5200) >>> _zz_379);
  assign _zz_5200 = _zz_5201;
  assign _zz_5201 = ($signed(_zz_5203) - $signed(_zz_376));
  assign _zz_5202 = ({9'd0,data_mid_2_19_real} <<< 9);
  assign _zz_5203 = {{9{_zz_5202[26]}}, _zz_5202};
  assign _zz_5204 = fixTo_452_dout;
  assign _zz_5205 = _zz_5206[35 : 0];
  assign _zz_5206 = _zz_5207;
  assign _zz_5207 = ($signed(_zz_5208) >>> _zz_379);
  assign _zz_5208 = _zz_5209;
  assign _zz_5209 = ($signed(_zz_5211) - $signed(_zz_377));
  assign _zz_5210 = ({9'd0,data_mid_2_19_imag} <<< 9);
  assign _zz_5211 = {{9{_zz_5210[26]}}, _zz_5210};
  assign _zz_5212 = fixTo_453_dout;
  assign _zz_5213 = _zz_5214[35 : 0];
  assign _zz_5214 = _zz_5215;
  assign _zz_5215 = ($signed(_zz_5216) >>> _zz_380);
  assign _zz_5216 = _zz_5217;
  assign _zz_5217 = ($signed(_zz_5219) + $signed(_zz_376));
  assign _zz_5218 = ({9'd0,data_mid_2_19_real} <<< 9);
  assign _zz_5219 = {{9{_zz_5218[26]}}, _zz_5218};
  assign _zz_5220 = fixTo_454_dout;
  assign _zz_5221 = _zz_5222[35 : 0];
  assign _zz_5222 = _zz_5223;
  assign _zz_5223 = ($signed(_zz_5224) >>> _zz_380);
  assign _zz_5224 = _zz_5225;
  assign _zz_5225 = ($signed(_zz_5227) + $signed(_zz_377));
  assign _zz_5226 = ({9'd0,data_mid_2_19_imag} <<< 9);
  assign _zz_5227 = {{9{_zz_5226[26]}}, _zz_5226};
  assign _zz_5228 = fixTo_455_dout;
  assign _zz_5229 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_5230 = ($signed(_zz_383) - $signed(_zz_5231));
  assign _zz_5231 = ($signed(_zz_5232) * $signed(twiddle_factor_table_3_imag));
  assign _zz_5232 = ($signed(data_mid_2_28_real) + $signed(data_mid_2_28_imag));
  assign _zz_5233 = fixTo_456_dout;
  assign _zz_5234 = ($signed(_zz_383) + $signed(_zz_5235));
  assign _zz_5235 = ($signed(_zz_5236) * $signed(twiddle_factor_table_3_real));
  assign _zz_5236 = ($signed(data_mid_2_28_imag) - $signed(data_mid_2_28_real));
  assign _zz_5237 = fixTo_457_dout;
  assign _zz_5238 = _zz_5239[35 : 0];
  assign _zz_5239 = _zz_5240;
  assign _zz_5240 = ($signed(_zz_5241) >>> _zz_384);
  assign _zz_5241 = _zz_5242;
  assign _zz_5242 = ($signed(_zz_5244) - $signed(_zz_381));
  assign _zz_5243 = ({9'd0,data_mid_2_24_real} <<< 9);
  assign _zz_5244 = {{9{_zz_5243[26]}}, _zz_5243};
  assign _zz_5245 = fixTo_458_dout;
  assign _zz_5246 = _zz_5247[35 : 0];
  assign _zz_5247 = _zz_5248;
  assign _zz_5248 = ($signed(_zz_5249) >>> _zz_384);
  assign _zz_5249 = _zz_5250;
  assign _zz_5250 = ($signed(_zz_5252) - $signed(_zz_382));
  assign _zz_5251 = ({9'd0,data_mid_2_24_imag} <<< 9);
  assign _zz_5252 = {{9{_zz_5251[26]}}, _zz_5251};
  assign _zz_5253 = fixTo_459_dout;
  assign _zz_5254 = _zz_5255[35 : 0];
  assign _zz_5255 = _zz_5256;
  assign _zz_5256 = ($signed(_zz_5257) >>> _zz_385);
  assign _zz_5257 = _zz_5258;
  assign _zz_5258 = ($signed(_zz_5260) + $signed(_zz_381));
  assign _zz_5259 = ({9'd0,data_mid_2_24_real} <<< 9);
  assign _zz_5260 = {{9{_zz_5259[26]}}, _zz_5259};
  assign _zz_5261 = fixTo_460_dout;
  assign _zz_5262 = _zz_5263[35 : 0];
  assign _zz_5263 = _zz_5264;
  assign _zz_5264 = ($signed(_zz_5265) >>> _zz_385);
  assign _zz_5265 = _zz_5266;
  assign _zz_5266 = ($signed(_zz_5268) + $signed(_zz_382));
  assign _zz_5267 = ({9'd0,data_mid_2_24_imag} <<< 9);
  assign _zz_5268 = {{9{_zz_5267[26]}}, _zz_5267};
  assign _zz_5269 = fixTo_461_dout;
  assign _zz_5270 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_5271 = ($signed(_zz_388) - $signed(_zz_5272));
  assign _zz_5272 = ($signed(_zz_5273) * $signed(twiddle_factor_table_4_imag));
  assign _zz_5273 = ($signed(data_mid_2_29_real) + $signed(data_mid_2_29_imag));
  assign _zz_5274 = fixTo_462_dout;
  assign _zz_5275 = ($signed(_zz_388) + $signed(_zz_5276));
  assign _zz_5276 = ($signed(_zz_5277) * $signed(twiddle_factor_table_4_real));
  assign _zz_5277 = ($signed(data_mid_2_29_imag) - $signed(data_mid_2_29_real));
  assign _zz_5278 = fixTo_463_dout;
  assign _zz_5279 = _zz_5280[35 : 0];
  assign _zz_5280 = _zz_5281;
  assign _zz_5281 = ($signed(_zz_5282) >>> _zz_389);
  assign _zz_5282 = _zz_5283;
  assign _zz_5283 = ($signed(_zz_5285) - $signed(_zz_386));
  assign _zz_5284 = ({9'd0,data_mid_2_25_real} <<< 9);
  assign _zz_5285 = {{9{_zz_5284[26]}}, _zz_5284};
  assign _zz_5286 = fixTo_464_dout;
  assign _zz_5287 = _zz_5288[35 : 0];
  assign _zz_5288 = _zz_5289;
  assign _zz_5289 = ($signed(_zz_5290) >>> _zz_389);
  assign _zz_5290 = _zz_5291;
  assign _zz_5291 = ($signed(_zz_5293) - $signed(_zz_387));
  assign _zz_5292 = ({9'd0,data_mid_2_25_imag} <<< 9);
  assign _zz_5293 = {{9{_zz_5292[26]}}, _zz_5292};
  assign _zz_5294 = fixTo_465_dout;
  assign _zz_5295 = _zz_5296[35 : 0];
  assign _zz_5296 = _zz_5297;
  assign _zz_5297 = ($signed(_zz_5298) >>> _zz_390);
  assign _zz_5298 = _zz_5299;
  assign _zz_5299 = ($signed(_zz_5301) + $signed(_zz_386));
  assign _zz_5300 = ({9'd0,data_mid_2_25_real} <<< 9);
  assign _zz_5301 = {{9{_zz_5300[26]}}, _zz_5300};
  assign _zz_5302 = fixTo_466_dout;
  assign _zz_5303 = _zz_5304[35 : 0];
  assign _zz_5304 = _zz_5305;
  assign _zz_5305 = ($signed(_zz_5306) >>> _zz_390);
  assign _zz_5306 = _zz_5307;
  assign _zz_5307 = ($signed(_zz_5309) + $signed(_zz_387));
  assign _zz_5308 = ({9'd0,data_mid_2_25_imag} <<< 9);
  assign _zz_5309 = {{9{_zz_5308[26]}}, _zz_5308};
  assign _zz_5310 = fixTo_467_dout;
  assign _zz_5311 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_5312 = ($signed(_zz_393) - $signed(_zz_5313));
  assign _zz_5313 = ($signed(_zz_5314) * $signed(twiddle_factor_table_5_imag));
  assign _zz_5314 = ($signed(data_mid_2_30_real) + $signed(data_mid_2_30_imag));
  assign _zz_5315 = fixTo_468_dout;
  assign _zz_5316 = ($signed(_zz_393) + $signed(_zz_5317));
  assign _zz_5317 = ($signed(_zz_5318) * $signed(twiddle_factor_table_5_real));
  assign _zz_5318 = ($signed(data_mid_2_30_imag) - $signed(data_mid_2_30_real));
  assign _zz_5319 = fixTo_469_dout;
  assign _zz_5320 = _zz_5321[35 : 0];
  assign _zz_5321 = _zz_5322;
  assign _zz_5322 = ($signed(_zz_5323) >>> _zz_394);
  assign _zz_5323 = _zz_5324;
  assign _zz_5324 = ($signed(_zz_5326) - $signed(_zz_391));
  assign _zz_5325 = ({9'd0,data_mid_2_26_real} <<< 9);
  assign _zz_5326 = {{9{_zz_5325[26]}}, _zz_5325};
  assign _zz_5327 = fixTo_470_dout;
  assign _zz_5328 = _zz_5329[35 : 0];
  assign _zz_5329 = _zz_5330;
  assign _zz_5330 = ($signed(_zz_5331) >>> _zz_394);
  assign _zz_5331 = _zz_5332;
  assign _zz_5332 = ($signed(_zz_5334) - $signed(_zz_392));
  assign _zz_5333 = ({9'd0,data_mid_2_26_imag} <<< 9);
  assign _zz_5334 = {{9{_zz_5333[26]}}, _zz_5333};
  assign _zz_5335 = fixTo_471_dout;
  assign _zz_5336 = _zz_5337[35 : 0];
  assign _zz_5337 = _zz_5338;
  assign _zz_5338 = ($signed(_zz_5339) >>> _zz_395);
  assign _zz_5339 = _zz_5340;
  assign _zz_5340 = ($signed(_zz_5342) + $signed(_zz_391));
  assign _zz_5341 = ({9'd0,data_mid_2_26_real} <<< 9);
  assign _zz_5342 = {{9{_zz_5341[26]}}, _zz_5341};
  assign _zz_5343 = fixTo_472_dout;
  assign _zz_5344 = _zz_5345[35 : 0];
  assign _zz_5345 = _zz_5346;
  assign _zz_5346 = ($signed(_zz_5347) >>> _zz_395);
  assign _zz_5347 = _zz_5348;
  assign _zz_5348 = ($signed(_zz_5350) + $signed(_zz_392));
  assign _zz_5349 = ({9'd0,data_mid_2_26_imag} <<< 9);
  assign _zz_5350 = {{9{_zz_5349[26]}}, _zz_5349};
  assign _zz_5351 = fixTo_473_dout;
  assign _zz_5352 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_5353 = ($signed(_zz_398) - $signed(_zz_5354));
  assign _zz_5354 = ($signed(_zz_5355) * $signed(twiddle_factor_table_6_imag));
  assign _zz_5355 = ($signed(data_mid_2_31_real) + $signed(data_mid_2_31_imag));
  assign _zz_5356 = fixTo_474_dout;
  assign _zz_5357 = ($signed(_zz_398) + $signed(_zz_5358));
  assign _zz_5358 = ($signed(_zz_5359) * $signed(twiddle_factor_table_6_real));
  assign _zz_5359 = ($signed(data_mid_2_31_imag) - $signed(data_mid_2_31_real));
  assign _zz_5360 = fixTo_475_dout;
  assign _zz_5361 = _zz_5362[35 : 0];
  assign _zz_5362 = _zz_5363;
  assign _zz_5363 = ($signed(_zz_5364) >>> _zz_399);
  assign _zz_5364 = _zz_5365;
  assign _zz_5365 = ($signed(_zz_5367) - $signed(_zz_396));
  assign _zz_5366 = ({9'd0,data_mid_2_27_real} <<< 9);
  assign _zz_5367 = {{9{_zz_5366[26]}}, _zz_5366};
  assign _zz_5368 = fixTo_476_dout;
  assign _zz_5369 = _zz_5370[35 : 0];
  assign _zz_5370 = _zz_5371;
  assign _zz_5371 = ($signed(_zz_5372) >>> _zz_399);
  assign _zz_5372 = _zz_5373;
  assign _zz_5373 = ($signed(_zz_5375) - $signed(_zz_397));
  assign _zz_5374 = ({9'd0,data_mid_2_27_imag} <<< 9);
  assign _zz_5375 = {{9{_zz_5374[26]}}, _zz_5374};
  assign _zz_5376 = fixTo_477_dout;
  assign _zz_5377 = _zz_5378[35 : 0];
  assign _zz_5378 = _zz_5379;
  assign _zz_5379 = ($signed(_zz_5380) >>> _zz_400);
  assign _zz_5380 = _zz_5381;
  assign _zz_5381 = ($signed(_zz_5383) + $signed(_zz_396));
  assign _zz_5382 = ({9'd0,data_mid_2_27_real} <<< 9);
  assign _zz_5383 = {{9{_zz_5382[26]}}, _zz_5382};
  assign _zz_5384 = fixTo_478_dout;
  assign _zz_5385 = _zz_5386[35 : 0];
  assign _zz_5386 = _zz_5387;
  assign _zz_5387 = ($signed(_zz_5388) >>> _zz_400);
  assign _zz_5388 = _zz_5389;
  assign _zz_5389 = ($signed(_zz_5391) + $signed(_zz_397));
  assign _zz_5390 = ({9'd0,data_mid_2_27_imag} <<< 9);
  assign _zz_5391 = {{9{_zz_5390[26]}}, _zz_5390};
  assign _zz_5392 = fixTo_479_dout;
  assign _zz_5393 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_5394 = ($signed(_zz_403) - $signed(_zz_5395));
  assign _zz_5395 = ($signed(_zz_5396) * $signed(twiddle_factor_table_3_imag));
  assign _zz_5396 = ($signed(data_mid_2_36_real) + $signed(data_mid_2_36_imag));
  assign _zz_5397 = fixTo_480_dout;
  assign _zz_5398 = ($signed(_zz_403) + $signed(_zz_5399));
  assign _zz_5399 = ($signed(_zz_5400) * $signed(twiddle_factor_table_3_real));
  assign _zz_5400 = ($signed(data_mid_2_36_imag) - $signed(data_mid_2_36_real));
  assign _zz_5401 = fixTo_481_dout;
  assign _zz_5402 = _zz_5403[35 : 0];
  assign _zz_5403 = _zz_5404;
  assign _zz_5404 = ($signed(_zz_5405) >>> _zz_404);
  assign _zz_5405 = _zz_5406;
  assign _zz_5406 = ($signed(_zz_5408) - $signed(_zz_401));
  assign _zz_5407 = ({9'd0,data_mid_2_32_real} <<< 9);
  assign _zz_5408 = {{9{_zz_5407[26]}}, _zz_5407};
  assign _zz_5409 = fixTo_482_dout;
  assign _zz_5410 = _zz_5411[35 : 0];
  assign _zz_5411 = _zz_5412;
  assign _zz_5412 = ($signed(_zz_5413) >>> _zz_404);
  assign _zz_5413 = _zz_5414;
  assign _zz_5414 = ($signed(_zz_5416) - $signed(_zz_402));
  assign _zz_5415 = ({9'd0,data_mid_2_32_imag} <<< 9);
  assign _zz_5416 = {{9{_zz_5415[26]}}, _zz_5415};
  assign _zz_5417 = fixTo_483_dout;
  assign _zz_5418 = _zz_5419[35 : 0];
  assign _zz_5419 = _zz_5420;
  assign _zz_5420 = ($signed(_zz_5421) >>> _zz_405);
  assign _zz_5421 = _zz_5422;
  assign _zz_5422 = ($signed(_zz_5424) + $signed(_zz_401));
  assign _zz_5423 = ({9'd0,data_mid_2_32_real} <<< 9);
  assign _zz_5424 = {{9{_zz_5423[26]}}, _zz_5423};
  assign _zz_5425 = fixTo_484_dout;
  assign _zz_5426 = _zz_5427[35 : 0];
  assign _zz_5427 = _zz_5428;
  assign _zz_5428 = ($signed(_zz_5429) >>> _zz_405);
  assign _zz_5429 = _zz_5430;
  assign _zz_5430 = ($signed(_zz_5432) + $signed(_zz_402));
  assign _zz_5431 = ({9'd0,data_mid_2_32_imag} <<< 9);
  assign _zz_5432 = {{9{_zz_5431[26]}}, _zz_5431};
  assign _zz_5433 = fixTo_485_dout;
  assign _zz_5434 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_5435 = ($signed(_zz_408) - $signed(_zz_5436));
  assign _zz_5436 = ($signed(_zz_5437) * $signed(twiddle_factor_table_4_imag));
  assign _zz_5437 = ($signed(data_mid_2_37_real) + $signed(data_mid_2_37_imag));
  assign _zz_5438 = fixTo_486_dout;
  assign _zz_5439 = ($signed(_zz_408) + $signed(_zz_5440));
  assign _zz_5440 = ($signed(_zz_5441) * $signed(twiddle_factor_table_4_real));
  assign _zz_5441 = ($signed(data_mid_2_37_imag) - $signed(data_mid_2_37_real));
  assign _zz_5442 = fixTo_487_dout;
  assign _zz_5443 = _zz_5444[35 : 0];
  assign _zz_5444 = _zz_5445;
  assign _zz_5445 = ($signed(_zz_5446) >>> _zz_409);
  assign _zz_5446 = _zz_5447;
  assign _zz_5447 = ($signed(_zz_5449) - $signed(_zz_406));
  assign _zz_5448 = ({9'd0,data_mid_2_33_real} <<< 9);
  assign _zz_5449 = {{9{_zz_5448[26]}}, _zz_5448};
  assign _zz_5450 = fixTo_488_dout;
  assign _zz_5451 = _zz_5452[35 : 0];
  assign _zz_5452 = _zz_5453;
  assign _zz_5453 = ($signed(_zz_5454) >>> _zz_409);
  assign _zz_5454 = _zz_5455;
  assign _zz_5455 = ($signed(_zz_5457) - $signed(_zz_407));
  assign _zz_5456 = ({9'd0,data_mid_2_33_imag} <<< 9);
  assign _zz_5457 = {{9{_zz_5456[26]}}, _zz_5456};
  assign _zz_5458 = fixTo_489_dout;
  assign _zz_5459 = _zz_5460[35 : 0];
  assign _zz_5460 = _zz_5461;
  assign _zz_5461 = ($signed(_zz_5462) >>> _zz_410);
  assign _zz_5462 = _zz_5463;
  assign _zz_5463 = ($signed(_zz_5465) + $signed(_zz_406));
  assign _zz_5464 = ({9'd0,data_mid_2_33_real} <<< 9);
  assign _zz_5465 = {{9{_zz_5464[26]}}, _zz_5464};
  assign _zz_5466 = fixTo_490_dout;
  assign _zz_5467 = _zz_5468[35 : 0];
  assign _zz_5468 = _zz_5469;
  assign _zz_5469 = ($signed(_zz_5470) >>> _zz_410);
  assign _zz_5470 = _zz_5471;
  assign _zz_5471 = ($signed(_zz_5473) + $signed(_zz_407));
  assign _zz_5472 = ({9'd0,data_mid_2_33_imag} <<< 9);
  assign _zz_5473 = {{9{_zz_5472[26]}}, _zz_5472};
  assign _zz_5474 = fixTo_491_dout;
  assign _zz_5475 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_5476 = ($signed(_zz_413) - $signed(_zz_5477));
  assign _zz_5477 = ($signed(_zz_5478) * $signed(twiddle_factor_table_5_imag));
  assign _zz_5478 = ($signed(data_mid_2_38_real) + $signed(data_mid_2_38_imag));
  assign _zz_5479 = fixTo_492_dout;
  assign _zz_5480 = ($signed(_zz_413) + $signed(_zz_5481));
  assign _zz_5481 = ($signed(_zz_5482) * $signed(twiddle_factor_table_5_real));
  assign _zz_5482 = ($signed(data_mid_2_38_imag) - $signed(data_mid_2_38_real));
  assign _zz_5483 = fixTo_493_dout;
  assign _zz_5484 = _zz_5485[35 : 0];
  assign _zz_5485 = _zz_5486;
  assign _zz_5486 = ($signed(_zz_5487) >>> _zz_414);
  assign _zz_5487 = _zz_5488;
  assign _zz_5488 = ($signed(_zz_5490) - $signed(_zz_411));
  assign _zz_5489 = ({9'd0,data_mid_2_34_real} <<< 9);
  assign _zz_5490 = {{9{_zz_5489[26]}}, _zz_5489};
  assign _zz_5491 = fixTo_494_dout;
  assign _zz_5492 = _zz_5493[35 : 0];
  assign _zz_5493 = _zz_5494;
  assign _zz_5494 = ($signed(_zz_5495) >>> _zz_414);
  assign _zz_5495 = _zz_5496;
  assign _zz_5496 = ($signed(_zz_5498) - $signed(_zz_412));
  assign _zz_5497 = ({9'd0,data_mid_2_34_imag} <<< 9);
  assign _zz_5498 = {{9{_zz_5497[26]}}, _zz_5497};
  assign _zz_5499 = fixTo_495_dout;
  assign _zz_5500 = _zz_5501[35 : 0];
  assign _zz_5501 = _zz_5502;
  assign _zz_5502 = ($signed(_zz_5503) >>> _zz_415);
  assign _zz_5503 = _zz_5504;
  assign _zz_5504 = ($signed(_zz_5506) + $signed(_zz_411));
  assign _zz_5505 = ({9'd0,data_mid_2_34_real} <<< 9);
  assign _zz_5506 = {{9{_zz_5505[26]}}, _zz_5505};
  assign _zz_5507 = fixTo_496_dout;
  assign _zz_5508 = _zz_5509[35 : 0];
  assign _zz_5509 = _zz_5510;
  assign _zz_5510 = ($signed(_zz_5511) >>> _zz_415);
  assign _zz_5511 = _zz_5512;
  assign _zz_5512 = ($signed(_zz_5514) + $signed(_zz_412));
  assign _zz_5513 = ({9'd0,data_mid_2_34_imag} <<< 9);
  assign _zz_5514 = {{9{_zz_5513[26]}}, _zz_5513};
  assign _zz_5515 = fixTo_497_dout;
  assign _zz_5516 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_5517 = ($signed(_zz_418) - $signed(_zz_5518));
  assign _zz_5518 = ($signed(_zz_5519) * $signed(twiddle_factor_table_6_imag));
  assign _zz_5519 = ($signed(data_mid_2_39_real) + $signed(data_mid_2_39_imag));
  assign _zz_5520 = fixTo_498_dout;
  assign _zz_5521 = ($signed(_zz_418) + $signed(_zz_5522));
  assign _zz_5522 = ($signed(_zz_5523) * $signed(twiddle_factor_table_6_real));
  assign _zz_5523 = ($signed(data_mid_2_39_imag) - $signed(data_mid_2_39_real));
  assign _zz_5524 = fixTo_499_dout;
  assign _zz_5525 = _zz_5526[35 : 0];
  assign _zz_5526 = _zz_5527;
  assign _zz_5527 = ($signed(_zz_5528) >>> _zz_419);
  assign _zz_5528 = _zz_5529;
  assign _zz_5529 = ($signed(_zz_5531) - $signed(_zz_416));
  assign _zz_5530 = ({9'd0,data_mid_2_35_real} <<< 9);
  assign _zz_5531 = {{9{_zz_5530[26]}}, _zz_5530};
  assign _zz_5532 = fixTo_500_dout;
  assign _zz_5533 = _zz_5534[35 : 0];
  assign _zz_5534 = _zz_5535;
  assign _zz_5535 = ($signed(_zz_5536) >>> _zz_419);
  assign _zz_5536 = _zz_5537;
  assign _zz_5537 = ($signed(_zz_5539) - $signed(_zz_417));
  assign _zz_5538 = ({9'd0,data_mid_2_35_imag} <<< 9);
  assign _zz_5539 = {{9{_zz_5538[26]}}, _zz_5538};
  assign _zz_5540 = fixTo_501_dout;
  assign _zz_5541 = _zz_5542[35 : 0];
  assign _zz_5542 = _zz_5543;
  assign _zz_5543 = ($signed(_zz_5544) >>> _zz_420);
  assign _zz_5544 = _zz_5545;
  assign _zz_5545 = ($signed(_zz_5547) + $signed(_zz_416));
  assign _zz_5546 = ({9'd0,data_mid_2_35_real} <<< 9);
  assign _zz_5547 = {{9{_zz_5546[26]}}, _zz_5546};
  assign _zz_5548 = fixTo_502_dout;
  assign _zz_5549 = _zz_5550[35 : 0];
  assign _zz_5550 = _zz_5551;
  assign _zz_5551 = ($signed(_zz_5552) >>> _zz_420);
  assign _zz_5552 = _zz_5553;
  assign _zz_5553 = ($signed(_zz_5555) + $signed(_zz_417));
  assign _zz_5554 = ({9'd0,data_mid_2_35_imag} <<< 9);
  assign _zz_5555 = {{9{_zz_5554[26]}}, _zz_5554};
  assign _zz_5556 = fixTo_503_dout;
  assign _zz_5557 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_5558 = ($signed(_zz_423) - $signed(_zz_5559));
  assign _zz_5559 = ($signed(_zz_5560) * $signed(twiddle_factor_table_3_imag));
  assign _zz_5560 = ($signed(data_mid_2_44_real) + $signed(data_mid_2_44_imag));
  assign _zz_5561 = fixTo_504_dout;
  assign _zz_5562 = ($signed(_zz_423) + $signed(_zz_5563));
  assign _zz_5563 = ($signed(_zz_5564) * $signed(twiddle_factor_table_3_real));
  assign _zz_5564 = ($signed(data_mid_2_44_imag) - $signed(data_mid_2_44_real));
  assign _zz_5565 = fixTo_505_dout;
  assign _zz_5566 = _zz_5567[35 : 0];
  assign _zz_5567 = _zz_5568;
  assign _zz_5568 = ($signed(_zz_5569) >>> _zz_424);
  assign _zz_5569 = _zz_5570;
  assign _zz_5570 = ($signed(_zz_5572) - $signed(_zz_421));
  assign _zz_5571 = ({9'd0,data_mid_2_40_real} <<< 9);
  assign _zz_5572 = {{9{_zz_5571[26]}}, _zz_5571};
  assign _zz_5573 = fixTo_506_dout;
  assign _zz_5574 = _zz_5575[35 : 0];
  assign _zz_5575 = _zz_5576;
  assign _zz_5576 = ($signed(_zz_5577) >>> _zz_424);
  assign _zz_5577 = _zz_5578;
  assign _zz_5578 = ($signed(_zz_5580) - $signed(_zz_422));
  assign _zz_5579 = ({9'd0,data_mid_2_40_imag} <<< 9);
  assign _zz_5580 = {{9{_zz_5579[26]}}, _zz_5579};
  assign _zz_5581 = fixTo_507_dout;
  assign _zz_5582 = _zz_5583[35 : 0];
  assign _zz_5583 = _zz_5584;
  assign _zz_5584 = ($signed(_zz_5585) >>> _zz_425);
  assign _zz_5585 = _zz_5586;
  assign _zz_5586 = ($signed(_zz_5588) + $signed(_zz_421));
  assign _zz_5587 = ({9'd0,data_mid_2_40_real} <<< 9);
  assign _zz_5588 = {{9{_zz_5587[26]}}, _zz_5587};
  assign _zz_5589 = fixTo_508_dout;
  assign _zz_5590 = _zz_5591[35 : 0];
  assign _zz_5591 = _zz_5592;
  assign _zz_5592 = ($signed(_zz_5593) >>> _zz_425);
  assign _zz_5593 = _zz_5594;
  assign _zz_5594 = ($signed(_zz_5596) + $signed(_zz_422));
  assign _zz_5595 = ({9'd0,data_mid_2_40_imag} <<< 9);
  assign _zz_5596 = {{9{_zz_5595[26]}}, _zz_5595};
  assign _zz_5597 = fixTo_509_dout;
  assign _zz_5598 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_5599 = ($signed(_zz_428) - $signed(_zz_5600));
  assign _zz_5600 = ($signed(_zz_5601) * $signed(twiddle_factor_table_4_imag));
  assign _zz_5601 = ($signed(data_mid_2_45_real) + $signed(data_mid_2_45_imag));
  assign _zz_5602 = fixTo_510_dout;
  assign _zz_5603 = ($signed(_zz_428) + $signed(_zz_5604));
  assign _zz_5604 = ($signed(_zz_5605) * $signed(twiddle_factor_table_4_real));
  assign _zz_5605 = ($signed(data_mid_2_45_imag) - $signed(data_mid_2_45_real));
  assign _zz_5606 = fixTo_511_dout;
  assign _zz_5607 = _zz_5608[35 : 0];
  assign _zz_5608 = _zz_5609;
  assign _zz_5609 = ($signed(_zz_5610) >>> _zz_429);
  assign _zz_5610 = _zz_5611;
  assign _zz_5611 = ($signed(_zz_5613) - $signed(_zz_426));
  assign _zz_5612 = ({9'd0,data_mid_2_41_real} <<< 9);
  assign _zz_5613 = {{9{_zz_5612[26]}}, _zz_5612};
  assign _zz_5614 = fixTo_512_dout;
  assign _zz_5615 = _zz_5616[35 : 0];
  assign _zz_5616 = _zz_5617;
  assign _zz_5617 = ($signed(_zz_5618) >>> _zz_429);
  assign _zz_5618 = _zz_5619;
  assign _zz_5619 = ($signed(_zz_5621) - $signed(_zz_427));
  assign _zz_5620 = ({9'd0,data_mid_2_41_imag} <<< 9);
  assign _zz_5621 = {{9{_zz_5620[26]}}, _zz_5620};
  assign _zz_5622 = fixTo_513_dout;
  assign _zz_5623 = _zz_5624[35 : 0];
  assign _zz_5624 = _zz_5625;
  assign _zz_5625 = ($signed(_zz_5626) >>> _zz_430);
  assign _zz_5626 = _zz_5627;
  assign _zz_5627 = ($signed(_zz_5629) + $signed(_zz_426));
  assign _zz_5628 = ({9'd0,data_mid_2_41_real} <<< 9);
  assign _zz_5629 = {{9{_zz_5628[26]}}, _zz_5628};
  assign _zz_5630 = fixTo_514_dout;
  assign _zz_5631 = _zz_5632[35 : 0];
  assign _zz_5632 = _zz_5633;
  assign _zz_5633 = ($signed(_zz_5634) >>> _zz_430);
  assign _zz_5634 = _zz_5635;
  assign _zz_5635 = ($signed(_zz_5637) + $signed(_zz_427));
  assign _zz_5636 = ({9'd0,data_mid_2_41_imag} <<< 9);
  assign _zz_5637 = {{9{_zz_5636[26]}}, _zz_5636};
  assign _zz_5638 = fixTo_515_dout;
  assign _zz_5639 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_5640 = ($signed(_zz_433) - $signed(_zz_5641));
  assign _zz_5641 = ($signed(_zz_5642) * $signed(twiddle_factor_table_5_imag));
  assign _zz_5642 = ($signed(data_mid_2_46_real) + $signed(data_mid_2_46_imag));
  assign _zz_5643 = fixTo_516_dout;
  assign _zz_5644 = ($signed(_zz_433) + $signed(_zz_5645));
  assign _zz_5645 = ($signed(_zz_5646) * $signed(twiddle_factor_table_5_real));
  assign _zz_5646 = ($signed(data_mid_2_46_imag) - $signed(data_mid_2_46_real));
  assign _zz_5647 = fixTo_517_dout;
  assign _zz_5648 = _zz_5649[35 : 0];
  assign _zz_5649 = _zz_5650;
  assign _zz_5650 = ($signed(_zz_5651) >>> _zz_434);
  assign _zz_5651 = _zz_5652;
  assign _zz_5652 = ($signed(_zz_5654) - $signed(_zz_431));
  assign _zz_5653 = ({9'd0,data_mid_2_42_real} <<< 9);
  assign _zz_5654 = {{9{_zz_5653[26]}}, _zz_5653};
  assign _zz_5655 = fixTo_518_dout;
  assign _zz_5656 = _zz_5657[35 : 0];
  assign _zz_5657 = _zz_5658;
  assign _zz_5658 = ($signed(_zz_5659) >>> _zz_434);
  assign _zz_5659 = _zz_5660;
  assign _zz_5660 = ($signed(_zz_5662) - $signed(_zz_432));
  assign _zz_5661 = ({9'd0,data_mid_2_42_imag} <<< 9);
  assign _zz_5662 = {{9{_zz_5661[26]}}, _zz_5661};
  assign _zz_5663 = fixTo_519_dout;
  assign _zz_5664 = _zz_5665[35 : 0];
  assign _zz_5665 = _zz_5666;
  assign _zz_5666 = ($signed(_zz_5667) >>> _zz_435);
  assign _zz_5667 = _zz_5668;
  assign _zz_5668 = ($signed(_zz_5670) + $signed(_zz_431));
  assign _zz_5669 = ({9'd0,data_mid_2_42_real} <<< 9);
  assign _zz_5670 = {{9{_zz_5669[26]}}, _zz_5669};
  assign _zz_5671 = fixTo_520_dout;
  assign _zz_5672 = _zz_5673[35 : 0];
  assign _zz_5673 = _zz_5674;
  assign _zz_5674 = ($signed(_zz_5675) >>> _zz_435);
  assign _zz_5675 = _zz_5676;
  assign _zz_5676 = ($signed(_zz_5678) + $signed(_zz_432));
  assign _zz_5677 = ({9'd0,data_mid_2_42_imag} <<< 9);
  assign _zz_5678 = {{9{_zz_5677[26]}}, _zz_5677};
  assign _zz_5679 = fixTo_521_dout;
  assign _zz_5680 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_5681 = ($signed(_zz_438) - $signed(_zz_5682));
  assign _zz_5682 = ($signed(_zz_5683) * $signed(twiddle_factor_table_6_imag));
  assign _zz_5683 = ($signed(data_mid_2_47_real) + $signed(data_mid_2_47_imag));
  assign _zz_5684 = fixTo_522_dout;
  assign _zz_5685 = ($signed(_zz_438) + $signed(_zz_5686));
  assign _zz_5686 = ($signed(_zz_5687) * $signed(twiddle_factor_table_6_real));
  assign _zz_5687 = ($signed(data_mid_2_47_imag) - $signed(data_mid_2_47_real));
  assign _zz_5688 = fixTo_523_dout;
  assign _zz_5689 = _zz_5690[35 : 0];
  assign _zz_5690 = _zz_5691;
  assign _zz_5691 = ($signed(_zz_5692) >>> _zz_439);
  assign _zz_5692 = _zz_5693;
  assign _zz_5693 = ($signed(_zz_5695) - $signed(_zz_436));
  assign _zz_5694 = ({9'd0,data_mid_2_43_real} <<< 9);
  assign _zz_5695 = {{9{_zz_5694[26]}}, _zz_5694};
  assign _zz_5696 = fixTo_524_dout;
  assign _zz_5697 = _zz_5698[35 : 0];
  assign _zz_5698 = _zz_5699;
  assign _zz_5699 = ($signed(_zz_5700) >>> _zz_439);
  assign _zz_5700 = _zz_5701;
  assign _zz_5701 = ($signed(_zz_5703) - $signed(_zz_437));
  assign _zz_5702 = ({9'd0,data_mid_2_43_imag} <<< 9);
  assign _zz_5703 = {{9{_zz_5702[26]}}, _zz_5702};
  assign _zz_5704 = fixTo_525_dout;
  assign _zz_5705 = _zz_5706[35 : 0];
  assign _zz_5706 = _zz_5707;
  assign _zz_5707 = ($signed(_zz_5708) >>> _zz_440);
  assign _zz_5708 = _zz_5709;
  assign _zz_5709 = ($signed(_zz_5711) + $signed(_zz_436));
  assign _zz_5710 = ({9'd0,data_mid_2_43_real} <<< 9);
  assign _zz_5711 = {{9{_zz_5710[26]}}, _zz_5710};
  assign _zz_5712 = fixTo_526_dout;
  assign _zz_5713 = _zz_5714[35 : 0];
  assign _zz_5714 = _zz_5715;
  assign _zz_5715 = ($signed(_zz_5716) >>> _zz_440);
  assign _zz_5716 = _zz_5717;
  assign _zz_5717 = ($signed(_zz_5719) + $signed(_zz_437));
  assign _zz_5718 = ({9'd0,data_mid_2_43_imag} <<< 9);
  assign _zz_5719 = {{9{_zz_5718[26]}}, _zz_5718};
  assign _zz_5720 = fixTo_527_dout;
  assign _zz_5721 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_5722 = ($signed(_zz_443) - $signed(_zz_5723));
  assign _zz_5723 = ($signed(_zz_5724) * $signed(twiddle_factor_table_3_imag));
  assign _zz_5724 = ($signed(data_mid_2_52_real) + $signed(data_mid_2_52_imag));
  assign _zz_5725 = fixTo_528_dout;
  assign _zz_5726 = ($signed(_zz_443) + $signed(_zz_5727));
  assign _zz_5727 = ($signed(_zz_5728) * $signed(twiddle_factor_table_3_real));
  assign _zz_5728 = ($signed(data_mid_2_52_imag) - $signed(data_mid_2_52_real));
  assign _zz_5729 = fixTo_529_dout;
  assign _zz_5730 = _zz_5731[35 : 0];
  assign _zz_5731 = _zz_5732;
  assign _zz_5732 = ($signed(_zz_5733) >>> _zz_444);
  assign _zz_5733 = _zz_5734;
  assign _zz_5734 = ($signed(_zz_5736) - $signed(_zz_441));
  assign _zz_5735 = ({9'd0,data_mid_2_48_real} <<< 9);
  assign _zz_5736 = {{9{_zz_5735[26]}}, _zz_5735};
  assign _zz_5737 = fixTo_530_dout;
  assign _zz_5738 = _zz_5739[35 : 0];
  assign _zz_5739 = _zz_5740;
  assign _zz_5740 = ($signed(_zz_5741) >>> _zz_444);
  assign _zz_5741 = _zz_5742;
  assign _zz_5742 = ($signed(_zz_5744) - $signed(_zz_442));
  assign _zz_5743 = ({9'd0,data_mid_2_48_imag} <<< 9);
  assign _zz_5744 = {{9{_zz_5743[26]}}, _zz_5743};
  assign _zz_5745 = fixTo_531_dout;
  assign _zz_5746 = _zz_5747[35 : 0];
  assign _zz_5747 = _zz_5748;
  assign _zz_5748 = ($signed(_zz_5749) >>> _zz_445);
  assign _zz_5749 = _zz_5750;
  assign _zz_5750 = ($signed(_zz_5752) + $signed(_zz_441));
  assign _zz_5751 = ({9'd0,data_mid_2_48_real} <<< 9);
  assign _zz_5752 = {{9{_zz_5751[26]}}, _zz_5751};
  assign _zz_5753 = fixTo_532_dout;
  assign _zz_5754 = _zz_5755[35 : 0];
  assign _zz_5755 = _zz_5756;
  assign _zz_5756 = ($signed(_zz_5757) >>> _zz_445);
  assign _zz_5757 = _zz_5758;
  assign _zz_5758 = ($signed(_zz_5760) + $signed(_zz_442));
  assign _zz_5759 = ({9'd0,data_mid_2_48_imag} <<< 9);
  assign _zz_5760 = {{9{_zz_5759[26]}}, _zz_5759};
  assign _zz_5761 = fixTo_533_dout;
  assign _zz_5762 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_5763 = ($signed(_zz_448) - $signed(_zz_5764));
  assign _zz_5764 = ($signed(_zz_5765) * $signed(twiddle_factor_table_4_imag));
  assign _zz_5765 = ($signed(data_mid_2_53_real) + $signed(data_mid_2_53_imag));
  assign _zz_5766 = fixTo_534_dout;
  assign _zz_5767 = ($signed(_zz_448) + $signed(_zz_5768));
  assign _zz_5768 = ($signed(_zz_5769) * $signed(twiddle_factor_table_4_real));
  assign _zz_5769 = ($signed(data_mid_2_53_imag) - $signed(data_mid_2_53_real));
  assign _zz_5770 = fixTo_535_dout;
  assign _zz_5771 = _zz_5772[35 : 0];
  assign _zz_5772 = _zz_5773;
  assign _zz_5773 = ($signed(_zz_5774) >>> _zz_449);
  assign _zz_5774 = _zz_5775;
  assign _zz_5775 = ($signed(_zz_5777) - $signed(_zz_446));
  assign _zz_5776 = ({9'd0,data_mid_2_49_real} <<< 9);
  assign _zz_5777 = {{9{_zz_5776[26]}}, _zz_5776};
  assign _zz_5778 = fixTo_536_dout;
  assign _zz_5779 = _zz_5780[35 : 0];
  assign _zz_5780 = _zz_5781;
  assign _zz_5781 = ($signed(_zz_5782) >>> _zz_449);
  assign _zz_5782 = _zz_5783;
  assign _zz_5783 = ($signed(_zz_5785) - $signed(_zz_447));
  assign _zz_5784 = ({9'd0,data_mid_2_49_imag} <<< 9);
  assign _zz_5785 = {{9{_zz_5784[26]}}, _zz_5784};
  assign _zz_5786 = fixTo_537_dout;
  assign _zz_5787 = _zz_5788[35 : 0];
  assign _zz_5788 = _zz_5789;
  assign _zz_5789 = ($signed(_zz_5790) >>> _zz_450);
  assign _zz_5790 = _zz_5791;
  assign _zz_5791 = ($signed(_zz_5793) + $signed(_zz_446));
  assign _zz_5792 = ({9'd0,data_mid_2_49_real} <<< 9);
  assign _zz_5793 = {{9{_zz_5792[26]}}, _zz_5792};
  assign _zz_5794 = fixTo_538_dout;
  assign _zz_5795 = _zz_5796[35 : 0];
  assign _zz_5796 = _zz_5797;
  assign _zz_5797 = ($signed(_zz_5798) >>> _zz_450);
  assign _zz_5798 = _zz_5799;
  assign _zz_5799 = ($signed(_zz_5801) + $signed(_zz_447));
  assign _zz_5800 = ({9'd0,data_mid_2_49_imag} <<< 9);
  assign _zz_5801 = {{9{_zz_5800[26]}}, _zz_5800};
  assign _zz_5802 = fixTo_539_dout;
  assign _zz_5803 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_5804 = ($signed(_zz_453) - $signed(_zz_5805));
  assign _zz_5805 = ($signed(_zz_5806) * $signed(twiddle_factor_table_5_imag));
  assign _zz_5806 = ($signed(data_mid_2_54_real) + $signed(data_mid_2_54_imag));
  assign _zz_5807 = fixTo_540_dout;
  assign _zz_5808 = ($signed(_zz_453) + $signed(_zz_5809));
  assign _zz_5809 = ($signed(_zz_5810) * $signed(twiddle_factor_table_5_real));
  assign _zz_5810 = ($signed(data_mid_2_54_imag) - $signed(data_mid_2_54_real));
  assign _zz_5811 = fixTo_541_dout;
  assign _zz_5812 = _zz_5813[35 : 0];
  assign _zz_5813 = _zz_5814;
  assign _zz_5814 = ($signed(_zz_5815) >>> _zz_454);
  assign _zz_5815 = _zz_5816;
  assign _zz_5816 = ($signed(_zz_5818) - $signed(_zz_451));
  assign _zz_5817 = ({9'd0,data_mid_2_50_real} <<< 9);
  assign _zz_5818 = {{9{_zz_5817[26]}}, _zz_5817};
  assign _zz_5819 = fixTo_542_dout;
  assign _zz_5820 = _zz_5821[35 : 0];
  assign _zz_5821 = _zz_5822;
  assign _zz_5822 = ($signed(_zz_5823) >>> _zz_454);
  assign _zz_5823 = _zz_5824;
  assign _zz_5824 = ($signed(_zz_5826) - $signed(_zz_452));
  assign _zz_5825 = ({9'd0,data_mid_2_50_imag} <<< 9);
  assign _zz_5826 = {{9{_zz_5825[26]}}, _zz_5825};
  assign _zz_5827 = fixTo_543_dout;
  assign _zz_5828 = _zz_5829[35 : 0];
  assign _zz_5829 = _zz_5830;
  assign _zz_5830 = ($signed(_zz_5831) >>> _zz_455);
  assign _zz_5831 = _zz_5832;
  assign _zz_5832 = ($signed(_zz_5834) + $signed(_zz_451));
  assign _zz_5833 = ({9'd0,data_mid_2_50_real} <<< 9);
  assign _zz_5834 = {{9{_zz_5833[26]}}, _zz_5833};
  assign _zz_5835 = fixTo_544_dout;
  assign _zz_5836 = _zz_5837[35 : 0];
  assign _zz_5837 = _zz_5838;
  assign _zz_5838 = ($signed(_zz_5839) >>> _zz_455);
  assign _zz_5839 = _zz_5840;
  assign _zz_5840 = ($signed(_zz_5842) + $signed(_zz_452));
  assign _zz_5841 = ({9'd0,data_mid_2_50_imag} <<< 9);
  assign _zz_5842 = {{9{_zz_5841[26]}}, _zz_5841};
  assign _zz_5843 = fixTo_545_dout;
  assign _zz_5844 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_5845 = ($signed(_zz_458) - $signed(_zz_5846));
  assign _zz_5846 = ($signed(_zz_5847) * $signed(twiddle_factor_table_6_imag));
  assign _zz_5847 = ($signed(data_mid_2_55_real) + $signed(data_mid_2_55_imag));
  assign _zz_5848 = fixTo_546_dout;
  assign _zz_5849 = ($signed(_zz_458) + $signed(_zz_5850));
  assign _zz_5850 = ($signed(_zz_5851) * $signed(twiddle_factor_table_6_real));
  assign _zz_5851 = ($signed(data_mid_2_55_imag) - $signed(data_mid_2_55_real));
  assign _zz_5852 = fixTo_547_dout;
  assign _zz_5853 = _zz_5854[35 : 0];
  assign _zz_5854 = _zz_5855;
  assign _zz_5855 = ($signed(_zz_5856) >>> _zz_459);
  assign _zz_5856 = _zz_5857;
  assign _zz_5857 = ($signed(_zz_5859) - $signed(_zz_456));
  assign _zz_5858 = ({9'd0,data_mid_2_51_real} <<< 9);
  assign _zz_5859 = {{9{_zz_5858[26]}}, _zz_5858};
  assign _zz_5860 = fixTo_548_dout;
  assign _zz_5861 = _zz_5862[35 : 0];
  assign _zz_5862 = _zz_5863;
  assign _zz_5863 = ($signed(_zz_5864) >>> _zz_459);
  assign _zz_5864 = _zz_5865;
  assign _zz_5865 = ($signed(_zz_5867) - $signed(_zz_457));
  assign _zz_5866 = ({9'd0,data_mid_2_51_imag} <<< 9);
  assign _zz_5867 = {{9{_zz_5866[26]}}, _zz_5866};
  assign _zz_5868 = fixTo_549_dout;
  assign _zz_5869 = _zz_5870[35 : 0];
  assign _zz_5870 = _zz_5871;
  assign _zz_5871 = ($signed(_zz_5872) >>> _zz_460);
  assign _zz_5872 = _zz_5873;
  assign _zz_5873 = ($signed(_zz_5875) + $signed(_zz_456));
  assign _zz_5874 = ({9'd0,data_mid_2_51_real} <<< 9);
  assign _zz_5875 = {{9{_zz_5874[26]}}, _zz_5874};
  assign _zz_5876 = fixTo_550_dout;
  assign _zz_5877 = _zz_5878[35 : 0];
  assign _zz_5878 = _zz_5879;
  assign _zz_5879 = ($signed(_zz_5880) >>> _zz_460);
  assign _zz_5880 = _zz_5881;
  assign _zz_5881 = ($signed(_zz_5883) + $signed(_zz_457));
  assign _zz_5882 = ({9'd0,data_mid_2_51_imag} <<< 9);
  assign _zz_5883 = {{9{_zz_5882[26]}}, _zz_5882};
  assign _zz_5884 = fixTo_551_dout;
  assign _zz_5885 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_5886 = ($signed(_zz_463) - $signed(_zz_5887));
  assign _zz_5887 = ($signed(_zz_5888) * $signed(twiddle_factor_table_3_imag));
  assign _zz_5888 = ($signed(data_mid_2_60_real) + $signed(data_mid_2_60_imag));
  assign _zz_5889 = fixTo_552_dout;
  assign _zz_5890 = ($signed(_zz_463) + $signed(_zz_5891));
  assign _zz_5891 = ($signed(_zz_5892) * $signed(twiddle_factor_table_3_real));
  assign _zz_5892 = ($signed(data_mid_2_60_imag) - $signed(data_mid_2_60_real));
  assign _zz_5893 = fixTo_553_dout;
  assign _zz_5894 = _zz_5895[35 : 0];
  assign _zz_5895 = _zz_5896;
  assign _zz_5896 = ($signed(_zz_5897) >>> _zz_464);
  assign _zz_5897 = _zz_5898;
  assign _zz_5898 = ($signed(_zz_5900) - $signed(_zz_461));
  assign _zz_5899 = ({9'd0,data_mid_2_56_real} <<< 9);
  assign _zz_5900 = {{9{_zz_5899[26]}}, _zz_5899};
  assign _zz_5901 = fixTo_554_dout;
  assign _zz_5902 = _zz_5903[35 : 0];
  assign _zz_5903 = _zz_5904;
  assign _zz_5904 = ($signed(_zz_5905) >>> _zz_464);
  assign _zz_5905 = _zz_5906;
  assign _zz_5906 = ($signed(_zz_5908) - $signed(_zz_462));
  assign _zz_5907 = ({9'd0,data_mid_2_56_imag} <<< 9);
  assign _zz_5908 = {{9{_zz_5907[26]}}, _zz_5907};
  assign _zz_5909 = fixTo_555_dout;
  assign _zz_5910 = _zz_5911[35 : 0];
  assign _zz_5911 = _zz_5912;
  assign _zz_5912 = ($signed(_zz_5913) >>> _zz_465);
  assign _zz_5913 = _zz_5914;
  assign _zz_5914 = ($signed(_zz_5916) + $signed(_zz_461));
  assign _zz_5915 = ({9'd0,data_mid_2_56_real} <<< 9);
  assign _zz_5916 = {{9{_zz_5915[26]}}, _zz_5915};
  assign _zz_5917 = fixTo_556_dout;
  assign _zz_5918 = _zz_5919[35 : 0];
  assign _zz_5919 = _zz_5920;
  assign _zz_5920 = ($signed(_zz_5921) >>> _zz_465);
  assign _zz_5921 = _zz_5922;
  assign _zz_5922 = ($signed(_zz_5924) + $signed(_zz_462));
  assign _zz_5923 = ({9'd0,data_mid_2_56_imag} <<< 9);
  assign _zz_5924 = {{9{_zz_5923[26]}}, _zz_5923};
  assign _zz_5925 = fixTo_557_dout;
  assign _zz_5926 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_5927 = ($signed(_zz_468) - $signed(_zz_5928));
  assign _zz_5928 = ($signed(_zz_5929) * $signed(twiddle_factor_table_4_imag));
  assign _zz_5929 = ($signed(data_mid_2_61_real) + $signed(data_mid_2_61_imag));
  assign _zz_5930 = fixTo_558_dout;
  assign _zz_5931 = ($signed(_zz_468) + $signed(_zz_5932));
  assign _zz_5932 = ($signed(_zz_5933) * $signed(twiddle_factor_table_4_real));
  assign _zz_5933 = ($signed(data_mid_2_61_imag) - $signed(data_mid_2_61_real));
  assign _zz_5934 = fixTo_559_dout;
  assign _zz_5935 = _zz_5936[35 : 0];
  assign _zz_5936 = _zz_5937;
  assign _zz_5937 = ($signed(_zz_5938) >>> _zz_469);
  assign _zz_5938 = _zz_5939;
  assign _zz_5939 = ($signed(_zz_5941) - $signed(_zz_466));
  assign _zz_5940 = ({9'd0,data_mid_2_57_real} <<< 9);
  assign _zz_5941 = {{9{_zz_5940[26]}}, _zz_5940};
  assign _zz_5942 = fixTo_560_dout;
  assign _zz_5943 = _zz_5944[35 : 0];
  assign _zz_5944 = _zz_5945;
  assign _zz_5945 = ($signed(_zz_5946) >>> _zz_469);
  assign _zz_5946 = _zz_5947;
  assign _zz_5947 = ($signed(_zz_5949) - $signed(_zz_467));
  assign _zz_5948 = ({9'd0,data_mid_2_57_imag} <<< 9);
  assign _zz_5949 = {{9{_zz_5948[26]}}, _zz_5948};
  assign _zz_5950 = fixTo_561_dout;
  assign _zz_5951 = _zz_5952[35 : 0];
  assign _zz_5952 = _zz_5953;
  assign _zz_5953 = ($signed(_zz_5954) >>> _zz_470);
  assign _zz_5954 = _zz_5955;
  assign _zz_5955 = ($signed(_zz_5957) + $signed(_zz_466));
  assign _zz_5956 = ({9'd0,data_mid_2_57_real} <<< 9);
  assign _zz_5957 = {{9{_zz_5956[26]}}, _zz_5956};
  assign _zz_5958 = fixTo_562_dout;
  assign _zz_5959 = _zz_5960[35 : 0];
  assign _zz_5960 = _zz_5961;
  assign _zz_5961 = ($signed(_zz_5962) >>> _zz_470);
  assign _zz_5962 = _zz_5963;
  assign _zz_5963 = ($signed(_zz_5965) + $signed(_zz_467));
  assign _zz_5964 = ({9'd0,data_mid_2_57_imag} <<< 9);
  assign _zz_5965 = {{9{_zz_5964[26]}}, _zz_5964};
  assign _zz_5966 = fixTo_563_dout;
  assign _zz_5967 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_5968 = ($signed(_zz_473) - $signed(_zz_5969));
  assign _zz_5969 = ($signed(_zz_5970) * $signed(twiddle_factor_table_5_imag));
  assign _zz_5970 = ($signed(data_mid_2_62_real) + $signed(data_mid_2_62_imag));
  assign _zz_5971 = fixTo_564_dout;
  assign _zz_5972 = ($signed(_zz_473) + $signed(_zz_5973));
  assign _zz_5973 = ($signed(_zz_5974) * $signed(twiddle_factor_table_5_real));
  assign _zz_5974 = ($signed(data_mid_2_62_imag) - $signed(data_mid_2_62_real));
  assign _zz_5975 = fixTo_565_dout;
  assign _zz_5976 = _zz_5977[35 : 0];
  assign _zz_5977 = _zz_5978;
  assign _zz_5978 = ($signed(_zz_5979) >>> _zz_474);
  assign _zz_5979 = _zz_5980;
  assign _zz_5980 = ($signed(_zz_5982) - $signed(_zz_471));
  assign _zz_5981 = ({9'd0,data_mid_2_58_real} <<< 9);
  assign _zz_5982 = {{9{_zz_5981[26]}}, _zz_5981};
  assign _zz_5983 = fixTo_566_dout;
  assign _zz_5984 = _zz_5985[35 : 0];
  assign _zz_5985 = _zz_5986;
  assign _zz_5986 = ($signed(_zz_5987) >>> _zz_474);
  assign _zz_5987 = _zz_5988;
  assign _zz_5988 = ($signed(_zz_5990) - $signed(_zz_472));
  assign _zz_5989 = ({9'd0,data_mid_2_58_imag} <<< 9);
  assign _zz_5990 = {{9{_zz_5989[26]}}, _zz_5989};
  assign _zz_5991 = fixTo_567_dout;
  assign _zz_5992 = _zz_5993[35 : 0];
  assign _zz_5993 = _zz_5994;
  assign _zz_5994 = ($signed(_zz_5995) >>> _zz_475);
  assign _zz_5995 = _zz_5996;
  assign _zz_5996 = ($signed(_zz_5998) + $signed(_zz_471));
  assign _zz_5997 = ({9'd0,data_mid_2_58_real} <<< 9);
  assign _zz_5998 = {{9{_zz_5997[26]}}, _zz_5997};
  assign _zz_5999 = fixTo_568_dout;
  assign _zz_6000 = _zz_6001[35 : 0];
  assign _zz_6001 = _zz_6002;
  assign _zz_6002 = ($signed(_zz_6003) >>> _zz_475);
  assign _zz_6003 = _zz_6004;
  assign _zz_6004 = ($signed(_zz_6006) + $signed(_zz_472));
  assign _zz_6005 = ({9'd0,data_mid_2_58_imag} <<< 9);
  assign _zz_6006 = {{9{_zz_6005[26]}}, _zz_6005};
  assign _zz_6007 = fixTo_569_dout;
  assign _zz_6008 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_6009 = ($signed(_zz_478) - $signed(_zz_6010));
  assign _zz_6010 = ($signed(_zz_6011) * $signed(twiddle_factor_table_6_imag));
  assign _zz_6011 = ($signed(data_mid_2_63_real) + $signed(data_mid_2_63_imag));
  assign _zz_6012 = fixTo_570_dout;
  assign _zz_6013 = ($signed(_zz_478) + $signed(_zz_6014));
  assign _zz_6014 = ($signed(_zz_6015) * $signed(twiddle_factor_table_6_real));
  assign _zz_6015 = ($signed(data_mid_2_63_imag) - $signed(data_mid_2_63_real));
  assign _zz_6016 = fixTo_571_dout;
  assign _zz_6017 = _zz_6018[35 : 0];
  assign _zz_6018 = _zz_6019;
  assign _zz_6019 = ($signed(_zz_6020) >>> _zz_479);
  assign _zz_6020 = _zz_6021;
  assign _zz_6021 = ($signed(_zz_6023) - $signed(_zz_476));
  assign _zz_6022 = ({9'd0,data_mid_2_59_real} <<< 9);
  assign _zz_6023 = {{9{_zz_6022[26]}}, _zz_6022};
  assign _zz_6024 = fixTo_572_dout;
  assign _zz_6025 = _zz_6026[35 : 0];
  assign _zz_6026 = _zz_6027;
  assign _zz_6027 = ($signed(_zz_6028) >>> _zz_479);
  assign _zz_6028 = _zz_6029;
  assign _zz_6029 = ($signed(_zz_6031) - $signed(_zz_477));
  assign _zz_6030 = ({9'd0,data_mid_2_59_imag} <<< 9);
  assign _zz_6031 = {{9{_zz_6030[26]}}, _zz_6030};
  assign _zz_6032 = fixTo_573_dout;
  assign _zz_6033 = _zz_6034[35 : 0];
  assign _zz_6034 = _zz_6035;
  assign _zz_6035 = ($signed(_zz_6036) >>> _zz_480);
  assign _zz_6036 = _zz_6037;
  assign _zz_6037 = ($signed(_zz_6039) + $signed(_zz_476));
  assign _zz_6038 = ({9'd0,data_mid_2_59_real} <<< 9);
  assign _zz_6039 = {{9{_zz_6038[26]}}, _zz_6038};
  assign _zz_6040 = fixTo_574_dout;
  assign _zz_6041 = _zz_6042[35 : 0];
  assign _zz_6042 = _zz_6043;
  assign _zz_6043 = ($signed(_zz_6044) >>> _zz_480);
  assign _zz_6044 = _zz_6045;
  assign _zz_6045 = ($signed(_zz_6047) + $signed(_zz_477));
  assign _zz_6046 = ({9'd0,data_mid_2_59_imag} <<< 9);
  assign _zz_6047 = {{9{_zz_6046[26]}}, _zz_6046};
  assign _zz_6048 = fixTo_575_dout;
  assign _zz_6049 = ($signed(twiddle_factor_table_7_real) + $signed(twiddle_factor_table_7_imag));
  assign _zz_6050 = ($signed(_zz_483) - $signed(_zz_6051));
  assign _zz_6051 = ($signed(_zz_6052) * $signed(twiddle_factor_table_7_imag));
  assign _zz_6052 = ($signed(data_mid_3_8_real) + $signed(data_mid_3_8_imag));
  assign _zz_6053 = fixTo_576_dout;
  assign _zz_6054 = ($signed(_zz_483) + $signed(_zz_6055));
  assign _zz_6055 = ($signed(_zz_6056) * $signed(twiddle_factor_table_7_real));
  assign _zz_6056 = ($signed(data_mid_3_8_imag) - $signed(data_mid_3_8_real));
  assign _zz_6057 = fixTo_577_dout;
  assign _zz_6058 = _zz_6059[35 : 0];
  assign _zz_6059 = _zz_6060;
  assign _zz_6060 = ($signed(_zz_6061) >>> _zz_484);
  assign _zz_6061 = _zz_6062;
  assign _zz_6062 = ($signed(_zz_6064) - $signed(_zz_481));
  assign _zz_6063 = ({9'd0,data_mid_3_0_real} <<< 9);
  assign _zz_6064 = {{9{_zz_6063[26]}}, _zz_6063};
  assign _zz_6065 = fixTo_578_dout;
  assign _zz_6066 = _zz_6067[35 : 0];
  assign _zz_6067 = _zz_6068;
  assign _zz_6068 = ($signed(_zz_6069) >>> _zz_484);
  assign _zz_6069 = _zz_6070;
  assign _zz_6070 = ($signed(_zz_6072) - $signed(_zz_482));
  assign _zz_6071 = ({9'd0,data_mid_3_0_imag} <<< 9);
  assign _zz_6072 = {{9{_zz_6071[26]}}, _zz_6071};
  assign _zz_6073 = fixTo_579_dout;
  assign _zz_6074 = _zz_6075[35 : 0];
  assign _zz_6075 = _zz_6076;
  assign _zz_6076 = ($signed(_zz_6077) >>> _zz_485);
  assign _zz_6077 = _zz_6078;
  assign _zz_6078 = ($signed(_zz_6080) + $signed(_zz_481));
  assign _zz_6079 = ({9'd0,data_mid_3_0_real} <<< 9);
  assign _zz_6080 = {{9{_zz_6079[26]}}, _zz_6079};
  assign _zz_6081 = fixTo_580_dout;
  assign _zz_6082 = _zz_6083[35 : 0];
  assign _zz_6083 = _zz_6084;
  assign _zz_6084 = ($signed(_zz_6085) >>> _zz_485);
  assign _zz_6085 = _zz_6086;
  assign _zz_6086 = ($signed(_zz_6088) + $signed(_zz_482));
  assign _zz_6087 = ({9'd0,data_mid_3_0_imag} <<< 9);
  assign _zz_6088 = {{9{_zz_6087[26]}}, _zz_6087};
  assign _zz_6089 = fixTo_581_dout;
  assign _zz_6090 = ($signed(twiddle_factor_table_8_real) + $signed(twiddle_factor_table_8_imag));
  assign _zz_6091 = ($signed(_zz_488) - $signed(_zz_6092));
  assign _zz_6092 = ($signed(_zz_6093) * $signed(twiddle_factor_table_8_imag));
  assign _zz_6093 = ($signed(data_mid_3_9_real) + $signed(data_mid_3_9_imag));
  assign _zz_6094 = fixTo_582_dout;
  assign _zz_6095 = ($signed(_zz_488) + $signed(_zz_6096));
  assign _zz_6096 = ($signed(_zz_6097) * $signed(twiddle_factor_table_8_real));
  assign _zz_6097 = ($signed(data_mid_3_9_imag) - $signed(data_mid_3_9_real));
  assign _zz_6098 = fixTo_583_dout;
  assign _zz_6099 = _zz_6100[35 : 0];
  assign _zz_6100 = _zz_6101;
  assign _zz_6101 = ($signed(_zz_6102) >>> _zz_489);
  assign _zz_6102 = _zz_6103;
  assign _zz_6103 = ($signed(_zz_6105) - $signed(_zz_486));
  assign _zz_6104 = ({9'd0,data_mid_3_1_real} <<< 9);
  assign _zz_6105 = {{9{_zz_6104[26]}}, _zz_6104};
  assign _zz_6106 = fixTo_584_dout;
  assign _zz_6107 = _zz_6108[35 : 0];
  assign _zz_6108 = _zz_6109;
  assign _zz_6109 = ($signed(_zz_6110) >>> _zz_489);
  assign _zz_6110 = _zz_6111;
  assign _zz_6111 = ($signed(_zz_6113) - $signed(_zz_487));
  assign _zz_6112 = ({9'd0,data_mid_3_1_imag} <<< 9);
  assign _zz_6113 = {{9{_zz_6112[26]}}, _zz_6112};
  assign _zz_6114 = fixTo_585_dout;
  assign _zz_6115 = _zz_6116[35 : 0];
  assign _zz_6116 = _zz_6117;
  assign _zz_6117 = ($signed(_zz_6118) >>> _zz_490);
  assign _zz_6118 = _zz_6119;
  assign _zz_6119 = ($signed(_zz_6121) + $signed(_zz_486));
  assign _zz_6120 = ({9'd0,data_mid_3_1_real} <<< 9);
  assign _zz_6121 = {{9{_zz_6120[26]}}, _zz_6120};
  assign _zz_6122 = fixTo_586_dout;
  assign _zz_6123 = _zz_6124[35 : 0];
  assign _zz_6124 = _zz_6125;
  assign _zz_6125 = ($signed(_zz_6126) >>> _zz_490);
  assign _zz_6126 = _zz_6127;
  assign _zz_6127 = ($signed(_zz_6129) + $signed(_zz_487));
  assign _zz_6128 = ({9'd0,data_mid_3_1_imag} <<< 9);
  assign _zz_6129 = {{9{_zz_6128[26]}}, _zz_6128};
  assign _zz_6130 = fixTo_587_dout;
  assign _zz_6131 = ($signed(twiddle_factor_table_9_real) + $signed(twiddle_factor_table_9_imag));
  assign _zz_6132 = ($signed(_zz_493) - $signed(_zz_6133));
  assign _zz_6133 = ($signed(_zz_6134) * $signed(twiddle_factor_table_9_imag));
  assign _zz_6134 = ($signed(data_mid_3_10_real) + $signed(data_mid_3_10_imag));
  assign _zz_6135 = fixTo_588_dout;
  assign _zz_6136 = ($signed(_zz_493) + $signed(_zz_6137));
  assign _zz_6137 = ($signed(_zz_6138) * $signed(twiddle_factor_table_9_real));
  assign _zz_6138 = ($signed(data_mid_3_10_imag) - $signed(data_mid_3_10_real));
  assign _zz_6139 = fixTo_589_dout;
  assign _zz_6140 = _zz_6141[35 : 0];
  assign _zz_6141 = _zz_6142;
  assign _zz_6142 = ($signed(_zz_6143) >>> _zz_494);
  assign _zz_6143 = _zz_6144;
  assign _zz_6144 = ($signed(_zz_6146) - $signed(_zz_491));
  assign _zz_6145 = ({9'd0,data_mid_3_2_real} <<< 9);
  assign _zz_6146 = {{9{_zz_6145[26]}}, _zz_6145};
  assign _zz_6147 = fixTo_590_dout;
  assign _zz_6148 = _zz_6149[35 : 0];
  assign _zz_6149 = _zz_6150;
  assign _zz_6150 = ($signed(_zz_6151) >>> _zz_494);
  assign _zz_6151 = _zz_6152;
  assign _zz_6152 = ($signed(_zz_6154) - $signed(_zz_492));
  assign _zz_6153 = ({9'd0,data_mid_3_2_imag} <<< 9);
  assign _zz_6154 = {{9{_zz_6153[26]}}, _zz_6153};
  assign _zz_6155 = fixTo_591_dout;
  assign _zz_6156 = _zz_6157[35 : 0];
  assign _zz_6157 = _zz_6158;
  assign _zz_6158 = ($signed(_zz_6159) >>> _zz_495);
  assign _zz_6159 = _zz_6160;
  assign _zz_6160 = ($signed(_zz_6162) + $signed(_zz_491));
  assign _zz_6161 = ({9'd0,data_mid_3_2_real} <<< 9);
  assign _zz_6162 = {{9{_zz_6161[26]}}, _zz_6161};
  assign _zz_6163 = fixTo_592_dout;
  assign _zz_6164 = _zz_6165[35 : 0];
  assign _zz_6165 = _zz_6166;
  assign _zz_6166 = ($signed(_zz_6167) >>> _zz_495);
  assign _zz_6167 = _zz_6168;
  assign _zz_6168 = ($signed(_zz_6170) + $signed(_zz_492));
  assign _zz_6169 = ({9'd0,data_mid_3_2_imag} <<< 9);
  assign _zz_6170 = {{9{_zz_6169[26]}}, _zz_6169};
  assign _zz_6171 = fixTo_593_dout;
  assign _zz_6172 = ($signed(twiddle_factor_table_10_real) + $signed(twiddle_factor_table_10_imag));
  assign _zz_6173 = ($signed(_zz_498) - $signed(_zz_6174));
  assign _zz_6174 = ($signed(_zz_6175) * $signed(twiddle_factor_table_10_imag));
  assign _zz_6175 = ($signed(data_mid_3_11_real) + $signed(data_mid_3_11_imag));
  assign _zz_6176 = fixTo_594_dout;
  assign _zz_6177 = ($signed(_zz_498) + $signed(_zz_6178));
  assign _zz_6178 = ($signed(_zz_6179) * $signed(twiddle_factor_table_10_real));
  assign _zz_6179 = ($signed(data_mid_3_11_imag) - $signed(data_mid_3_11_real));
  assign _zz_6180 = fixTo_595_dout;
  assign _zz_6181 = _zz_6182[35 : 0];
  assign _zz_6182 = _zz_6183;
  assign _zz_6183 = ($signed(_zz_6184) >>> _zz_499);
  assign _zz_6184 = _zz_6185;
  assign _zz_6185 = ($signed(_zz_6187) - $signed(_zz_496));
  assign _zz_6186 = ({9'd0,data_mid_3_3_real} <<< 9);
  assign _zz_6187 = {{9{_zz_6186[26]}}, _zz_6186};
  assign _zz_6188 = fixTo_596_dout;
  assign _zz_6189 = _zz_6190[35 : 0];
  assign _zz_6190 = _zz_6191;
  assign _zz_6191 = ($signed(_zz_6192) >>> _zz_499);
  assign _zz_6192 = _zz_6193;
  assign _zz_6193 = ($signed(_zz_6195) - $signed(_zz_497));
  assign _zz_6194 = ({9'd0,data_mid_3_3_imag} <<< 9);
  assign _zz_6195 = {{9{_zz_6194[26]}}, _zz_6194};
  assign _zz_6196 = fixTo_597_dout;
  assign _zz_6197 = _zz_6198[35 : 0];
  assign _zz_6198 = _zz_6199;
  assign _zz_6199 = ($signed(_zz_6200) >>> _zz_500);
  assign _zz_6200 = _zz_6201;
  assign _zz_6201 = ($signed(_zz_6203) + $signed(_zz_496));
  assign _zz_6202 = ({9'd0,data_mid_3_3_real} <<< 9);
  assign _zz_6203 = {{9{_zz_6202[26]}}, _zz_6202};
  assign _zz_6204 = fixTo_598_dout;
  assign _zz_6205 = _zz_6206[35 : 0];
  assign _zz_6206 = _zz_6207;
  assign _zz_6207 = ($signed(_zz_6208) >>> _zz_500);
  assign _zz_6208 = _zz_6209;
  assign _zz_6209 = ($signed(_zz_6211) + $signed(_zz_497));
  assign _zz_6210 = ({9'd0,data_mid_3_3_imag} <<< 9);
  assign _zz_6211 = {{9{_zz_6210[26]}}, _zz_6210};
  assign _zz_6212 = fixTo_599_dout;
  assign _zz_6213 = ($signed(twiddle_factor_table_11_real) + $signed(twiddle_factor_table_11_imag));
  assign _zz_6214 = ($signed(_zz_503) - $signed(_zz_6215));
  assign _zz_6215 = ($signed(_zz_6216) * $signed(twiddle_factor_table_11_imag));
  assign _zz_6216 = ($signed(data_mid_3_12_real) + $signed(data_mid_3_12_imag));
  assign _zz_6217 = fixTo_600_dout;
  assign _zz_6218 = ($signed(_zz_503) + $signed(_zz_6219));
  assign _zz_6219 = ($signed(_zz_6220) * $signed(twiddle_factor_table_11_real));
  assign _zz_6220 = ($signed(data_mid_3_12_imag) - $signed(data_mid_3_12_real));
  assign _zz_6221 = fixTo_601_dout;
  assign _zz_6222 = _zz_6223[35 : 0];
  assign _zz_6223 = _zz_6224;
  assign _zz_6224 = ($signed(_zz_6225) >>> _zz_504);
  assign _zz_6225 = _zz_6226;
  assign _zz_6226 = ($signed(_zz_6228) - $signed(_zz_501));
  assign _zz_6227 = ({9'd0,data_mid_3_4_real} <<< 9);
  assign _zz_6228 = {{9{_zz_6227[26]}}, _zz_6227};
  assign _zz_6229 = fixTo_602_dout;
  assign _zz_6230 = _zz_6231[35 : 0];
  assign _zz_6231 = _zz_6232;
  assign _zz_6232 = ($signed(_zz_6233) >>> _zz_504);
  assign _zz_6233 = _zz_6234;
  assign _zz_6234 = ($signed(_zz_6236) - $signed(_zz_502));
  assign _zz_6235 = ({9'd0,data_mid_3_4_imag} <<< 9);
  assign _zz_6236 = {{9{_zz_6235[26]}}, _zz_6235};
  assign _zz_6237 = fixTo_603_dout;
  assign _zz_6238 = _zz_6239[35 : 0];
  assign _zz_6239 = _zz_6240;
  assign _zz_6240 = ($signed(_zz_6241) >>> _zz_505);
  assign _zz_6241 = _zz_6242;
  assign _zz_6242 = ($signed(_zz_6244) + $signed(_zz_501));
  assign _zz_6243 = ({9'd0,data_mid_3_4_real} <<< 9);
  assign _zz_6244 = {{9{_zz_6243[26]}}, _zz_6243};
  assign _zz_6245 = fixTo_604_dout;
  assign _zz_6246 = _zz_6247[35 : 0];
  assign _zz_6247 = _zz_6248;
  assign _zz_6248 = ($signed(_zz_6249) >>> _zz_505);
  assign _zz_6249 = _zz_6250;
  assign _zz_6250 = ($signed(_zz_6252) + $signed(_zz_502));
  assign _zz_6251 = ({9'd0,data_mid_3_4_imag} <<< 9);
  assign _zz_6252 = {{9{_zz_6251[26]}}, _zz_6251};
  assign _zz_6253 = fixTo_605_dout;
  assign _zz_6254 = ($signed(twiddle_factor_table_12_real) + $signed(twiddle_factor_table_12_imag));
  assign _zz_6255 = ($signed(_zz_508) - $signed(_zz_6256));
  assign _zz_6256 = ($signed(_zz_6257) * $signed(twiddle_factor_table_12_imag));
  assign _zz_6257 = ($signed(data_mid_3_13_real) + $signed(data_mid_3_13_imag));
  assign _zz_6258 = fixTo_606_dout;
  assign _zz_6259 = ($signed(_zz_508) + $signed(_zz_6260));
  assign _zz_6260 = ($signed(_zz_6261) * $signed(twiddle_factor_table_12_real));
  assign _zz_6261 = ($signed(data_mid_3_13_imag) - $signed(data_mid_3_13_real));
  assign _zz_6262 = fixTo_607_dout;
  assign _zz_6263 = _zz_6264[35 : 0];
  assign _zz_6264 = _zz_6265;
  assign _zz_6265 = ($signed(_zz_6266) >>> _zz_509);
  assign _zz_6266 = _zz_6267;
  assign _zz_6267 = ($signed(_zz_6269) - $signed(_zz_506));
  assign _zz_6268 = ({9'd0,data_mid_3_5_real} <<< 9);
  assign _zz_6269 = {{9{_zz_6268[26]}}, _zz_6268};
  assign _zz_6270 = fixTo_608_dout;
  assign _zz_6271 = _zz_6272[35 : 0];
  assign _zz_6272 = _zz_6273;
  assign _zz_6273 = ($signed(_zz_6274) >>> _zz_509);
  assign _zz_6274 = _zz_6275;
  assign _zz_6275 = ($signed(_zz_6277) - $signed(_zz_507));
  assign _zz_6276 = ({9'd0,data_mid_3_5_imag} <<< 9);
  assign _zz_6277 = {{9{_zz_6276[26]}}, _zz_6276};
  assign _zz_6278 = fixTo_609_dout;
  assign _zz_6279 = _zz_6280[35 : 0];
  assign _zz_6280 = _zz_6281;
  assign _zz_6281 = ($signed(_zz_6282) >>> _zz_510);
  assign _zz_6282 = _zz_6283;
  assign _zz_6283 = ($signed(_zz_6285) + $signed(_zz_506));
  assign _zz_6284 = ({9'd0,data_mid_3_5_real} <<< 9);
  assign _zz_6285 = {{9{_zz_6284[26]}}, _zz_6284};
  assign _zz_6286 = fixTo_610_dout;
  assign _zz_6287 = _zz_6288[35 : 0];
  assign _zz_6288 = _zz_6289;
  assign _zz_6289 = ($signed(_zz_6290) >>> _zz_510);
  assign _zz_6290 = _zz_6291;
  assign _zz_6291 = ($signed(_zz_6293) + $signed(_zz_507));
  assign _zz_6292 = ({9'd0,data_mid_3_5_imag} <<< 9);
  assign _zz_6293 = {{9{_zz_6292[26]}}, _zz_6292};
  assign _zz_6294 = fixTo_611_dout;
  assign _zz_6295 = ($signed(twiddle_factor_table_13_real) + $signed(twiddle_factor_table_13_imag));
  assign _zz_6296 = ($signed(_zz_513) - $signed(_zz_6297));
  assign _zz_6297 = ($signed(_zz_6298) * $signed(twiddle_factor_table_13_imag));
  assign _zz_6298 = ($signed(data_mid_3_14_real) + $signed(data_mid_3_14_imag));
  assign _zz_6299 = fixTo_612_dout;
  assign _zz_6300 = ($signed(_zz_513) + $signed(_zz_6301));
  assign _zz_6301 = ($signed(_zz_6302) * $signed(twiddle_factor_table_13_real));
  assign _zz_6302 = ($signed(data_mid_3_14_imag) - $signed(data_mid_3_14_real));
  assign _zz_6303 = fixTo_613_dout;
  assign _zz_6304 = _zz_6305[35 : 0];
  assign _zz_6305 = _zz_6306;
  assign _zz_6306 = ($signed(_zz_6307) >>> _zz_514);
  assign _zz_6307 = _zz_6308;
  assign _zz_6308 = ($signed(_zz_6310) - $signed(_zz_511));
  assign _zz_6309 = ({9'd0,data_mid_3_6_real} <<< 9);
  assign _zz_6310 = {{9{_zz_6309[26]}}, _zz_6309};
  assign _zz_6311 = fixTo_614_dout;
  assign _zz_6312 = _zz_6313[35 : 0];
  assign _zz_6313 = _zz_6314;
  assign _zz_6314 = ($signed(_zz_6315) >>> _zz_514);
  assign _zz_6315 = _zz_6316;
  assign _zz_6316 = ($signed(_zz_6318) - $signed(_zz_512));
  assign _zz_6317 = ({9'd0,data_mid_3_6_imag} <<< 9);
  assign _zz_6318 = {{9{_zz_6317[26]}}, _zz_6317};
  assign _zz_6319 = fixTo_615_dout;
  assign _zz_6320 = _zz_6321[35 : 0];
  assign _zz_6321 = _zz_6322;
  assign _zz_6322 = ($signed(_zz_6323) >>> _zz_515);
  assign _zz_6323 = _zz_6324;
  assign _zz_6324 = ($signed(_zz_6326) + $signed(_zz_511));
  assign _zz_6325 = ({9'd0,data_mid_3_6_real} <<< 9);
  assign _zz_6326 = {{9{_zz_6325[26]}}, _zz_6325};
  assign _zz_6327 = fixTo_616_dout;
  assign _zz_6328 = _zz_6329[35 : 0];
  assign _zz_6329 = _zz_6330;
  assign _zz_6330 = ($signed(_zz_6331) >>> _zz_515);
  assign _zz_6331 = _zz_6332;
  assign _zz_6332 = ($signed(_zz_6334) + $signed(_zz_512));
  assign _zz_6333 = ({9'd0,data_mid_3_6_imag} <<< 9);
  assign _zz_6334 = {{9{_zz_6333[26]}}, _zz_6333};
  assign _zz_6335 = fixTo_617_dout;
  assign _zz_6336 = ($signed(twiddle_factor_table_14_real) + $signed(twiddle_factor_table_14_imag));
  assign _zz_6337 = ($signed(_zz_518) - $signed(_zz_6338));
  assign _zz_6338 = ($signed(_zz_6339) * $signed(twiddle_factor_table_14_imag));
  assign _zz_6339 = ($signed(data_mid_3_15_real) + $signed(data_mid_3_15_imag));
  assign _zz_6340 = fixTo_618_dout;
  assign _zz_6341 = ($signed(_zz_518) + $signed(_zz_6342));
  assign _zz_6342 = ($signed(_zz_6343) * $signed(twiddle_factor_table_14_real));
  assign _zz_6343 = ($signed(data_mid_3_15_imag) - $signed(data_mid_3_15_real));
  assign _zz_6344 = fixTo_619_dout;
  assign _zz_6345 = _zz_6346[35 : 0];
  assign _zz_6346 = _zz_6347;
  assign _zz_6347 = ($signed(_zz_6348) >>> _zz_519);
  assign _zz_6348 = _zz_6349;
  assign _zz_6349 = ($signed(_zz_6351) - $signed(_zz_516));
  assign _zz_6350 = ({9'd0,data_mid_3_7_real} <<< 9);
  assign _zz_6351 = {{9{_zz_6350[26]}}, _zz_6350};
  assign _zz_6352 = fixTo_620_dout;
  assign _zz_6353 = _zz_6354[35 : 0];
  assign _zz_6354 = _zz_6355;
  assign _zz_6355 = ($signed(_zz_6356) >>> _zz_519);
  assign _zz_6356 = _zz_6357;
  assign _zz_6357 = ($signed(_zz_6359) - $signed(_zz_517));
  assign _zz_6358 = ({9'd0,data_mid_3_7_imag} <<< 9);
  assign _zz_6359 = {{9{_zz_6358[26]}}, _zz_6358};
  assign _zz_6360 = fixTo_621_dout;
  assign _zz_6361 = _zz_6362[35 : 0];
  assign _zz_6362 = _zz_6363;
  assign _zz_6363 = ($signed(_zz_6364) >>> _zz_520);
  assign _zz_6364 = _zz_6365;
  assign _zz_6365 = ($signed(_zz_6367) + $signed(_zz_516));
  assign _zz_6366 = ({9'd0,data_mid_3_7_real} <<< 9);
  assign _zz_6367 = {{9{_zz_6366[26]}}, _zz_6366};
  assign _zz_6368 = fixTo_622_dout;
  assign _zz_6369 = _zz_6370[35 : 0];
  assign _zz_6370 = _zz_6371;
  assign _zz_6371 = ($signed(_zz_6372) >>> _zz_520);
  assign _zz_6372 = _zz_6373;
  assign _zz_6373 = ($signed(_zz_6375) + $signed(_zz_517));
  assign _zz_6374 = ({9'd0,data_mid_3_7_imag} <<< 9);
  assign _zz_6375 = {{9{_zz_6374[26]}}, _zz_6374};
  assign _zz_6376 = fixTo_623_dout;
  assign _zz_6377 = ($signed(twiddle_factor_table_7_real) + $signed(twiddle_factor_table_7_imag));
  assign _zz_6378 = ($signed(_zz_523) - $signed(_zz_6379));
  assign _zz_6379 = ($signed(_zz_6380) * $signed(twiddle_factor_table_7_imag));
  assign _zz_6380 = ($signed(data_mid_3_24_real) + $signed(data_mid_3_24_imag));
  assign _zz_6381 = fixTo_624_dout;
  assign _zz_6382 = ($signed(_zz_523) + $signed(_zz_6383));
  assign _zz_6383 = ($signed(_zz_6384) * $signed(twiddle_factor_table_7_real));
  assign _zz_6384 = ($signed(data_mid_3_24_imag) - $signed(data_mid_3_24_real));
  assign _zz_6385 = fixTo_625_dout;
  assign _zz_6386 = _zz_6387[35 : 0];
  assign _zz_6387 = _zz_6388;
  assign _zz_6388 = ($signed(_zz_6389) >>> _zz_524);
  assign _zz_6389 = _zz_6390;
  assign _zz_6390 = ($signed(_zz_6392) - $signed(_zz_521));
  assign _zz_6391 = ({9'd0,data_mid_3_16_real} <<< 9);
  assign _zz_6392 = {{9{_zz_6391[26]}}, _zz_6391};
  assign _zz_6393 = fixTo_626_dout;
  assign _zz_6394 = _zz_6395[35 : 0];
  assign _zz_6395 = _zz_6396;
  assign _zz_6396 = ($signed(_zz_6397) >>> _zz_524);
  assign _zz_6397 = _zz_6398;
  assign _zz_6398 = ($signed(_zz_6400) - $signed(_zz_522));
  assign _zz_6399 = ({9'd0,data_mid_3_16_imag} <<< 9);
  assign _zz_6400 = {{9{_zz_6399[26]}}, _zz_6399};
  assign _zz_6401 = fixTo_627_dout;
  assign _zz_6402 = _zz_6403[35 : 0];
  assign _zz_6403 = _zz_6404;
  assign _zz_6404 = ($signed(_zz_6405) >>> _zz_525);
  assign _zz_6405 = _zz_6406;
  assign _zz_6406 = ($signed(_zz_6408) + $signed(_zz_521));
  assign _zz_6407 = ({9'd0,data_mid_3_16_real} <<< 9);
  assign _zz_6408 = {{9{_zz_6407[26]}}, _zz_6407};
  assign _zz_6409 = fixTo_628_dout;
  assign _zz_6410 = _zz_6411[35 : 0];
  assign _zz_6411 = _zz_6412;
  assign _zz_6412 = ($signed(_zz_6413) >>> _zz_525);
  assign _zz_6413 = _zz_6414;
  assign _zz_6414 = ($signed(_zz_6416) + $signed(_zz_522));
  assign _zz_6415 = ({9'd0,data_mid_3_16_imag} <<< 9);
  assign _zz_6416 = {{9{_zz_6415[26]}}, _zz_6415};
  assign _zz_6417 = fixTo_629_dout;
  assign _zz_6418 = ($signed(twiddle_factor_table_8_real) + $signed(twiddle_factor_table_8_imag));
  assign _zz_6419 = ($signed(_zz_528) - $signed(_zz_6420));
  assign _zz_6420 = ($signed(_zz_6421) * $signed(twiddle_factor_table_8_imag));
  assign _zz_6421 = ($signed(data_mid_3_25_real) + $signed(data_mid_3_25_imag));
  assign _zz_6422 = fixTo_630_dout;
  assign _zz_6423 = ($signed(_zz_528) + $signed(_zz_6424));
  assign _zz_6424 = ($signed(_zz_6425) * $signed(twiddle_factor_table_8_real));
  assign _zz_6425 = ($signed(data_mid_3_25_imag) - $signed(data_mid_3_25_real));
  assign _zz_6426 = fixTo_631_dout;
  assign _zz_6427 = _zz_6428[35 : 0];
  assign _zz_6428 = _zz_6429;
  assign _zz_6429 = ($signed(_zz_6430) >>> _zz_529);
  assign _zz_6430 = _zz_6431;
  assign _zz_6431 = ($signed(_zz_6433) - $signed(_zz_526));
  assign _zz_6432 = ({9'd0,data_mid_3_17_real} <<< 9);
  assign _zz_6433 = {{9{_zz_6432[26]}}, _zz_6432};
  assign _zz_6434 = fixTo_632_dout;
  assign _zz_6435 = _zz_6436[35 : 0];
  assign _zz_6436 = _zz_6437;
  assign _zz_6437 = ($signed(_zz_6438) >>> _zz_529);
  assign _zz_6438 = _zz_6439;
  assign _zz_6439 = ($signed(_zz_6441) - $signed(_zz_527));
  assign _zz_6440 = ({9'd0,data_mid_3_17_imag} <<< 9);
  assign _zz_6441 = {{9{_zz_6440[26]}}, _zz_6440};
  assign _zz_6442 = fixTo_633_dout;
  assign _zz_6443 = _zz_6444[35 : 0];
  assign _zz_6444 = _zz_6445;
  assign _zz_6445 = ($signed(_zz_6446) >>> _zz_530);
  assign _zz_6446 = _zz_6447;
  assign _zz_6447 = ($signed(_zz_6449) + $signed(_zz_526));
  assign _zz_6448 = ({9'd0,data_mid_3_17_real} <<< 9);
  assign _zz_6449 = {{9{_zz_6448[26]}}, _zz_6448};
  assign _zz_6450 = fixTo_634_dout;
  assign _zz_6451 = _zz_6452[35 : 0];
  assign _zz_6452 = _zz_6453;
  assign _zz_6453 = ($signed(_zz_6454) >>> _zz_530);
  assign _zz_6454 = _zz_6455;
  assign _zz_6455 = ($signed(_zz_6457) + $signed(_zz_527));
  assign _zz_6456 = ({9'd0,data_mid_3_17_imag} <<< 9);
  assign _zz_6457 = {{9{_zz_6456[26]}}, _zz_6456};
  assign _zz_6458 = fixTo_635_dout;
  assign _zz_6459 = ($signed(twiddle_factor_table_9_real) + $signed(twiddle_factor_table_9_imag));
  assign _zz_6460 = ($signed(_zz_533) - $signed(_zz_6461));
  assign _zz_6461 = ($signed(_zz_6462) * $signed(twiddle_factor_table_9_imag));
  assign _zz_6462 = ($signed(data_mid_3_26_real) + $signed(data_mid_3_26_imag));
  assign _zz_6463 = fixTo_636_dout;
  assign _zz_6464 = ($signed(_zz_533) + $signed(_zz_6465));
  assign _zz_6465 = ($signed(_zz_6466) * $signed(twiddle_factor_table_9_real));
  assign _zz_6466 = ($signed(data_mid_3_26_imag) - $signed(data_mid_3_26_real));
  assign _zz_6467 = fixTo_637_dout;
  assign _zz_6468 = _zz_6469[35 : 0];
  assign _zz_6469 = _zz_6470;
  assign _zz_6470 = ($signed(_zz_6471) >>> _zz_534);
  assign _zz_6471 = _zz_6472;
  assign _zz_6472 = ($signed(_zz_6474) - $signed(_zz_531));
  assign _zz_6473 = ({9'd0,data_mid_3_18_real} <<< 9);
  assign _zz_6474 = {{9{_zz_6473[26]}}, _zz_6473};
  assign _zz_6475 = fixTo_638_dout;
  assign _zz_6476 = _zz_6477[35 : 0];
  assign _zz_6477 = _zz_6478;
  assign _zz_6478 = ($signed(_zz_6479) >>> _zz_534);
  assign _zz_6479 = _zz_6480;
  assign _zz_6480 = ($signed(_zz_6482) - $signed(_zz_532));
  assign _zz_6481 = ({9'd0,data_mid_3_18_imag} <<< 9);
  assign _zz_6482 = {{9{_zz_6481[26]}}, _zz_6481};
  assign _zz_6483 = fixTo_639_dout;
  assign _zz_6484 = _zz_6485[35 : 0];
  assign _zz_6485 = _zz_6486;
  assign _zz_6486 = ($signed(_zz_6487) >>> _zz_535);
  assign _zz_6487 = _zz_6488;
  assign _zz_6488 = ($signed(_zz_6490) + $signed(_zz_531));
  assign _zz_6489 = ({9'd0,data_mid_3_18_real} <<< 9);
  assign _zz_6490 = {{9{_zz_6489[26]}}, _zz_6489};
  assign _zz_6491 = fixTo_640_dout;
  assign _zz_6492 = _zz_6493[35 : 0];
  assign _zz_6493 = _zz_6494;
  assign _zz_6494 = ($signed(_zz_6495) >>> _zz_535);
  assign _zz_6495 = _zz_6496;
  assign _zz_6496 = ($signed(_zz_6498) + $signed(_zz_532));
  assign _zz_6497 = ({9'd0,data_mid_3_18_imag} <<< 9);
  assign _zz_6498 = {{9{_zz_6497[26]}}, _zz_6497};
  assign _zz_6499 = fixTo_641_dout;
  assign _zz_6500 = ($signed(twiddle_factor_table_10_real) + $signed(twiddle_factor_table_10_imag));
  assign _zz_6501 = ($signed(_zz_538) - $signed(_zz_6502));
  assign _zz_6502 = ($signed(_zz_6503) * $signed(twiddle_factor_table_10_imag));
  assign _zz_6503 = ($signed(data_mid_3_27_real) + $signed(data_mid_3_27_imag));
  assign _zz_6504 = fixTo_642_dout;
  assign _zz_6505 = ($signed(_zz_538) + $signed(_zz_6506));
  assign _zz_6506 = ($signed(_zz_6507) * $signed(twiddle_factor_table_10_real));
  assign _zz_6507 = ($signed(data_mid_3_27_imag) - $signed(data_mid_3_27_real));
  assign _zz_6508 = fixTo_643_dout;
  assign _zz_6509 = _zz_6510[35 : 0];
  assign _zz_6510 = _zz_6511;
  assign _zz_6511 = ($signed(_zz_6512) >>> _zz_539);
  assign _zz_6512 = _zz_6513;
  assign _zz_6513 = ($signed(_zz_6515) - $signed(_zz_536));
  assign _zz_6514 = ({9'd0,data_mid_3_19_real} <<< 9);
  assign _zz_6515 = {{9{_zz_6514[26]}}, _zz_6514};
  assign _zz_6516 = fixTo_644_dout;
  assign _zz_6517 = _zz_6518[35 : 0];
  assign _zz_6518 = _zz_6519;
  assign _zz_6519 = ($signed(_zz_6520) >>> _zz_539);
  assign _zz_6520 = _zz_6521;
  assign _zz_6521 = ($signed(_zz_6523) - $signed(_zz_537));
  assign _zz_6522 = ({9'd0,data_mid_3_19_imag} <<< 9);
  assign _zz_6523 = {{9{_zz_6522[26]}}, _zz_6522};
  assign _zz_6524 = fixTo_645_dout;
  assign _zz_6525 = _zz_6526[35 : 0];
  assign _zz_6526 = _zz_6527;
  assign _zz_6527 = ($signed(_zz_6528) >>> _zz_540);
  assign _zz_6528 = _zz_6529;
  assign _zz_6529 = ($signed(_zz_6531) + $signed(_zz_536));
  assign _zz_6530 = ({9'd0,data_mid_3_19_real} <<< 9);
  assign _zz_6531 = {{9{_zz_6530[26]}}, _zz_6530};
  assign _zz_6532 = fixTo_646_dout;
  assign _zz_6533 = _zz_6534[35 : 0];
  assign _zz_6534 = _zz_6535;
  assign _zz_6535 = ($signed(_zz_6536) >>> _zz_540);
  assign _zz_6536 = _zz_6537;
  assign _zz_6537 = ($signed(_zz_6539) + $signed(_zz_537));
  assign _zz_6538 = ({9'd0,data_mid_3_19_imag} <<< 9);
  assign _zz_6539 = {{9{_zz_6538[26]}}, _zz_6538};
  assign _zz_6540 = fixTo_647_dout;
  assign _zz_6541 = ($signed(twiddle_factor_table_11_real) + $signed(twiddle_factor_table_11_imag));
  assign _zz_6542 = ($signed(_zz_543) - $signed(_zz_6543));
  assign _zz_6543 = ($signed(_zz_6544) * $signed(twiddle_factor_table_11_imag));
  assign _zz_6544 = ($signed(data_mid_3_28_real) + $signed(data_mid_3_28_imag));
  assign _zz_6545 = fixTo_648_dout;
  assign _zz_6546 = ($signed(_zz_543) + $signed(_zz_6547));
  assign _zz_6547 = ($signed(_zz_6548) * $signed(twiddle_factor_table_11_real));
  assign _zz_6548 = ($signed(data_mid_3_28_imag) - $signed(data_mid_3_28_real));
  assign _zz_6549 = fixTo_649_dout;
  assign _zz_6550 = _zz_6551[35 : 0];
  assign _zz_6551 = _zz_6552;
  assign _zz_6552 = ($signed(_zz_6553) >>> _zz_544);
  assign _zz_6553 = _zz_6554;
  assign _zz_6554 = ($signed(_zz_6556) - $signed(_zz_541));
  assign _zz_6555 = ({9'd0,data_mid_3_20_real} <<< 9);
  assign _zz_6556 = {{9{_zz_6555[26]}}, _zz_6555};
  assign _zz_6557 = fixTo_650_dout;
  assign _zz_6558 = _zz_6559[35 : 0];
  assign _zz_6559 = _zz_6560;
  assign _zz_6560 = ($signed(_zz_6561) >>> _zz_544);
  assign _zz_6561 = _zz_6562;
  assign _zz_6562 = ($signed(_zz_6564) - $signed(_zz_542));
  assign _zz_6563 = ({9'd0,data_mid_3_20_imag} <<< 9);
  assign _zz_6564 = {{9{_zz_6563[26]}}, _zz_6563};
  assign _zz_6565 = fixTo_651_dout;
  assign _zz_6566 = _zz_6567[35 : 0];
  assign _zz_6567 = _zz_6568;
  assign _zz_6568 = ($signed(_zz_6569) >>> _zz_545);
  assign _zz_6569 = _zz_6570;
  assign _zz_6570 = ($signed(_zz_6572) + $signed(_zz_541));
  assign _zz_6571 = ({9'd0,data_mid_3_20_real} <<< 9);
  assign _zz_6572 = {{9{_zz_6571[26]}}, _zz_6571};
  assign _zz_6573 = fixTo_652_dout;
  assign _zz_6574 = _zz_6575[35 : 0];
  assign _zz_6575 = _zz_6576;
  assign _zz_6576 = ($signed(_zz_6577) >>> _zz_545);
  assign _zz_6577 = _zz_6578;
  assign _zz_6578 = ($signed(_zz_6580) + $signed(_zz_542));
  assign _zz_6579 = ({9'd0,data_mid_3_20_imag} <<< 9);
  assign _zz_6580 = {{9{_zz_6579[26]}}, _zz_6579};
  assign _zz_6581 = fixTo_653_dout;
  assign _zz_6582 = ($signed(twiddle_factor_table_12_real) + $signed(twiddle_factor_table_12_imag));
  assign _zz_6583 = ($signed(_zz_548) - $signed(_zz_6584));
  assign _zz_6584 = ($signed(_zz_6585) * $signed(twiddle_factor_table_12_imag));
  assign _zz_6585 = ($signed(data_mid_3_29_real) + $signed(data_mid_3_29_imag));
  assign _zz_6586 = fixTo_654_dout;
  assign _zz_6587 = ($signed(_zz_548) + $signed(_zz_6588));
  assign _zz_6588 = ($signed(_zz_6589) * $signed(twiddle_factor_table_12_real));
  assign _zz_6589 = ($signed(data_mid_3_29_imag) - $signed(data_mid_3_29_real));
  assign _zz_6590 = fixTo_655_dout;
  assign _zz_6591 = _zz_6592[35 : 0];
  assign _zz_6592 = _zz_6593;
  assign _zz_6593 = ($signed(_zz_6594) >>> _zz_549);
  assign _zz_6594 = _zz_6595;
  assign _zz_6595 = ($signed(_zz_6597) - $signed(_zz_546));
  assign _zz_6596 = ({9'd0,data_mid_3_21_real} <<< 9);
  assign _zz_6597 = {{9{_zz_6596[26]}}, _zz_6596};
  assign _zz_6598 = fixTo_656_dout;
  assign _zz_6599 = _zz_6600[35 : 0];
  assign _zz_6600 = _zz_6601;
  assign _zz_6601 = ($signed(_zz_6602) >>> _zz_549);
  assign _zz_6602 = _zz_6603;
  assign _zz_6603 = ($signed(_zz_6605) - $signed(_zz_547));
  assign _zz_6604 = ({9'd0,data_mid_3_21_imag} <<< 9);
  assign _zz_6605 = {{9{_zz_6604[26]}}, _zz_6604};
  assign _zz_6606 = fixTo_657_dout;
  assign _zz_6607 = _zz_6608[35 : 0];
  assign _zz_6608 = _zz_6609;
  assign _zz_6609 = ($signed(_zz_6610) >>> _zz_550);
  assign _zz_6610 = _zz_6611;
  assign _zz_6611 = ($signed(_zz_6613) + $signed(_zz_546));
  assign _zz_6612 = ({9'd0,data_mid_3_21_real} <<< 9);
  assign _zz_6613 = {{9{_zz_6612[26]}}, _zz_6612};
  assign _zz_6614 = fixTo_658_dout;
  assign _zz_6615 = _zz_6616[35 : 0];
  assign _zz_6616 = _zz_6617;
  assign _zz_6617 = ($signed(_zz_6618) >>> _zz_550);
  assign _zz_6618 = _zz_6619;
  assign _zz_6619 = ($signed(_zz_6621) + $signed(_zz_547));
  assign _zz_6620 = ({9'd0,data_mid_3_21_imag} <<< 9);
  assign _zz_6621 = {{9{_zz_6620[26]}}, _zz_6620};
  assign _zz_6622 = fixTo_659_dout;
  assign _zz_6623 = ($signed(twiddle_factor_table_13_real) + $signed(twiddle_factor_table_13_imag));
  assign _zz_6624 = ($signed(_zz_553) - $signed(_zz_6625));
  assign _zz_6625 = ($signed(_zz_6626) * $signed(twiddle_factor_table_13_imag));
  assign _zz_6626 = ($signed(data_mid_3_30_real) + $signed(data_mid_3_30_imag));
  assign _zz_6627 = fixTo_660_dout;
  assign _zz_6628 = ($signed(_zz_553) + $signed(_zz_6629));
  assign _zz_6629 = ($signed(_zz_6630) * $signed(twiddle_factor_table_13_real));
  assign _zz_6630 = ($signed(data_mid_3_30_imag) - $signed(data_mid_3_30_real));
  assign _zz_6631 = fixTo_661_dout;
  assign _zz_6632 = _zz_6633[35 : 0];
  assign _zz_6633 = _zz_6634;
  assign _zz_6634 = ($signed(_zz_6635) >>> _zz_554);
  assign _zz_6635 = _zz_6636;
  assign _zz_6636 = ($signed(_zz_6638) - $signed(_zz_551));
  assign _zz_6637 = ({9'd0,data_mid_3_22_real} <<< 9);
  assign _zz_6638 = {{9{_zz_6637[26]}}, _zz_6637};
  assign _zz_6639 = fixTo_662_dout;
  assign _zz_6640 = _zz_6641[35 : 0];
  assign _zz_6641 = _zz_6642;
  assign _zz_6642 = ($signed(_zz_6643) >>> _zz_554);
  assign _zz_6643 = _zz_6644;
  assign _zz_6644 = ($signed(_zz_6646) - $signed(_zz_552));
  assign _zz_6645 = ({9'd0,data_mid_3_22_imag} <<< 9);
  assign _zz_6646 = {{9{_zz_6645[26]}}, _zz_6645};
  assign _zz_6647 = fixTo_663_dout;
  assign _zz_6648 = _zz_6649[35 : 0];
  assign _zz_6649 = _zz_6650;
  assign _zz_6650 = ($signed(_zz_6651) >>> _zz_555);
  assign _zz_6651 = _zz_6652;
  assign _zz_6652 = ($signed(_zz_6654) + $signed(_zz_551));
  assign _zz_6653 = ({9'd0,data_mid_3_22_real} <<< 9);
  assign _zz_6654 = {{9{_zz_6653[26]}}, _zz_6653};
  assign _zz_6655 = fixTo_664_dout;
  assign _zz_6656 = _zz_6657[35 : 0];
  assign _zz_6657 = _zz_6658;
  assign _zz_6658 = ($signed(_zz_6659) >>> _zz_555);
  assign _zz_6659 = _zz_6660;
  assign _zz_6660 = ($signed(_zz_6662) + $signed(_zz_552));
  assign _zz_6661 = ({9'd0,data_mid_3_22_imag} <<< 9);
  assign _zz_6662 = {{9{_zz_6661[26]}}, _zz_6661};
  assign _zz_6663 = fixTo_665_dout;
  assign _zz_6664 = ($signed(twiddle_factor_table_14_real) + $signed(twiddle_factor_table_14_imag));
  assign _zz_6665 = ($signed(_zz_558) - $signed(_zz_6666));
  assign _zz_6666 = ($signed(_zz_6667) * $signed(twiddle_factor_table_14_imag));
  assign _zz_6667 = ($signed(data_mid_3_31_real) + $signed(data_mid_3_31_imag));
  assign _zz_6668 = fixTo_666_dout;
  assign _zz_6669 = ($signed(_zz_558) + $signed(_zz_6670));
  assign _zz_6670 = ($signed(_zz_6671) * $signed(twiddle_factor_table_14_real));
  assign _zz_6671 = ($signed(data_mid_3_31_imag) - $signed(data_mid_3_31_real));
  assign _zz_6672 = fixTo_667_dout;
  assign _zz_6673 = _zz_6674[35 : 0];
  assign _zz_6674 = _zz_6675;
  assign _zz_6675 = ($signed(_zz_6676) >>> _zz_559);
  assign _zz_6676 = _zz_6677;
  assign _zz_6677 = ($signed(_zz_6679) - $signed(_zz_556));
  assign _zz_6678 = ({9'd0,data_mid_3_23_real} <<< 9);
  assign _zz_6679 = {{9{_zz_6678[26]}}, _zz_6678};
  assign _zz_6680 = fixTo_668_dout;
  assign _zz_6681 = _zz_6682[35 : 0];
  assign _zz_6682 = _zz_6683;
  assign _zz_6683 = ($signed(_zz_6684) >>> _zz_559);
  assign _zz_6684 = _zz_6685;
  assign _zz_6685 = ($signed(_zz_6687) - $signed(_zz_557));
  assign _zz_6686 = ({9'd0,data_mid_3_23_imag} <<< 9);
  assign _zz_6687 = {{9{_zz_6686[26]}}, _zz_6686};
  assign _zz_6688 = fixTo_669_dout;
  assign _zz_6689 = _zz_6690[35 : 0];
  assign _zz_6690 = _zz_6691;
  assign _zz_6691 = ($signed(_zz_6692) >>> _zz_560);
  assign _zz_6692 = _zz_6693;
  assign _zz_6693 = ($signed(_zz_6695) + $signed(_zz_556));
  assign _zz_6694 = ({9'd0,data_mid_3_23_real} <<< 9);
  assign _zz_6695 = {{9{_zz_6694[26]}}, _zz_6694};
  assign _zz_6696 = fixTo_670_dout;
  assign _zz_6697 = _zz_6698[35 : 0];
  assign _zz_6698 = _zz_6699;
  assign _zz_6699 = ($signed(_zz_6700) >>> _zz_560);
  assign _zz_6700 = _zz_6701;
  assign _zz_6701 = ($signed(_zz_6703) + $signed(_zz_557));
  assign _zz_6702 = ({9'd0,data_mid_3_23_imag} <<< 9);
  assign _zz_6703 = {{9{_zz_6702[26]}}, _zz_6702};
  assign _zz_6704 = fixTo_671_dout;
  assign _zz_6705 = ($signed(twiddle_factor_table_7_real) + $signed(twiddle_factor_table_7_imag));
  assign _zz_6706 = ($signed(_zz_563) - $signed(_zz_6707));
  assign _zz_6707 = ($signed(_zz_6708) * $signed(twiddle_factor_table_7_imag));
  assign _zz_6708 = ($signed(data_mid_3_40_real) + $signed(data_mid_3_40_imag));
  assign _zz_6709 = fixTo_672_dout;
  assign _zz_6710 = ($signed(_zz_563) + $signed(_zz_6711));
  assign _zz_6711 = ($signed(_zz_6712) * $signed(twiddle_factor_table_7_real));
  assign _zz_6712 = ($signed(data_mid_3_40_imag) - $signed(data_mid_3_40_real));
  assign _zz_6713 = fixTo_673_dout;
  assign _zz_6714 = _zz_6715[35 : 0];
  assign _zz_6715 = _zz_6716;
  assign _zz_6716 = ($signed(_zz_6717) >>> _zz_564);
  assign _zz_6717 = _zz_6718;
  assign _zz_6718 = ($signed(_zz_6720) - $signed(_zz_561));
  assign _zz_6719 = ({9'd0,data_mid_3_32_real} <<< 9);
  assign _zz_6720 = {{9{_zz_6719[26]}}, _zz_6719};
  assign _zz_6721 = fixTo_674_dout;
  assign _zz_6722 = _zz_6723[35 : 0];
  assign _zz_6723 = _zz_6724;
  assign _zz_6724 = ($signed(_zz_6725) >>> _zz_564);
  assign _zz_6725 = _zz_6726;
  assign _zz_6726 = ($signed(_zz_6728) - $signed(_zz_562));
  assign _zz_6727 = ({9'd0,data_mid_3_32_imag} <<< 9);
  assign _zz_6728 = {{9{_zz_6727[26]}}, _zz_6727};
  assign _zz_6729 = fixTo_675_dout;
  assign _zz_6730 = _zz_6731[35 : 0];
  assign _zz_6731 = _zz_6732;
  assign _zz_6732 = ($signed(_zz_6733) >>> _zz_565);
  assign _zz_6733 = _zz_6734;
  assign _zz_6734 = ($signed(_zz_6736) + $signed(_zz_561));
  assign _zz_6735 = ({9'd0,data_mid_3_32_real} <<< 9);
  assign _zz_6736 = {{9{_zz_6735[26]}}, _zz_6735};
  assign _zz_6737 = fixTo_676_dout;
  assign _zz_6738 = _zz_6739[35 : 0];
  assign _zz_6739 = _zz_6740;
  assign _zz_6740 = ($signed(_zz_6741) >>> _zz_565);
  assign _zz_6741 = _zz_6742;
  assign _zz_6742 = ($signed(_zz_6744) + $signed(_zz_562));
  assign _zz_6743 = ({9'd0,data_mid_3_32_imag} <<< 9);
  assign _zz_6744 = {{9{_zz_6743[26]}}, _zz_6743};
  assign _zz_6745 = fixTo_677_dout;
  assign _zz_6746 = ($signed(twiddle_factor_table_8_real) + $signed(twiddle_factor_table_8_imag));
  assign _zz_6747 = ($signed(_zz_568) - $signed(_zz_6748));
  assign _zz_6748 = ($signed(_zz_6749) * $signed(twiddle_factor_table_8_imag));
  assign _zz_6749 = ($signed(data_mid_3_41_real) + $signed(data_mid_3_41_imag));
  assign _zz_6750 = fixTo_678_dout;
  assign _zz_6751 = ($signed(_zz_568) + $signed(_zz_6752));
  assign _zz_6752 = ($signed(_zz_6753) * $signed(twiddle_factor_table_8_real));
  assign _zz_6753 = ($signed(data_mid_3_41_imag) - $signed(data_mid_3_41_real));
  assign _zz_6754 = fixTo_679_dout;
  assign _zz_6755 = _zz_6756[35 : 0];
  assign _zz_6756 = _zz_6757;
  assign _zz_6757 = ($signed(_zz_6758) >>> _zz_569);
  assign _zz_6758 = _zz_6759;
  assign _zz_6759 = ($signed(_zz_6761) - $signed(_zz_566));
  assign _zz_6760 = ({9'd0,data_mid_3_33_real} <<< 9);
  assign _zz_6761 = {{9{_zz_6760[26]}}, _zz_6760};
  assign _zz_6762 = fixTo_680_dout;
  assign _zz_6763 = _zz_6764[35 : 0];
  assign _zz_6764 = _zz_6765;
  assign _zz_6765 = ($signed(_zz_6766) >>> _zz_569);
  assign _zz_6766 = _zz_6767;
  assign _zz_6767 = ($signed(_zz_6769) - $signed(_zz_567));
  assign _zz_6768 = ({9'd0,data_mid_3_33_imag} <<< 9);
  assign _zz_6769 = {{9{_zz_6768[26]}}, _zz_6768};
  assign _zz_6770 = fixTo_681_dout;
  assign _zz_6771 = _zz_6772[35 : 0];
  assign _zz_6772 = _zz_6773;
  assign _zz_6773 = ($signed(_zz_6774) >>> _zz_570);
  assign _zz_6774 = _zz_6775;
  assign _zz_6775 = ($signed(_zz_6777) + $signed(_zz_566));
  assign _zz_6776 = ({9'd0,data_mid_3_33_real} <<< 9);
  assign _zz_6777 = {{9{_zz_6776[26]}}, _zz_6776};
  assign _zz_6778 = fixTo_682_dout;
  assign _zz_6779 = _zz_6780[35 : 0];
  assign _zz_6780 = _zz_6781;
  assign _zz_6781 = ($signed(_zz_6782) >>> _zz_570);
  assign _zz_6782 = _zz_6783;
  assign _zz_6783 = ($signed(_zz_6785) + $signed(_zz_567));
  assign _zz_6784 = ({9'd0,data_mid_3_33_imag} <<< 9);
  assign _zz_6785 = {{9{_zz_6784[26]}}, _zz_6784};
  assign _zz_6786 = fixTo_683_dout;
  assign _zz_6787 = ($signed(twiddle_factor_table_9_real) + $signed(twiddle_factor_table_9_imag));
  assign _zz_6788 = ($signed(_zz_573) - $signed(_zz_6789));
  assign _zz_6789 = ($signed(_zz_6790) * $signed(twiddle_factor_table_9_imag));
  assign _zz_6790 = ($signed(data_mid_3_42_real) + $signed(data_mid_3_42_imag));
  assign _zz_6791 = fixTo_684_dout;
  assign _zz_6792 = ($signed(_zz_573) + $signed(_zz_6793));
  assign _zz_6793 = ($signed(_zz_6794) * $signed(twiddle_factor_table_9_real));
  assign _zz_6794 = ($signed(data_mid_3_42_imag) - $signed(data_mid_3_42_real));
  assign _zz_6795 = fixTo_685_dout;
  assign _zz_6796 = _zz_6797[35 : 0];
  assign _zz_6797 = _zz_6798;
  assign _zz_6798 = ($signed(_zz_6799) >>> _zz_574);
  assign _zz_6799 = _zz_6800;
  assign _zz_6800 = ($signed(_zz_6802) - $signed(_zz_571));
  assign _zz_6801 = ({9'd0,data_mid_3_34_real} <<< 9);
  assign _zz_6802 = {{9{_zz_6801[26]}}, _zz_6801};
  assign _zz_6803 = fixTo_686_dout;
  assign _zz_6804 = _zz_6805[35 : 0];
  assign _zz_6805 = _zz_6806;
  assign _zz_6806 = ($signed(_zz_6807) >>> _zz_574);
  assign _zz_6807 = _zz_6808;
  assign _zz_6808 = ($signed(_zz_6810) - $signed(_zz_572));
  assign _zz_6809 = ({9'd0,data_mid_3_34_imag} <<< 9);
  assign _zz_6810 = {{9{_zz_6809[26]}}, _zz_6809};
  assign _zz_6811 = fixTo_687_dout;
  assign _zz_6812 = _zz_6813[35 : 0];
  assign _zz_6813 = _zz_6814;
  assign _zz_6814 = ($signed(_zz_6815) >>> _zz_575);
  assign _zz_6815 = _zz_6816;
  assign _zz_6816 = ($signed(_zz_6818) + $signed(_zz_571));
  assign _zz_6817 = ({9'd0,data_mid_3_34_real} <<< 9);
  assign _zz_6818 = {{9{_zz_6817[26]}}, _zz_6817};
  assign _zz_6819 = fixTo_688_dout;
  assign _zz_6820 = _zz_6821[35 : 0];
  assign _zz_6821 = _zz_6822;
  assign _zz_6822 = ($signed(_zz_6823) >>> _zz_575);
  assign _zz_6823 = _zz_6824;
  assign _zz_6824 = ($signed(_zz_6826) + $signed(_zz_572));
  assign _zz_6825 = ({9'd0,data_mid_3_34_imag} <<< 9);
  assign _zz_6826 = {{9{_zz_6825[26]}}, _zz_6825};
  assign _zz_6827 = fixTo_689_dout;
  assign _zz_6828 = ($signed(twiddle_factor_table_10_real) + $signed(twiddle_factor_table_10_imag));
  assign _zz_6829 = ($signed(_zz_578) - $signed(_zz_6830));
  assign _zz_6830 = ($signed(_zz_6831) * $signed(twiddle_factor_table_10_imag));
  assign _zz_6831 = ($signed(data_mid_3_43_real) + $signed(data_mid_3_43_imag));
  assign _zz_6832 = fixTo_690_dout;
  assign _zz_6833 = ($signed(_zz_578) + $signed(_zz_6834));
  assign _zz_6834 = ($signed(_zz_6835) * $signed(twiddle_factor_table_10_real));
  assign _zz_6835 = ($signed(data_mid_3_43_imag) - $signed(data_mid_3_43_real));
  assign _zz_6836 = fixTo_691_dout;
  assign _zz_6837 = _zz_6838[35 : 0];
  assign _zz_6838 = _zz_6839;
  assign _zz_6839 = ($signed(_zz_6840) >>> _zz_579);
  assign _zz_6840 = _zz_6841;
  assign _zz_6841 = ($signed(_zz_6843) - $signed(_zz_576));
  assign _zz_6842 = ({9'd0,data_mid_3_35_real} <<< 9);
  assign _zz_6843 = {{9{_zz_6842[26]}}, _zz_6842};
  assign _zz_6844 = fixTo_692_dout;
  assign _zz_6845 = _zz_6846[35 : 0];
  assign _zz_6846 = _zz_6847;
  assign _zz_6847 = ($signed(_zz_6848) >>> _zz_579);
  assign _zz_6848 = _zz_6849;
  assign _zz_6849 = ($signed(_zz_6851) - $signed(_zz_577));
  assign _zz_6850 = ({9'd0,data_mid_3_35_imag} <<< 9);
  assign _zz_6851 = {{9{_zz_6850[26]}}, _zz_6850};
  assign _zz_6852 = fixTo_693_dout;
  assign _zz_6853 = _zz_6854[35 : 0];
  assign _zz_6854 = _zz_6855;
  assign _zz_6855 = ($signed(_zz_6856) >>> _zz_580);
  assign _zz_6856 = _zz_6857;
  assign _zz_6857 = ($signed(_zz_6859) + $signed(_zz_576));
  assign _zz_6858 = ({9'd0,data_mid_3_35_real} <<< 9);
  assign _zz_6859 = {{9{_zz_6858[26]}}, _zz_6858};
  assign _zz_6860 = fixTo_694_dout;
  assign _zz_6861 = _zz_6862[35 : 0];
  assign _zz_6862 = _zz_6863;
  assign _zz_6863 = ($signed(_zz_6864) >>> _zz_580);
  assign _zz_6864 = _zz_6865;
  assign _zz_6865 = ($signed(_zz_6867) + $signed(_zz_577));
  assign _zz_6866 = ({9'd0,data_mid_3_35_imag} <<< 9);
  assign _zz_6867 = {{9{_zz_6866[26]}}, _zz_6866};
  assign _zz_6868 = fixTo_695_dout;
  assign _zz_6869 = ($signed(twiddle_factor_table_11_real) + $signed(twiddle_factor_table_11_imag));
  assign _zz_6870 = ($signed(_zz_583) - $signed(_zz_6871));
  assign _zz_6871 = ($signed(_zz_6872) * $signed(twiddle_factor_table_11_imag));
  assign _zz_6872 = ($signed(data_mid_3_44_real) + $signed(data_mid_3_44_imag));
  assign _zz_6873 = fixTo_696_dout;
  assign _zz_6874 = ($signed(_zz_583) + $signed(_zz_6875));
  assign _zz_6875 = ($signed(_zz_6876) * $signed(twiddle_factor_table_11_real));
  assign _zz_6876 = ($signed(data_mid_3_44_imag) - $signed(data_mid_3_44_real));
  assign _zz_6877 = fixTo_697_dout;
  assign _zz_6878 = _zz_6879[35 : 0];
  assign _zz_6879 = _zz_6880;
  assign _zz_6880 = ($signed(_zz_6881) >>> _zz_584);
  assign _zz_6881 = _zz_6882;
  assign _zz_6882 = ($signed(_zz_6884) - $signed(_zz_581));
  assign _zz_6883 = ({9'd0,data_mid_3_36_real} <<< 9);
  assign _zz_6884 = {{9{_zz_6883[26]}}, _zz_6883};
  assign _zz_6885 = fixTo_698_dout;
  assign _zz_6886 = _zz_6887[35 : 0];
  assign _zz_6887 = _zz_6888;
  assign _zz_6888 = ($signed(_zz_6889) >>> _zz_584);
  assign _zz_6889 = _zz_6890;
  assign _zz_6890 = ($signed(_zz_6892) - $signed(_zz_582));
  assign _zz_6891 = ({9'd0,data_mid_3_36_imag} <<< 9);
  assign _zz_6892 = {{9{_zz_6891[26]}}, _zz_6891};
  assign _zz_6893 = fixTo_699_dout;
  assign _zz_6894 = _zz_6895[35 : 0];
  assign _zz_6895 = _zz_6896;
  assign _zz_6896 = ($signed(_zz_6897) >>> _zz_585);
  assign _zz_6897 = _zz_6898;
  assign _zz_6898 = ($signed(_zz_6900) + $signed(_zz_581));
  assign _zz_6899 = ({9'd0,data_mid_3_36_real} <<< 9);
  assign _zz_6900 = {{9{_zz_6899[26]}}, _zz_6899};
  assign _zz_6901 = fixTo_700_dout;
  assign _zz_6902 = _zz_6903[35 : 0];
  assign _zz_6903 = _zz_6904;
  assign _zz_6904 = ($signed(_zz_6905) >>> _zz_585);
  assign _zz_6905 = _zz_6906;
  assign _zz_6906 = ($signed(_zz_6908) + $signed(_zz_582));
  assign _zz_6907 = ({9'd0,data_mid_3_36_imag} <<< 9);
  assign _zz_6908 = {{9{_zz_6907[26]}}, _zz_6907};
  assign _zz_6909 = fixTo_701_dout;
  assign _zz_6910 = ($signed(twiddle_factor_table_12_real) + $signed(twiddle_factor_table_12_imag));
  assign _zz_6911 = ($signed(_zz_588) - $signed(_zz_6912));
  assign _zz_6912 = ($signed(_zz_6913) * $signed(twiddle_factor_table_12_imag));
  assign _zz_6913 = ($signed(data_mid_3_45_real) + $signed(data_mid_3_45_imag));
  assign _zz_6914 = fixTo_702_dout;
  assign _zz_6915 = ($signed(_zz_588) + $signed(_zz_6916));
  assign _zz_6916 = ($signed(_zz_6917) * $signed(twiddle_factor_table_12_real));
  assign _zz_6917 = ($signed(data_mid_3_45_imag) - $signed(data_mid_3_45_real));
  assign _zz_6918 = fixTo_703_dout;
  assign _zz_6919 = _zz_6920[35 : 0];
  assign _zz_6920 = _zz_6921;
  assign _zz_6921 = ($signed(_zz_6922) >>> _zz_589);
  assign _zz_6922 = _zz_6923;
  assign _zz_6923 = ($signed(_zz_6925) - $signed(_zz_586));
  assign _zz_6924 = ({9'd0,data_mid_3_37_real} <<< 9);
  assign _zz_6925 = {{9{_zz_6924[26]}}, _zz_6924};
  assign _zz_6926 = fixTo_704_dout;
  assign _zz_6927 = _zz_6928[35 : 0];
  assign _zz_6928 = _zz_6929;
  assign _zz_6929 = ($signed(_zz_6930) >>> _zz_589);
  assign _zz_6930 = _zz_6931;
  assign _zz_6931 = ($signed(_zz_6933) - $signed(_zz_587));
  assign _zz_6932 = ({9'd0,data_mid_3_37_imag} <<< 9);
  assign _zz_6933 = {{9{_zz_6932[26]}}, _zz_6932};
  assign _zz_6934 = fixTo_705_dout;
  assign _zz_6935 = _zz_6936[35 : 0];
  assign _zz_6936 = _zz_6937;
  assign _zz_6937 = ($signed(_zz_6938) >>> _zz_590);
  assign _zz_6938 = _zz_6939;
  assign _zz_6939 = ($signed(_zz_6941) + $signed(_zz_586));
  assign _zz_6940 = ({9'd0,data_mid_3_37_real} <<< 9);
  assign _zz_6941 = {{9{_zz_6940[26]}}, _zz_6940};
  assign _zz_6942 = fixTo_706_dout;
  assign _zz_6943 = _zz_6944[35 : 0];
  assign _zz_6944 = _zz_6945;
  assign _zz_6945 = ($signed(_zz_6946) >>> _zz_590);
  assign _zz_6946 = _zz_6947;
  assign _zz_6947 = ($signed(_zz_6949) + $signed(_zz_587));
  assign _zz_6948 = ({9'd0,data_mid_3_37_imag} <<< 9);
  assign _zz_6949 = {{9{_zz_6948[26]}}, _zz_6948};
  assign _zz_6950 = fixTo_707_dout;
  assign _zz_6951 = ($signed(twiddle_factor_table_13_real) + $signed(twiddle_factor_table_13_imag));
  assign _zz_6952 = ($signed(_zz_593) - $signed(_zz_6953));
  assign _zz_6953 = ($signed(_zz_6954) * $signed(twiddle_factor_table_13_imag));
  assign _zz_6954 = ($signed(data_mid_3_46_real) + $signed(data_mid_3_46_imag));
  assign _zz_6955 = fixTo_708_dout;
  assign _zz_6956 = ($signed(_zz_593) + $signed(_zz_6957));
  assign _zz_6957 = ($signed(_zz_6958) * $signed(twiddle_factor_table_13_real));
  assign _zz_6958 = ($signed(data_mid_3_46_imag) - $signed(data_mid_3_46_real));
  assign _zz_6959 = fixTo_709_dout;
  assign _zz_6960 = _zz_6961[35 : 0];
  assign _zz_6961 = _zz_6962;
  assign _zz_6962 = ($signed(_zz_6963) >>> _zz_594);
  assign _zz_6963 = _zz_6964;
  assign _zz_6964 = ($signed(_zz_6966) - $signed(_zz_591));
  assign _zz_6965 = ({9'd0,data_mid_3_38_real} <<< 9);
  assign _zz_6966 = {{9{_zz_6965[26]}}, _zz_6965};
  assign _zz_6967 = fixTo_710_dout;
  assign _zz_6968 = _zz_6969[35 : 0];
  assign _zz_6969 = _zz_6970;
  assign _zz_6970 = ($signed(_zz_6971) >>> _zz_594);
  assign _zz_6971 = _zz_6972;
  assign _zz_6972 = ($signed(_zz_6974) - $signed(_zz_592));
  assign _zz_6973 = ({9'd0,data_mid_3_38_imag} <<< 9);
  assign _zz_6974 = {{9{_zz_6973[26]}}, _zz_6973};
  assign _zz_6975 = fixTo_711_dout;
  assign _zz_6976 = _zz_6977[35 : 0];
  assign _zz_6977 = _zz_6978;
  assign _zz_6978 = ($signed(_zz_6979) >>> _zz_595);
  assign _zz_6979 = _zz_6980;
  assign _zz_6980 = ($signed(_zz_6982) + $signed(_zz_591));
  assign _zz_6981 = ({9'd0,data_mid_3_38_real} <<< 9);
  assign _zz_6982 = {{9{_zz_6981[26]}}, _zz_6981};
  assign _zz_6983 = fixTo_712_dout;
  assign _zz_6984 = _zz_6985[35 : 0];
  assign _zz_6985 = _zz_6986;
  assign _zz_6986 = ($signed(_zz_6987) >>> _zz_595);
  assign _zz_6987 = _zz_6988;
  assign _zz_6988 = ($signed(_zz_6990) + $signed(_zz_592));
  assign _zz_6989 = ({9'd0,data_mid_3_38_imag} <<< 9);
  assign _zz_6990 = {{9{_zz_6989[26]}}, _zz_6989};
  assign _zz_6991 = fixTo_713_dout;
  assign _zz_6992 = ($signed(twiddle_factor_table_14_real) + $signed(twiddle_factor_table_14_imag));
  assign _zz_6993 = ($signed(_zz_598) - $signed(_zz_6994));
  assign _zz_6994 = ($signed(_zz_6995) * $signed(twiddle_factor_table_14_imag));
  assign _zz_6995 = ($signed(data_mid_3_47_real) + $signed(data_mid_3_47_imag));
  assign _zz_6996 = fixTo_714_dout;
  assign _zz_6997 = ($signed(_zz_598) + $signed(_zz_6998));
  assign _zz_6998 = ($signed(_zz_6999) * $signed(twiddle_factor_table_14_real));
  assign _zz_6999 = ($signed(data_mid_3_47_imag) - $signed(data_mid_3_47_real));
  assign _zz_7000 = fixTo_715_dout;
  assign _zz_7001 = _zz_7002[35 : 0];
  assign _zz_7002 = _zz_7003;
  assign _zz_7003 = ($signed(_zz_7004) >>> _zz_599);
  assign _zz_7004 = _zz_7005;
  assign _zz_7005 = ($signed(_zz_7007) - $signed(_zz_596));
  assign _zz_7006 = ({9'd0,data_mid_3_39_real} <<< 9);
  assign _zz_7007 = {{9{_zz_7006[26]}}, _zz_7006};
  assign _zz_7008 = fixTo_716_dout;
  assign _zz_7009 = _zz_7010[35 : 0];
  assign _zz_7010 = _zz_7011;
  assign _zz_7011 = ($signed(_zz_7012) >>> _zz_599);
  assign _zz_7012 = _zz_7013;
  assign _zz_7013 = ($signed(_zz_7015) - $signed(_zz_597));
  assign _zz_7014 = ({9'd0,data_mid_3_39_imag} <<< 9);
  assign _zz_7015 = {{9{_zz_7014[26]}}, _zz_7014};
  assign _zz_7016 = fixTo_717_dout;
  assign _zz_7017 = _zz_7018[35 : 0];
  assign _zz_7018 = _zz_7019;
  assign _zz_7019 = ($signed(_zz_7020) >>> _zz_600);
  assign _zz_7020 = _zz_7021;
  assign _zz_7021 = ($signed(_zz_7023) + $signed(_zz_596));
  assign _zz_7022 = ({9'd0,data_mid_3_39_real} <<< 9);
  assign _zz_7023 = {{9{_zz_7022[26]}}, _zz_7022};
  assign _zz_7024 = fixTo_718_dout;
  assign _zz_7025 = _zz_7026[35 : 0];
  assign _zz_7026 = _zz_7027;
  assign _zz_7027 = ($signed(_zz_7028) >>> _zz_600);
  assign _zz_7028 = _zz_7029;
  assign _zz_7029 = ($signed(_zz_7031) + $signed(_zz_597));
  assign _zz_7030 = ({9'd0,data_mid_3_39_imag} <<< 9);
  assign _zz_7031 = {{9{_zz_7030[26]}}, _zz_7030};
  assign _zz_7032 = fixTo_719_dout;
  assign _zz_7033 = ($signed(twiddle_factor_table_7_real) + $signed(twiddle_factor_table_7_imag));
  assign _zz_7034 = ($signed(_zz_603) - $signed(_zz_7035));
  assign _zz_7035 = ($signed(_zz_7036) * $signed(twiddle_factor_table_7_imag));
  assign _zz_7036 = ($signed(data_mid_3_56_real) + $signed(data_mid_3_56_imag));
  assign _zz_7037 = fixTo_720_dout;
  assign _zz_7038 = ($signed(_zz_603) + $signed(_zz_7039));
  assign _zz_7039 = ($signed(_zz_7040) * $signed(twiddle_factor_table_7_real));
  assign _zz_7040 = ($signed(data_mid_3_56_imag) - $signed(data_mid_3_56_real));
  assign _zz_7041 = fixTo_721_dout;
  assign _zz_7042 = _zz_7043[35 : 0];
  assign _zz_7043 = _zz_7044;
  assign _zz_7044 = ($signed(_zz_7045) >>> _zz_604);
  assign _zz_7045 = _zz_7046;
  assign _zz_7046 = ($signed(_zz_7048) - $signed(_zz_601));
  assign _zz_7047 = ({9'd0,data_mid_3_48_real} <<< 9);
  assign _zz_7048 = {{9{_zz_7047[26]}}, _zz_7047};
  assign _zz_7049 = fixTo_722_dout;
  assign _zz_7050 = _zz_7051[35 : 0];
  assign _zz_7051 = _zz_7052;
  assign _zz_7052 = ($signed(_zz_7053) >>> _zz_604);
  assign _zz_7053 = _zz_7054;
  assign _zz_7054 = ($signed(_zz_7056) - $signed(_zz_602));
  assign _zz_7055 = ({9'd0,data_mid_3_48_imag} <<< 9);
  assign _zz_7056 = {{9{_zz_7055[26]}}, _zz_7055};
  assign _zz_7057 = fixTo_723_dout;
  assign _zz_7058 = _zz_7059[35 : 0];
  assign _zz_7059 = _zz_7060;
  assign _zz_7060 = ($signed(_zz_7061) >>> _zz_605);
  assign _zz_7061 = _zz_7062;
  assign _zz_7062 = ($signed(_zz_7064) + $signed(_zz_601));
  assign _zz_7063 = ({9'd0,data_mid_3_48_real} <<< 9);
  assign _zz_7064 = {{9{_zz_7063[26]}}, _zz_7063};
  assign _zz_7065 = fixTo_724_dout;
  assign _zz_7066 = _zz_7067[35 : 0];
  assign _zz_7067 = _zz_7068;
  assign _zz_7068 = ($signed(_zz_7069) >>> _zz_605);
  assign _zz_7069 = _zz_7070;
  assign _zz_7070 = ($signed(_zz_7072) + $signed(_zz_602));
  assign _zz_7071 = ({9'd0,data_mid_3_48_imag} <<< 9);
  assign _zz_7072 = {{9{_zz_7071[26]}}, _zz_7071};
  assign _zz_7073 = fixTo_725_dout;
  assign _zz_7074 = ($signed(twiddle_factor_table_8_real) + $signed(twiddle_factor_table_8_imag));
  assign _zz_7075 = ($signed(_zz_608) - $signed(_zz_7076));
  assign _zz_7076 = ($signed(_zz_7077) * $signed(twiddle_factor_table_8_imag));
  assign _zz_7077 = ($signed(data_mid_3_57_real) + $signed(data_mid_3_57_imag));
  assign _zz_7078 = fixTo_726_dout;
  assign _zz_7079 = ($signed(_zz_608) + $signed(_zz_7080));
  assign _zz_7080 = ($signed(_zz_7081) * $signed(twiddle_factor_table_8_real));
  assign _zz_7081 = ($signed(data_mid_3_57_imag) - $signed(data_mid_3_57_real));
  assign _zz_7082 = fixTo_727_dout;
  assign _zz_7083 = _zz_7084[35 : 0];
  assign _zz_7084 = _zz_7085;
  assign _zz_7085 = ($signed(_zz_7086) >>> _zz_609);
  assign _zz_7086 = _zz_7087;
  assign _zz_7087 = ($signed(_zz_7089) - $signed(_zz_606));
  assign _zz_7088 = ({9'd0,data_mid_3_49_real} <<< 9);
  assign _zz_7089 = {{9{_zz_7088[26]}}, _zz_7088};
  assign _zz_7090 = fixTo_728_dout;
  assign _zz_7091 = _zz_7092[35 : 0];
  assign _zz_7092 = _zz_7093;
  assign _zz_7093 = ($signed(_zz_7094) >>> _zz_609);
  assign _zz_7094 = _zz_7095;
  assign _zz_7095 = ($signed(_zz_7097) - $signed(_zz_607));
  assign _zz_7096 = ({9'd0,data_mid_3_49_imag} <<< 9);
  assign _zz_7097 = {{9{_zz_7096[26]}}, _zz_7096};
  assign _zz_7098 = fixTo_729_dout;
  assign _zz_7099 = _zz_7100[35 : 0];
  assign _zz_7100 = _zz_7101;
  assign _zz_7101 = ($signed(_zz_7102) >>> _zz_610);
  assign _zz_7102 = _zz_7103;
  assign _zz_7103 = ($signed(_zz_7105) + $signed(_zz_606));
  assign _zz_7104 = ({9'd0,data_mid_3_49_real} <<< 9);
  assign _zz_7105 = {{9{_zz_7104[26]}}, _zz_7104};
  assign _zz_7106 = fixTo_730_dout;
  assign _zz_7107 = _zz_7108[35 : 0];
  assign _zz_7108 = _zz_7109;
  assign _zz_7109 = ($signed(_zz_7110) >>> _zz_610);
  assign _zz_7110 = _zz_7111;
  assign _zz_7111 = ($signed(_zz_7113) + $signed(_zz_607));
  assign _zz_7112 = ({9'd0,data_mid_3_49_imag} <<< 9);
  assign _zz_7113 = {{9{_zz_7112[26]}}, _zz_7112};
  assign _zz_7114 = fixTo_731_dout;
  assign _zz_7115 = ($signed(twiddle_factor_table_9_real) + $signed(twiddle_factor_table_9_imag));
  assign _zz_7116 = ($signed(_zz_613) - $signed(_zz_7117));
  assign _zz_7117 = ($signed(_zz_7118) * $signed(twiddle_factor_table_9_imag));
  assign _zz_7118 = ($signed(data_mid_3_58_real) + $signed(data_mid_3_58_imag));
  assign _zz_7119 = fixTo_732_dout;
  assign _zz_7120 = ($signed(_zz_613) + $signed(_zz_7121));
  assign _zz_7121 = ($signed(_zz_7122) * $signed(twiddle_factor_table_9_real));
  assign _zz_7122 = ($signed(data_mid_3_58_imag) - $signed(data_mid_3_58_real));
  assign _zz_7123 = fixTo_733_dout;
  assign _zz_7124 = _zz_7125[35 : 0];
  assign _zz_7125 = _zz_7126;
  assign _zz_7126 = ($signed(_zz_7127) >>> _zz_614);
  assign _zz_7127 = _zz_7128;
  assign _zz_7128 = ($signed(_zz_7130) - $signed(_zz_611));
  assign _zz_7129 = ({9'd0,data_mid_3_50_real} <<< 9);
  assign _zz_7130 = {{9{_zz_7129[26]}}, _zz_7129};
  assign _zz_7131 = fixTo_734_dout;
  assign _zz_7132 = _zz_7133[35 : 0];
  assign _zz_7133 = _zz_7134;
  assign _zz_7134 = ($signed(_zz_7135) >>> _zz_614);
  assign _zz_7135 = _zz_7136;
  assign _zz_7136 = ($signed(_zz_7138) - $signed(_zz_612));
  assign _zz_7137 = ({9'd0,data_mid_3_50_imag} <<< 9);
  assign _zz_7138 = {{9{_zz_7137[26]}}, _zz_7137};
  assign _zz_7139 = fixTo_735_dout;
  assign _zz_7140 = _zz_7141[35 : 0];
  assign _zz_7141 = _zz_7142;
  assign _zz_7142 = ($signed(_zz_7143) >>> _zz_615);
  assign _zz_7143 = _zz_7144;
  assign _zz_7144 = ($signed(_zz_7146) + $signed(_zz_611));
  assign _zz_7145 = ({9'd0,data_mid_3_50_real} <<< 9);
  assign _zz_7146 = {{9{_zz_7145[26]}}, _zz_7145};
  assign _zz_7147 = fixTo_736_dout;
  assign _zz_7148 = _zz_7149[35 : 0];
  assign _zz_7149 = _zz_7150;
  assign _zz_7150 = ($signed(_zz_7151) >>> _zz_615);
  assign _zz_7151 = _zz_7152;
  assign _zz_7152 = ($signed(_zz_7154) + $signed(_zz_612));
  assign _zz_7153 = ({9'd0,data_mid_3_50_imag} <<< 9);
  assign _zz_7154 = {{9{_zz_7153[26]}}, _zz_7153};
  assign _zz_7155 = fixTo_737_dout;
  assign _zz_7156 = ($signed(twiddle_factor_table_10_real) + $signed(twiddle_factor_table_10_imag));
  assign _zz_7157 = ($signed(_zz_618) - $signed(_zz_7158));
  assign _zz_7158 = ($signed(_zz_7159) * $signed(twiddle_factor_table_10_imag));
  assign _zz_7159 = ($signed(data_mid_3_59_real) + $signed(data_mid_3_59_imag));
  assign _zz_7160 = fixTo_738_dout;
  assign _zz_7161 = ($signed(_zz_618) + $signed(_zz_7162));
  assign _zz_7162 = ($signed(_zz_7163) * $signed(twiddle_factor_table_10_real));
  assign _zz_7163 = ($signed(data_mid_3_59_imag) - $signed(data_mid_3_59_real));
  assign _zz_7164 = fixTo_739_dout;
  assign _zz_7165 = _zz_7166[35 : 0];
  assign _zz_7166 = _zz_7167;
  assign _zz_7167 = ($signed(_zz_7168) >>> _zz_619);
  assign _zz_7168 = _zz_7169;
  assign _zz_7169 = ($signed(_zz_7171) - $signed(_zz_616));
  assign _zz_7170 = ({9'd0,data_mid_3_51_real} <<< 9);
  assign _zz_7171 = {{9{_zz_7170[26]}}, _zz_7170};
  assign _zz_7172 = fixTo_740_dout;
  assign _zz_7173 = _zz_7174[35 : 0];
  assign _zz_7174 = _zz_7175;
  assign _zz_7175 = ($signed(_zz_7176) >>> _zz_619);
  assign _zz_7176 = _zz_7177;
  assign _zz_7177 = ($signed(_zz_7179) - $signed(_zz_617));
  assign _zz_7178 = ({9'd0,data_mid_3_51_imag} <<< 9);
  assign _zz_7179 = {{9{_zz_7178[26]}}, _zz_7178};
  assign _zz_7180 = fixTo_741_dout;
  assign _zz_7181 = _zz_7182[35 : 0];
  assign _zz_7182 = _zz_7183;
  assign _zz_7183 = ($signed(_zz_7184) >>> _zz_620);
  assign _zz_7184 = _zz_7185;
  assign _zz_7185 = ($signed(_zz_7187) + $signed(_zz_616));
  assign _zz_7186 = ({9'd0,data_mid_3_51_real} <<< 9);
  assign _zz_7187 = {{9{_zz_7186[26]}}, _zz_7186};
  assign _zz_7188 = fixTo_742_dout;
  assign _zz_7189 = _zz_7190[35 : 0];
  assign _zz_7190 = _zz_7191;
  assign _zz_7191 = ($signed(_zz_7192) >>> _zz_620);
  assign _zz_7192 = _zz_7193;
  assign _zz_7193 = ($signed(_zz_7195) + $signed(_zz_617));
  assign _zz_7194 = ({9'd0,data_mid_3_51_imag} <<< 9);
  assign _zz_7195 = {{9{_zz_7194[26]}}, _zz_7194};
  assign _zz_7196 = fixTo_743_dout;
  assign _zz_7197 = ($signed(twiddle_factor_table_11_real) + $signed(twiddle_factor_table_11_imag));
  assign _zz_7198 = ($signed(_zz_623) - $signed(_zz_7199));
  assign _zz_7199 = ($signed(_zz_7200) * $signed(twiddle_factor_table_11_imag));
  assign _zz_7200 = ($signed(data_mid_3_60_real) + $signed(data_mid_3_60_imag));
  assign _zz_7201 = fixTo_744_dout;
  assign _zz_7202 = ($signed(_zz_623) + $signed(_zz_7203));
  assign _zz_7203 = ($signed(_zz_7204) * $signed(twiddle_factor_table_11_real));
  assign _zz_7204 = ($signed(data_mid_3_60_imag) - $signed(data_mid_3_60_real));
  assign _zz_7205 = fixTo_745_dout;
  assign _zz_7206 = _zz_7207[35 : 0];
  assign _zz_7207 = _zz_7208;
  assign _zz_7208 = ($signed(_zz_7209) >>> _zz_624);
  assign _zz_7209 = _zz_7210;
  assign _zz_7210 = ($signed(_zz_7212) - $signed(_zz_621));
  assign _zz_7211 = ({9'd0,data_mid_3_52_real} <<< 9);
  assign _zz_7212 = {{9{_zz_7211[26]}}, _zz_7211};
  assign _zz_7213 = fixTo_746_dout;
  assign _zz_7214 = _zz_7215[35 : 0];
  assign _zz_7215 = _zz_7216;
  assign _zz_7216 = ($signed(_zz_7217) >>> _zz_624);
  assign _zz_7217 = _zz_7218;
  assign _zz_7218 = ($signed(_zz_7220) - $signed(_zz_622));
  assign _zz_7219 = ({9'd0,data_mid_3_52_imag} <<< 9);
  assign _zz_7220 = {{9{_zz_7219[26]}}, _zz_7219};
  assign _zz_7221 = fixTo_747_dout;
  assign _zz_7222 = _zz_7223[35 : 0];
  assign _zz_7223 = _zz_7224;
  assign _zz_7224 = ($signed(_zz_7225) >>> _zz_625);
  assign _zz_7225 = _zz_7226;
  assign _zz_7226 = ($signed(_zz_7228) + $signed(_zz_621));
  assign _zz_7227 = ({9'd0,data_mid_3_52_real} <<< 9);
  assign _zz_7228 = {{9{_zz_7227[26]}}, _zz_7227};
  assign _zz_7229 = fixTo_748_dout;
  assign _zz_7230 = _zz_7231[35 : 0];
  assign _zz_7231 = _zz_7232;
  assign _zz_7232 = ($signed(_zz_7233) >>> _zz_625);
  assign _zz_7233 = _zz_7234;
  assign _zz_7234 = ($signed(_zz_7236) + $signed(_zz_622));
  assign _zz_7235 = ({9'd0,data_mid_3_52_imag} <<< 9);
  assign _zz_7236 = {{9{_zz_7235[26]}}, _zz_7235};
  assign _zz_7237 = fixTo_749_dout;
  assign _zz_7238 = ($signed(twiddle_factor_table_12_real) + $signed(twiddle_factor_table_12_imag));
  assign _zz_7239 = ($signed(_zz_628) - $signed(_zz_7240));
  assign _zz_7240 = ($signed(_zz_7241) * $signed(twiddle_factor_table_12_imag));
  assign _zz_7241 = ($signed(data_mid_3_61_real) + $signed(data_mid_3_61_imag));
  assign _zz_7242 = fixTo_750_dout;
  assign _zz_7243 = ($signed(_zz_628) + $signed(_zz_7244));
  assign _zz_7244 = ($signed(_zz_7245) * $signed(twiddle_factor_table_12_real));
  assign _zz_7245 = ($signed(data_mid_3_61_imag) - $signed(data_mid_3_61_real));
  assign _zz_7246 = fixTo_751_dout;
  assign _zz_7247 = _zz_7248[35 : 0];
  assign _zz_7248 = _zz_7249;
  assign _zz_7249 = ($signed(_zz_7250) >>> _zz_629);
  assign _zz_7250 = _zz_7251;
  assign _zz_7251 = ($signed(_zz_7253) - $signed(_zz_626));
  assign _zz_7252 = ({9'd0,data_mid_3_53_real} <<< 9);
  assign _zz_7253 = {{9{_zz_7252[26]}}, _zz_7252};
  assign _zz_7254 = fixTo_752_dout;
  assign _zz_7255 = _zz_7256[35 : 0];
  assign _zz_7256 = _zz_7257;
  assign _zz_7257 = ($signed(_zz_7258) >>> _zz_629);
  assign _zz_7258 = _zz_7259;
  assign _zz_7259 = ($signed(_zz_7261) - $signed(_zz_627));
  assign _zz_7260 = ({9'd0,data_mid_3_53_imag} <<< 9);
  assign _zz_7261 = {{9{_zz_7260[26]}}, _zz_7260};
  assign _zz_7262 = fixTo_753_dout;
  assign _zz_7263 = _zz_7264[35 : 0];
  assign _zz_7264 = _zz_7265;
  assign _zz_7265 = ($signed(_zz_7266) >>> _zz_630);
  assign _zz_7266 = _zz_7267;
  assign _zz_7267 = ($signed(_zz_7269) + $signed(_zz_626));
  assign _zz_7268 = ({9'd0,data_mid_3_53_real} <<< 9);
  assign _zz_7269 = {{9{_zz_7268[26]}}, _zz_7268};
  assign _zz_7270 = fixTo_754_dout;
  assign _zz_7271 = _zz_7272[35 : 0];
  assign _zz_7272 = _zz_7273;
  assign _zz_7273 = ($signed(_zz_7274) >>> _zz_630);
  assign _zz_7274 = _zz_7275;
  assign _zz_7275 = ($signed(_zz_7277) + $signed(_zz_627));
  assign _zz_7276 = ({9'd0,data_mid_3_53_imag} <<< 9);
  assign _zz_7277 = {{9{_zz_7276[26]}}, _zz_7276};
  assign _zz_7278 = fixTo_755_dout;
  assign _zz_7279 = ($signed(twiddle_factor_table_13_real) + $signed(twiddle_factor_table_13_imag));
  assign _zz_7280 = ($signed(_zz_633) - $signed(_zz_7281));
  assign _zz_7281 = ($signed(_zz_7282) * $signed(twiddle_factor_table_13_imag));
  assign _zz_7282 = ($signed(data_mid_3_62_real) + $signed(data_mid_3_62_imag));
  assign _zz_7283 = fixTo_756_dout;
  assign _zz_7284 = ($signed(_zz_633) + $signed(_zz_7285));
  assign _zz_7285 = ($signed(_zz_7286) * $signed(twiddle_factor_table_13_real));
  assign _zz_7286 = ($signed(data_mid_3_62_imag) - $signed(data_mid_3_62_real));
  assign _zz_7287 = fixTo_757_dout;
  assign _zz_7288 = _zz_7289[35 : 0];
  assign _zz_7289 = _zz_7290;
  assign _zz_7290 = ($signed(_zz_7291) >>> _zz_634);
  assign _zz_7291 = _zz_7292;
  assign _zz_7292 = ($signed(_zz_7294) - $signed(_zz_631));
  assign _zz_7293 = ({9'd0,data_mid_3_54_real} <<< 9);
  assign _zz_7294 = {{9{_zz_7293[26]}}, _zz_7293};
  assign _zz_7295 = fixTo_758_dout;
  assign _zz_7296 = _zz_7297[35 : 0];
  assign _zz_7297 = _zz_7298;
  assign _zz_7298 = ($signed(_zz_7299) >>> _zz_634);
  assign _zz_7299 = _zz_7300;
  assign _zz_7300 = ($signed(_zz_7302) - $signed(_zz_632));
  assign _zz_7301 = ({9'd0,data_mid_3_54_imag} <<< 9);
  assign _zz_7302 = {{9{_zz_7301[26]}}, _zz_7301};
  assign _zz_7303 = fixTo_759_dout;
  assign _zz_7304 = _zz_7305[35 : 0];
  assign _zz_7305 = _zz_7306;
  assign _zz_7306 = ($signed(_zz_7307) >>> _zz_635);
  assign _zz_7307 = _zz_7308;
  assign _zz_7308 = ($signed(_zz_7310) + $signed(_zz_631));
  assign _zz_7309 = ({9'd0,data_mid_3_54_real} <<< 9);
  assign _zz_7310 = {{9{_zz_7309[26]}}, _zz_7309};
  assign _zz_7311 = fixTo_760_dout;
  assign _zz_7312 = _zz_7313[35 : 0];
  assign _zz_7313 = _zz_7314;
  assign _zz_7314 = ($signed(_zz_7315) >>> _zz_635);
  assign _zz_7315 = _zz_7316;
  assign _zz_7316 = ($signed(_zz_7318) + $signed(_zz_632));
  assign _zz_7317 = ({9'd0,data_mid_3_54_imag} <<< 9);
  assign _zz_7318 = {{9{_zz_7317[26]}}, _zz_7317};
  assign _zz_7319 = fixTo_761_dout;
  assign _zz_7320 = ($signed(twiddle_factor_table_14_real) + $signed(twiddle_factor_table_14_imag));
  assign _zz_7321 = ($signed(_zz_638) - $signed(_zz_7322));
  assign _zz_7322 = ($signed(_zz_7323) * $signed(twiddle_factor_table_14_imag));
  assign _zz_7323 = ($signed(data_mid_3_63_real) + $signed(data_mid_3_63_imag));
  assign _zz_7324 = fixTo_762_dout;
  assign _zz_7325 = ($signed(_zz_638) + $signed(_zz_7326));
  assign _zz_7326 = ($signed(_zz_7327) * $signed(twiddle_factor_table_14_real));
  assign _zz_7327 = ($signed(data_mid_3_63_imag) - $signed(data_mid_3_63_real));
  assign _zz_7328 = fixTo_763_dout;
  assign _zz_7329 = _zz_7330[35 : 0];
  assign _zz_7330 = _zz_7331;
  assign _zz_7331 = ($signed(_zz_7332) >>> _zz_639);
  assign _zz_7332 = _zz_7333;
  assign _zz_7333 = ($signed(_zz_7335) - $signed(_zz_636));
  assign _zz_7334 = ({9'd0,data_mid_3_55_real} <<< 9);
  assign _zz_7335 = {{9{_zz_7334[26]}}, _zz_7334};
  assign _zz_7336 = fixTo_764_dout;
  assign _zz_7337 = _zz_7338[35 : 0];
  assign _zz_7338 = _zz_7339;
  assign _zz_7339 = ($signed(_zz_7340) >>> _zz_639);
  assign _zz_7340 = _zz_7341;
  assign _zz_7341 = ($signed(_zz_7343) - $signed(_zz_637));
  assign _zz_7342 = ({9'd0,data_mid_3_55_imag} <<< 9);
  assign _zz_7343 = {{9{_zz_7342[26]}}, _zz_7342};
  assign _zz_7344 = fixTo_765_dout;
  assign _zz_7345 = _zz_7346[35 : 0];
  assign _zz_7346 = _zz_7347;
  assign _zz_7347 = ($signed(_zz_7348) >>> _zz_640);
  assign _zz_7348 = _zz_7349;
  assign _zz_7349 = ($signed(_zz_7351) + $signed(_zz_636));
  assign _zz_7350 = ({9'd0,data_mid_3_55_real} <<< 9);
  assign _zz_7351 = {{9{_zz_7350[26]}}, _zz_7350};
  assign _zz_7352 = fixTo_766_dout;
  assign _zz_7353 = _zz_7354[35 : 0];
  assign _zz_7354 = _zz_7355;
  assign _zz_7355 = ($signed(_zz_7356) >>> _zz_640);
  assign _zz_7356 = _zz_7357;
  assign _zz_7357 = ($signed(_zz_7359) + $signed(_zz_637));
  assign _zz_7358 = ({9'd0,data_mid_3_55_imag} <<< 9);
  assign _zz_7359 = {{9{_zz_7358[26]}}, _zz_7358};
  assign _zz_7360 = fixTo_767_dout;
  assign _zz_7361 = ($signed(twiddle_factor_table_15_real) + $signed(twiddle_factor_table_15_imag));
  assign _zz_7362 = ($signed(_zz_643) - $signed(_zz_7363));
  assign _zz_7363 = ($signed(_zz_7364) * $signed(twiddle_factor_table_15_imag));
  assign _zz_7364 = ($signed(data_mid_4_16_real) + $signed(data_mid_4_16_imag));
  assign _zz_7365 = fixTo_768_dout;
  assign _zz_7366 = ($signed(_zz_643) + $signed(_zz_7367));
  assign _zz_7367 = ($signed(_zz_7368) * $signed(twiddle_factor_table_15_real));
  assign _zz_7368 = ($signed(data_mid_4_16_imag) - $signed(data_mid_4_16_real));
  assign _zz_7369 = fixTo_769_dout;
  assign _zz_7370 = _zz_7371[35 : 0];
  assign _zz_7371 = _zz_7372;
  assign _zz_7372 = ($signed(_zz_7373) >>> _zz_644);
  assign _zz_7373 = _zz_7374;
  assign _zz_7374 = ($signed(_zz_7376) - $signed(_zz_641));
  assign _zz_7375 = ({9'd0,data_mid_4_0_real} <<< 9);
  assign _zz_7376 = {{9{_zz_7375[26]}}, _zz_7375};
  assign _zz_7377 = fixTo_770_dout;
  assign _zz_7378 = _zz_7379[35 : 0];
  assign _zz_7379 = _zz_7380;
  assign _zz_7380 = ($signed(_zz_7381) >>> _zz_644);
  assign _zz_7381 = _zz_7382;
  assign _zz_7382 = ($signed(_zz_7384) - $signed(_zz_642));
  assign _zz_7383 = ({9'd0,data_mid_4_0_imag} <<< 9);
  assign _zz_7384 = {{9{_zz_7383[26]}}, _zz_7383};
  assign _zz_7385 = fixTo_771_dout;
  assign _zz_7386 = _zz_7387[35 : 0];
  assign _zz_7387 = _zz_7388;
  assign _zz_7388 = ($signed(_zz_7389) >>> _zz_645);
  assign _zz_7389 = _zz_7390;
  assign _zz_7390 = ($signed(_zz_7392) + $signed(_zz_641));
  assign _zz_7391 = ({9'd0,data_mid_4_0_real} <<< 9);
  assign _zz_7392 = {{9{_zz_7391[26]}}, _zz_7391};
  assign _zz_7393 = fixTo_772_dout;
  assign _zz_7394 = _zz_7395[35 : 0];
  assign _zz_7395 = _zz_7396;
  assign _zz_7396 = ($signed(_zz_7397) >>> _zz_645);
  assign _zz_7397 = _zz_7398;
  assign _zz_7398 = ($signed(_zz_7400) + $signed(_zz_642));
  assign _zz_7399 = ({9'd0,data_mid_4_0_imag} <<< 9);
  assign _zz_7400 = {{9{_zz_7399[26]}}, _zz_7399};
  assign _zz_7401 = fixTo_773_dout;
  assign _zz_7402 = ($signed(twiddle_factor_table_16_real) + $signed(twiddle_factor_table_16_imag));
  assign _zz_7403 = ($signed(_zz_648) - $signed(_zz_7404));
  assign _zz_7404 = ($signed(_zz_7405) * $signed(twiddle_factor_table_16_imag));
  assign _zz_7405 = ($signed(data_mid_4_17_real) + $signed(data_mid_4_17_imag));
  assign _zz_7406 = fixTo_774_dout;
  assign _zz_7407 = ($signed(_zz_648) + $signed(_zz_7408));
  assign _zz_7408 = ($signed(_zz_7409) * $signed(twiddle_factor_table_16_real));
  assign _zz_7409 = ($signed(data_mid_4_17_imag) - $signed(data_mid_4_17_real));
  assign _zz_7410 = fixTo_775_dout;
  assign _zz_7411 = _zz_7412[35 : 0];
  assign _zz_7412 = _zz_7413;
  assign _zz_7413 = ($signed(_zz_7414) >>> _zz_649);
  assign _zz_7414 = _zz_7415;
  assign _zz_7415 = ($signed(_zz_7417) - $signed(_zz_646));
  assign _zz_7416 = ({9'd0,data_mid_4_1_real} <<< 9);
  assign _zz_7417 = {{9{_zz_7416[26]}}, _zz_7416};
  assign _zz_7418 = fixTo_776_dout;
  assign _zz_7419 = _zz_7420[35 : 0];
  assign _zz_7420 = _zz_7421;
  assign _zz_7421 = ($signed(_zz_7422) >>> _zz_649);
  assign _zz_7422 = _zz_7423;
  assign _zz_7423 = ($signed(_zz_7425) - $signed(_zz_647));
  assign _zz_7424 = ({9'd0,data_mid_4_1_imag} <<< 9);
  assign _zz_7425 = {{9{_zz_7424[26]}}, _zz_7424};
  assign _zz_7426 = fixTo_777_dout;
  assign _zz_7427 = _zz_7428[35 : 0];
  assign _zz_7428 = _zz_7429;
  assign _zz_7429 = ($signed(_zz_7430) >>> _zz_650);
  assign _zz_7430 = _zz_7431;
  assign _zz_7431 = ($signed(_zz_7433) + $signed(_zz_646));
  assign _zz_7432 = ({9'd0,data_mid_4_1_real} <<< 9);
  assign _zz_7433 = {{9{_zz_7432[26]}}, _zz_7432};
  assign _zz_7434 = fixTo_778_dout;
  assign _zz_7435 = _zz_7436[35 : 0];
  assign _zz_7436 = _zz_7437;
  assign _zz_7437 = ($signed(_zz_7438) >>> _zz_650);
  assign _zz_7438 = _zz_7439;
  assign _zz_7439 = ($signed(_zz_7441) + $signed(_zz_647));
  assign _zz_7440 = ({9'd0,data_mid_4_1_imag} <<< 9);
  assign _zz_7441 = {{9{_zz_7440[26]}}, _zz_7440};
  assign _zz_7442 = fixTo_779_dout;
  assign _zz_7443 = ($signed(twiddle_factor_table_17_real) + $signed(twiddle_factor_table_17_imag));
  assign _zz_7444 = ($signed(_zz_653) - $signed(_zz_7445));
  assign _zz_7445 = ($signed(_zz_7446) * $signed(twiddle_factor_table_17_imag));
  assign _zz_7446 = ($signed(data_mid_4_18_real) + $signed(data_mid_4_18_imag));
  assign _zz_7447 = fixTo_780_dout;
  assign _zz_7448 = ($signed(_zz_653) + $signed(_zz_7449));
  assign _zz_7449 = ($signed(_zz_7450) * $signed(twiddle_factor_table_17_real));
  assign _zz_7450 = ($signed(data_mid_4_18_imag) - $signed(data_mid_4_18_real));
  assign _zz_7451 = fixTo_781_dout;
  assign _zz_7452 = _zz_7453[35 : 0];
  assign _zz_7453 = _zz_7454;
  assign _zz_7454 = ($signed(_zz_7455) >>> _zz_654);
  assign _zz_7455 = _zz_7456;
  assign _zz_7456 = ($signed(_zz_7458) - $signed(_zz_651));
  assign _zz_7457 = ({9'd0,data_mid_4_2_real} <<< 9);
  assign _zz_7458 = {{9{_zz_7457[26]}}, _zz_7457};
  assign _zz_7459 = fixTo_782_dout;
  assign _zz_7460 = _zz_7461[35 : 0];
  assign _zz_7461 = _zz_7462;
  assign _zz_7462 = ($signed(_zz_7463) >>> _zz_654);
  assign _zz_7463 = _zz_7464;
  assign _zz_7464 = ($signed(_zz_7466) - $signed(_zz_652));
  assign _zz_7465 = ({9'd0,data_mid_4_2_imag} <<< 9);
  assign _zz_7466 = {{9{_zz_7465[26]}}, _zz_7465};
  assign _zz_7467 = fixTo_783_dout;
  assign _zz_7468 = _zz_7469[35 : 0];
  assign _zz_7469 = _zz_7470;
  assign _zz_7470 = ($signed(_zz_7471) >>> _zz_655);
  assign _zz_7471 = _zz_7472;
  assign _zz_7472 = ($signed(_zz_7474) + $signed(_zz_651));
  assign _zz_7473 = ({9'd0,data_mid_4_2_real} <<< 9);
  assign _zz_7474 = {{9{_zz_7473[26]}}, _zz_7473};
  assign _zz_7475 = fixTo_784_dout;
  assign _zz_7476 = _zz_7477[35 : 0];
  assign _zz_7477 = _zz_7478;
  assign _zz_7478 = ($signed(_zz_7479) >>> _zz_655);
  assign _zz_7479 = _zz_7480;
  assign _zz_7480 = ($signed(_zz_7482) + $signed(_zz_652));
  assign _zz_7481 = ({9'd0,data_mid_4_2_imag} <<< 9);
  assign _zz_7482 = {{9{_zz_7481[26]}}, _zz_7481};
  assign _zz_7483 = fixTo_785_dout;
  assign _zz_7484 = ($signed(twiddle_factor_table_18_real) + $signed(twiddle_factor_table_18_imag));
  assign _zz_7485 = ($signed(_zz_658) - $signed(_zz_7486));
  assign _zz_7486 = ($signed(_zz_7487) * $signed(twiddle_factor_table_18_imag));
  assign _zz_7487 = ($signed(data_mid_4_19_real) + $signed(data_mid_4_19_imag));
  assign _zz_7488 = fixTo_786_dout;
  assign _zz_7489 = ($signed(_zz_658) + $signed(_zz_7490));
  assign _zz_7490 = ($signed(_zz_7491) * $signed(twiddle_factor_table_18_real));
  assign _zz_7491 = ($signed(data_mid_4_19_imag) - $signed(data_mid_4_19_real));
  assign _zz_7492 = fixTo_787_dout;
  assign _zz_7493 = _zz_7494[35 : 0];
  assign _zz_7494 = _zz_7495;
  assign _zz_7495 = ($signed(_zz_7496) >>> _zz_659);
  assign _zz_7496 = _zz_7497;
  assign _zz_7497 = ($signed(_zz_7499) - $signed(_zz_656));
  assign _zz_7498 = ({9'd0,data_mid_4_3_real} <<< 9);
  assign _zz_7499 = {{9{_zz_7498[26]}}, _zz_7498};
  assign _zz_7500 = fixTo_788_dout;
  assign _zz_7501 = _zz_7502[35 : 0];
  assign _zz_7502 = _zz_7503;
  assign _zz_7503 = ($signed(_zz_7504) >>> _zz_659);
  assign _zz_7504 = _zz_7505;
  assign _zz_7505 = ($signed(_zz_7507) - $signed(_zz_657));
  assign _zz_7506 = ({9'd0,data_mid_4_3_imag} <<< 9);
  assign _zz_7507 = {{9{_zz_7506[26]}}, _zz_7506};
  assign _zz_7508 = fixTo_789_dout;
  assign _zz_7509 = _zz_7510[35 : 0];
  assign _zz_7510 = _zz_7511;
  assign _zz_7511 = ($signed(_zz_7512) >>> _zz_660);
  assign _zz_7512 = _zz_7513;
  assign _zz_7513 = ($signed(_zz_7515) + $signed(_zz_656));
  assign _zz_7514 = ({9'd0,data_mid_4_3_real} <<< 9);
  assign _zz_7515 = {{9{_zz_7514[26]}}, _zz_7514};
  assign _zz_7516 = fixTo_790_dout;
  assign _zz_7517 = _zz_7518[35 : 0];
  assign _zz_7518 = _zz_7519;
  assign _zz_7519 = ($signed(_zz_7520) >>> _zz_660);
  assign _zz_7520 = _zz_7521;
  assign _zz_7521 = ($signed(_zz_7523) + $signed(_zz_657));
  assign _zz_7522 = ({9'd0,data_mid_4_3_imag} <<< 9);
  assign _zz_7523 = {{9{_zz_7522[26]}}, _zz_7522};
  assign _zz_7524 = fixTo_791_dout;
  assign _zz_7525 = ($signed(twiddle_factor_table_19_real) + $signed(twiddle_factor_table_19_imag));
  assign _zz_7526 = ($signed(_zz_663) - $signed(_zz_7527));
  assign _zz_7527 = ($signed(_zz_7528) * $signed(twiddle_factor_table_19_imag));
  assign _zz_7528 = ($signed(data_mid_4_20_real) + $signed(data_mid_4_20_imag));
  assign _zz_7529 = fixTo_792_dout;
  assign _zz_7530 = ($signed(_zz_663) + $signed(_zz_7531));
  assign _zz_7531 = ($signed(_zz_7532) * $signed(twiddle_factor_table_19_real));
  assign _zz_7532 = ($signed(data_mid_4_20_imag) - $signed(data_mid_4_20_real));
  assign _zz_7533 = fixTo_793_dout;
  assign _zz_7534 = _zz_7535[35 : 0];
  assign _zz_7535 = _zz_7536;
  assign _zz_7536 = ($signed(_zz_7537) >>> _zz_664);
  assign _zz_7537 = _zz_7538;
  assign _zz_7538 = ($signed(_zz_7540) - $signed(_zz_661));
  assign _zz_7539 = ({9'd0,data_mid_4_4_real} <<< 9);
  assign _zz_7540 = {{9{_zz_7539[26]}}, _zz_7539};
  assign _zz_7541 = fixTo_794_dout;
  assign _zz_7542 = _zz_7543[35 : 0];
  assign _zz_7543 = _zz_7544;
  assign _zz_7544 = ($signed(_zz_7545) >>> _zz_664);
  assign _zz_7545 = _zz_7546;
  assign _zz_7546 = ($signed(_zz_7548) - $signed(_zz_662));
  assign _zz_7547 = ({9'd0,data_mid_4_4_imag} <<< 9);
  assign _zz_7548 = {{9{_zz_7547[26]}}, _zz_7547};
  assign _zz_7549 = fixTo_795_dout;
  assign _zz_7550 = _zz_7551[35 : 0];
  assign _zz_7551 = _zz_7552;
  assign _zz_7552 = ($signed(_zz_7553) >>> _zz_665);
  assign _zz_7553 = _zz_7554;
  assign _zz_7554 = ($signed(_zz_7556) + $signed(_zz_661));
  assign _zz_7555 = ({9'd0,data_mid_4_4_real} <<< 9);
  assign _zz_7556 = {{9{_zz_7555[26]}}, _zz_7555};
  assign _zz_7557 = fixTo_796_dout;
  assign _zz_7558 = _zz_7559[35 : 0];
  assign _zz_7559 = _zz_7560;
  assign _zz_7560 = ($signed(_zz_7561) >>> _zz_665);
  assign _zz_7561 = _zz_7562;
  assign _zz_7562 = ($signed(_zz_7564) + $signed(_zz_662));
  assign _zz_7563 = ({9'd0,data_mid_4_4_imag} <<< 9);
  assign _zz_7564 = {{9{_zz_7563[26]}}, _zz_7563};
  assign _zz_7565 = fixTo_797_dout;
  assign _zz_7566 = ($signed(twiddle_factor_table_20_real) + $signed(twiddle_factor_table_20_imag));
  assign _zz_7567 = ($signed(_zz_668) - $signed(_zz_7568));
  assign _zz_7568 = ($signed(_zz_7569) * $signed(twiddle_factor_table_20_imag));
  assign _zz_7569 = ($signed(data_mid_4_21_real) + $signed(data_mid_4_21_imag));
  assign _zz_7570 = fixTo_798_dout;
  assign _zz_7571 = ($signed(_zz_668) + $signed(_zz_7572));
  assign _zz_7572 = ($signed(_zz_7573) * $signed(twiddle_factor_table_20_real));
  assign _zz_7573 = ($signed(data_mid_4_21_imag) - $signed(data_mid_4_21_real));
  assign _zz_7574 = fixTo_799_dout;
  assign _zz_7575 = _zz_7576[35 : 0];
  assign _zz_7576 = _zz_7577;
  assign _zz_7577 = ($signed(_zz_7578) >>> _zz_669);
  assign _zz_7578 = _zz_7579;
  assign _zz_7579 = ($signed(_zz_7581) - $signed(_zz_666));
  assign _zz_7580 = ({9'd0,data_mid_4_5_real} <<< 9);
  assign _zz_7581 = {{9{_zz_7580[26]}}, _zz_7580};
  assign _zz_7582 = fixTo_800_dout;
  assign _zz_7583 = _zz_7584[35 : 0];
  assign _zz_7584 = _zz_7585;
  assign _zz_7585 = ($signed(_zz_7586) >>> _zz_669);
  assign _zz_7586 = _zz_7587;
  assign _zz_7587 = ($signed(_zz_7589) - $signed(_zz_667));
  assign _zz_7588 = ({9'd0,data_mid_4_5_imag} <<< 9);
  assign _zz_7589 = {{9{_zz_7588[26]}}, _zz_7588};
  assign _zz_7590 = fixTo_801_dout;
  assign _zz_7591 = _zz_7592[35 : 0];
  assign _zz_7592 = _zz_7593;
  assign _zz_7593 = ($signed(_zz_7594) >>> _zz_670);
  assign _zz_7594 = _zz_7595;
  assign _zz_7595 = ($signed(_zz_7597) + $signed(_zz_666));
  assign _zz_7596 = ({9'd0,data_mid_4_5_real} <<< 9);
  assign _zz_7597 = {{9{_zz_7596[26]}}, _zz_7596};
  assign _zz_7598 = fixTo_802_dout;
  assign _zz_7599 = _zz_7600[35 : 0];
  assign _zz_7600 = _zz_7601;
  assign _zz_7601 = ($signed(_zz_7602) >>> _zz_670);
  assign _zz_7602 = _zz_7603;
  assign _zz_7603 = ($signed(_zz_7605) + $signed(_zz_667));
  assign _zz_7604 = ({9'd0,data_mid_4_5_imag} <<< 9);
  assign _zz_7605 = {{9{_zz_7604[26]}}, _zz_7604};
  assign _zz_7606 = fixTo_803_dout;
  assign _zz_7607 = ($signed(twiddle_factor_table_21_real) + $signed(twiddle_factor_table_21_imag));
  assign _zz_7608 = ($signed(_zz_673) - $signed(_zz_7609));
  assign _zz_7609 = ($signed(_zz_7610) * $signed(twiddle_factor_table_21_imag));
  assign _zz_7610 = ($signed(data_mid_4_22_real) + $signed(data_mid_4_22_imag));
  assign _zz_7611 = fixTo_804_dout;
  assign _zz_7612 = ($signed(_zz_673) + $signed(_zz_7613));
  assign _zz_7613 = ($signed(_zz_7614) * $signed(twiddle_factor_table_21_real));
  assign _zz_7614 = ($signed(data_mid_4_22_imag) - $signed(data_mid_4_22_real));
  assign _zz_7615 = fixTo_805_dout;
  assign _zz_7616 = _zz_7617[35 : 0];
  assign _zz_7617 = _zz_7618;
  assign _zz_7618 = ($signed(_zz_7619) >>> _zz_674);
  assign _zz_7619 = _zz_7620;
  assign _zz_7620 = ($signed(_zz_7622) - $signed(_zz_671));
  assign _zz_7621 = ({9'd0,data_mid_4_6_real} <<< 9);
  assign _zz_7622 = {{9{_zz_7621[26]}}, _zz_7621};
  assign _zz_7623 = fixTo_806_dout;
  assign _zz_7624 = _zz_7625[35 : 0];
  assign _zz_7625 = _zz_7626;
  assign _zz_7626 = ($signed(_zz_7627) >>> _zz_674);
  assign _zz_7627 = _zz_7628;
  assign _zz_7628 = ($signed(_zz_7630) - $signed(_zz_672));
  assign _zz_7629 = ({9'd0,data_mid_4_6_imag} <<< 9);
  assign _zz_7630 = {{9{_zz_7629[26]}}, _zz_7629};
  assign _zz_7631 = fixTo_807_dout;
  assign _zz_7632 = _zz_7633[35 : 0];
  assign _zz_7633 = _zz_7634;
  assign _zz_7634 = ($signed(_zz_7635) >>> _zz_675);
  assign _zz_7635 = _zz_7636;
  assign _zz_7636 = ($signed(_zz_7638) + $signed(_zz_671));
  assign _zz_7637 = ({9'd0,data_mid_4_6_real} <<< 9);
  assign _zz_7638 = {{9{_zz_7637[26]}}, _zz_7637};
  assign _zz_7639 = fixTo_808_dout;
  assign _zz_7640 = _zz_7641[35 : 0];
  assign _zz_7641 = _zz_7642;
  assign _zz_7642 = ($signed(_zz_7643) >>> _zz_675);
  assign _zz_7643 = _zz_7644;
  assign _zz_7644 = ($signed(_zz_7646) + $signed(_zz_672));
  assign _zz_7645 = ({9'd0,data_mid_4_6_imag} <<< 9);
  assign _zz_7646 = {{9{_zz_7645[26]}}, _zz_7645};
  assign _zz_7647 = fixTo_809_dout;
  assign _zz_7648 = ($signed(twiddle_factor_table_22_real) + $signed(twiddle_factor_table_22_imag));
  assign _zz_7649 = ($signed(_zz_678) - $signed(_zz_7650));
  assign _zz_7650 = ($signed(_zz_7651) * $signed(twiddle_factor_table_22_imag));
  assign _zz_7651 = ($signed(data_mid_4_23_real) + $signed(data_mid_4_23_imag));
  assign _zz_7652 = fixTo_810_dout;
  assign _zz_7653 = ($signed(_zz_678) + $signed(_zz_7654));
  assign _zz_7654 = ($signed(_zz_7655) * $signed(twiddle_factor_table_22_real));
  assign _zz_7655 = ($signed(data_mid_4_23_imag) - $signed(data_mid_4_23_real));
  assign _zz_7656 = fixTo_811_dout;
  assign _zz_7657 = _zz_7658[35 : 0];
  assign _zz_7658 = _zz_7659;
  assign _zz_7659 = ($signed(_zz_7660) >>> _zz_679);
  assign _zz_7660 = _zz_7661;
  assign _zz_7661 = ($signed(_zz_7663) - $signed(_zz_676));
  assign _zz_7662 = ({9'd0,data_mid_4_7_real} <<< 9);
  assign _zz_7663 = {{9{_zz_7662[26]}}, _zz_7662};
  assign _zz_7664 = fixTo_812_dout;
  assign _zz_7665 = _zz_7666[35 : 0];
  assign _zz_7666 = _zz_7667;
  assign _zz_7667 = ($signed(_zz_7668) >>> _zz_679);
  assign _zz_7668 = _zz_7669;
  assign _zz_7669 = ($signed(_zz_7671) - $signed(_zz_677));
  assign _zz_7670 = ({9'd0,data_mid_4_7_imag} <<< 9);
  assign _zz_7671 = {{9{_zz_7670[26]}}, _zz_7670};
  assign _zz_7672 = fixTo_813_dout;
  assign _zz_7673 = _zz_7674[35 : 0];
  assign _zz_7674 = _zz_7675;
  assign _zz_7675 = ($signed(_zz_7676) >>> _zz_680);
  assign _zz_7676 = _zz_7677;
  assign _zz_7677 = ($signed(_zz_7679) + $signed(_zz_676));
  assign _zz_7678 = ({9'd0,data_mid_4_7_real} <<< 9);
  assign _zz_7679 = {{9{_zz_7678[26]}}, _zz_7678};
  assign _zz_7680 = fixTo_814_dout;
  assign _zz_7681 = _zz_7682[35 : 0];
  assign _zz_7682 = _zz_7683;
  assign _zz_7683 = ($signed(_zz_7684) >>> _zz_680);
  assign _zz_7684 = _zz_7685;
  assign _zz_7685 = ($signed(_zz_7687) + $signed(_zz_677));
  assign _zz_7686 = ({9'd0,data_mid_4_7_imag} <<< 9);
  assign _zz_7687 = {{9{_zz_7686[26]}}, _zz_7686};
  assign _zz_7688 = fixTo_815_dout;
  assign _zz_7689 = ($signed(twiddle_factor_table_23_real) + $signed(twiddle_factor_table_23_imag));
  assign _zz_7690 = ($signed(_zz_683) - $signed(_zz_7691));
  assign _zz_7691 = ($signed(_zz_7692) * $signed(twiddle_factor_table_23_imag));
  assign _zz_7692 = ($signed(data_mid_4_24_real) + $signed(data_mid_4_24_imag));
  assign _zz_7693 = fixTo_816_dout;
  assign _zz_7694 = ($signed(_zz_683) + $signed(_zz_7695));
  assign _zz_7695 = ($signed(_zz_7696) * $signed(twiddle_factor_table_23_real));
  assign _zz_7696 = ($signed(data_mid_4_24_imag) - $signed(data_mid_4_24_real));
  assign _zz_7697 = fixTo_817_dout;
  assign _zz_7698 = _zz_7699[35 : 0];
  assign _zz_7699 = _zz_7700;
  assign _zz_7700 = ($signed(_zz_7701) >>> _zz_684);
  assign _zz_7701 = _zz_7702;
  assign _zz_7702 = ($signed(_zz_7704) - $signed(_zz_681));
  assign _zz_7703 = ({9'd0,data_mid_4_8_real} <<< 9);
  assign _zz_7704 = {{9{_zz_7703[26]}}, _zz_7703};
  assign _zz_7705 = fixTo_818_dout;
  assign _zz_7706 = _zz_7707[35 : 0];
  assign _zz_7707 = _zz_7708;
  assign _zz_7708 = ($signed(_zz_7709) >>> _zz_684);
  assign _zz_7709 = _zz_7710;
  assign _zz_7710 = ($signed(_zz_7712) - $signed(_zz_682));
  assign _zz_7711 = ({9'd0,data_mid_4_8_imag} <<< 9);
  assign _zz_7712 = {{9{_zz_7711[26]}}, _zz_7711};
  assign _zz_7713 = fixTo_819_dout;
  assign _zz_7714 = _zz_7715[35 : 0];
  assign _zz_7715 = _zz_7716;
  assign _zz_7716 = ($signed(_zz_7717) >>> _zz_685);
  assign _zz_7717 = _zz_7718;
  assign _zz_7718 = ($signed(_zz_7720) + $signed(_zz_681));
  assign _zz_7719 = ({9'd0,data_mid_4_8_real} <<< 9);
  assign _zz_7720 = {{9{_zz_7719[26]}}, _zz_7719};
  assign _zz_7721 = fixTo_820_dout;
  assign _zz_7722 = _zz_7723[35 : 0];
  assign _zz_7723 = _zz_7724;
  assign _zz_7724 = ($signed(_zz_7725) >>> _zz_685);
  assign _zz_7725 = _zz_7726;
  assign _zz_7726 = ($signed(_zz_7728) + $signed(_zz_682));
  assign _zz_7727 = ({9'd0,data_mid_4_8_imag} <<< 9);
  assign _zz_7728 = {{9{_zz_7727[26]}}, _zz_7727};
  assign _zz_7729 = fixTo_821_dout;
  assign _zz_7730 = ($signed(twiddle_factor_table_24_real) + $signed(twiddle_factor_table_24_imag));
  assign _zz_7731 = ($signed(_zz_688) - $signed(_zz_7732));
  assign _zz_7732 = ($signed(_zz_7733) * $signed(twiddle_factor_table_24_imag));
  assign _zz_7733 = ($signed(data_mid_4_25_real) + $signed(data_mid_4_25_imag));
  assign _zz_7734 = fixTo_822_dout;
  assign _zz_7735 = ($signed(_zz_688) + $signed(_zz_7736));
  assign _zz_7736 = ($signed(_zz_7737) * $signed(twiddle_factor_table_24_real));
  assign _zz_7737 = ($signed(data_mid_4_25_imag) - $signed(data_mid_4_25_real));
  assign _zz_7738 = fixTo_823_dout;
  assign _zz_7739 = _zz_7740[35 : 0];
  assign _zz_7740 = _zz_7741;
  assign _zz_7741 = ($signed(_zz_7742) >>> _zz_689);
  assign _zz_7742 = _zz_7743;
  assign _zz_7743 = ($signed(_zz_7745) - $signed(_zz_686));
  assign _zz_7744 = ({9'd0,data_mid_4_9_real} <<< 9);
  assign _zz_7745 = {{9{_zz_7744[26]}}, _zz_7744};
  assign _zz_7746 = fixTo_824_dout;
  assign _zz_7747 = _zz_7748[35 : 0];
  assign _zz_7748 = _zz_7749;
  assign _zz_7749 = ($signed(_zz_7750) >>> _zz_689);
  assign _zz_7750 = _zz_7751;
  assign _zz_7751 = ($signed(_zz_7753) - $signed(_zz_687));
  assign _zz_7752 = ({9'd0,data_mid_4_9_imag} <<< 9);
  assign _zz_7753 = {{9{_zz_7752[26]}}, _zz_7752};
  assign _zz_7754 = fixTo_825_dout;
  assign _zz_7755 = _zz_7756[35 : 0];
  assign _zz_7756 = _zz_7757;
  assign _zz_7757 = ($signed(_zz_7758) >>> _zz_690);
  assign _zz_7758 = _zz_7759;
  assign _zz_7759 = ($signed(_zz_7761) + $signed(_zz_686));
  assign _zz_7760 = ({9'd0,data_mid_4_9_real} <<< 9);
  assign _zz_7761 = {{9{_zz_7760[26]}}, _zz_7760};
  assign _zz_7762 = fixTo_826_dout;
  assign _zz_7763 = _zz_7764[35 : 0];
  assign _zz_7764 = _zz_7765;
  assign _zz_7765 = ($signed(_zz_7766) >>> _zz_690);
  assign _zz_7766 = _zz_7767;
  assign _zz_7767 = ($signed(_zz_7769) + $signed(_zz_687));
  assign _zz_7768 = ({9'd0,data_mid_4_9_imag} <<< 9);
  assign _zz_7769 = {{9{_zz_7768[26]}}, _zz_7768};
  assign _zz_7770 = fixTo_827_dout;
  assign _zz_7771 = ($signed(twiddle_factor_table_25_real) + $signed(twiddle_factor_table_25_imag));
  assign _zz_7772 = ($signed(_zz_693) - $signed(_zz_7773));
  assign _zz_7773 = ($signed(_zz_7774) * $signed(twiddle_factor_table_25_imag));
  assign _zz_7774 = ($signed(data_mid_4_26_real) + $signed(data_mid_4_26_imag));
  assign _zz_7775 = fixTo_828_dout;
  assign _zz_7776 = ($signed(_zz_693) + $signed(_zz_7777));
  assign _zz_7777 = ($signed(_zz_7778) * $signed(twiddle_factor_table_25_real));
  assign _zz_7778 = ($signed(data_mid_4_26_imag) - $signed(data_mid_4_26_real));
  assign _zz_7779 = fixTo_829_dout;
  assign _zz_7780 = _zz_7781[35 : 0];
  assign _zz_7781 = _zz_7782;
  assign _zz_7782 = ($signed(_zz_7783) >>> _zz_694);
  assign _zz_7783 = _zz_7784;
  assign _zz_7784 = ($signed(_zz_7786) - $signed(_zz_691));
  assign _zz_7785 = ({9'd0,data_mid_4_10_real} <<< 9);
  assign _zz_7786 = {{9{_zz_7785[26]}}, _zz_7785};
  assign _zz_7787 = fixTo_830_dout;
  assign _zz_7788 = _zz_7789[35 : 0];
  assign _zz_7789 = _zz_7790;
  assign _zz_7790 = ($signed(_zz_7791) >>> _zz_694);
  assign _zz_7791 = _zz_7792;
  assign _zz_7792 = ($signed(_zz_7794) - $signed(_zz_692));
  assign _zz_7793 = ({9'd0,data_mid_4_10_imag} <<< 9);
  assign _zz_7794 = {{9{_zz_7793[26]}}, _zz_7793};
  assign _zz_7795 = fixTo_831_dout;
  assign _zz_7796 = _zz_7797[35 : 0];
  assign _zz_7797 = _zz_7798;
  assign _zz_7798 = ($signed(_zz_7799) >>> _zz_695);
  assign _zz_7799 = _zz_7800;
  assign _zz_7800 = ($signed(_zz_7802) + $signed(_zz_691));
  assign _zz_7801 = ({9'd0,data_mid_4_10_real} <<< 9);
  assign _zz_7802 = {{9{_zz_7801[26]}}, _zz_7801};
  assign _zz_7803 = fixTo_832_dout;
  assign _zz_7804 = _zz_7805[35 : 0];
  assign _zz_7805 = _zz_7806;
  assign _zz_7806 = ($signed(_zz_7807) >>> _zz_695);
  assign _zz_7807 = _zz_7808;
  assign _zz_7808 = ($signed(_zz_7810) + $signed(_zz_692));
  assign _zz_7809 = ({9'd0,data_mid_4_10_imag} <<< 9);
  assign _zz_7810 = {{9{_zz_7809[26]}}, _zz_7809};
  assign _zz_7811 = fixTo_833_dout;
  assign _zz_7812 = ($signed(twiddle_factor_table_26_real) + $signed(twiddle_factor_table_26_imag));
  assign _zz_7813 = ($signed(_zz_698) - $signed(_zz_7814));
  assign _zz_7814 = ($signed(_zz_7815) * $signed(twiddle_factor_table_26_imag));
  assign _zz_7815 = ($signed(data_mid_4_27_real) + $signed(data_mid_4_27_imag));
  assign _zz_7816 = fixTo_834_dout;
  assign _zz_7817 = ($signed(_zz_698) + $signed(_zz_7818));
  assign _zz_7818 = ($signed(_zz_7819) * $signed(twiddle_factor_table_26_real));
  assign _zz_7819 = ($signed(data_mid_4_27_imag) - $signed(data_mid_4_27_real));
  assign _zz_7820 = fixTo_835_dout;
  assign _zz_7821 = _zz_7822[35 : 0];
  assign _zz_7822 = _zz_7823;
  assign _zz_7823 = ($signed(_zz_7824) >>> _zz_699);
  assign _zz_7824 = _zz_7825;
  assign _zz_7825 = ($signed(_zz_7827) - $signed(_zz_696));
  assign _zz_7826 = ({9'd0,data_mid_4_11_real} <<< 9);
  assign _zz_7827 = {{9{_zz_7826[26]}}, _zz_7826};
  assign _zz_7828 = fixTo_836_dout;
  assign _zz_7829 = _zz_7830[35 : 0];
  assign _zz_7830 = _zz_7831;
  assign _zz_7831 = ($signed(_zz_7832) >>> _zz_699);
  assign _zz_7832 = _zz_7833;
  assign _zz_7833 = ($signed(_zz_7835) - $signed(_zz_697));
  assign _zz_7834 = ({9'd0,data_mid_4_11_imag} <<< 9);
  assign _zz_7835 = {{9{_zz_7834[26]}}, _zz_7834};
  assign _zz_7836 = fixTo_837_dout;
  assign _zz_7837 = _zz_7838[35 : 0];
  assign _zz_7838 = _zz_7839;
  assign _zz_7839 = ($signed(_zz_7840) >>> _zz_700);
  assign _zz_7840 = _zz_7841;
  assign _zz_7841 = ($signed(_zz_7843) + $signed(_zz_696));
  assign _zz_7842 = ({9'd0,data_mid_4_11_real} <<< 9);
  assign _zz_7843 = {{9{_zz_7842[26]}}, _zz_7842};
  assign _zz_7844 = fixTo_838_dout;
  assign _zz_7845 = _zz_7846[35 : 0];
  assign _zz_7846 = _zz_7847;
  assign _zz_7847 = ($signed(_zz_7848) >>> _zz_700);
  assign _zz_7848 = _zz_7849;
  assign _zz_7849 = ($signed(_zz_7851) + $signed(_zz_697));
  assign _zz_7850 = ({9'd0,data_mid_4_11_imag} <<< 9);
  assign _zz_7851 = {{9{_zz_7850[26]}}, _zz_7850};
  assign _zz_7852 = fixTo_839_dout;
  assign _zz_7853 = ($signed(twiddle_factor_table_27_real) + $signed(twiddle_factor_table_27_imag));
  assign _zz_7854 = ($signed(_zz_703) - $signed(_zz_7855));
  assign _zz_7855 = ($signed(_zz_7856) * $signed(twiddle_factor_table_27_imag));
  assign _zz_7856 = ($signed(data_mid_4_28_real) + $signed(data_mid_4_28_imag));
  assign _zz_7857 = fixTo_840_dout;
  assign _zz_7858 = ($signed(_zz_703) + $signed(_zz_7859));
  assign _zz_7859 = ($signed(_zz_7860) * $signed(twiddle_factor_table_27_real));
  assign _zz_7860 = ($signed(data_mid_4_28_imag) - $signed(data_mid_4_28_real));
  assign _zz_7861 = fixTo_841_dout;
  assign _zz_7862 = _zz_7863[35 : 0];
  assign _zz_7863 = _zz_7864;
  assign _zz_7864 = ($signed(_zz_7865) >>> _zz_704);
  assign _zz_7865 = _zz_7866;
  assign _zz_7866 = ($signed(_zz_7868) - $signed(_zz_701));
  assign _zz_7867 = ({9'd0,data_mid_4_12_real} <<< 9);
  assign _zz_7868 = {{9{_zz_7867[26]}}, _zz_7867};
  assign _zz_7869 = fixTo_842_dout;
  assign _zz_7870 = _zz_7871[35 : 0];
  assign _zz_7871 = _zz_7872;
  assign _zz_7872 = ($signed(_zz_7873) >>> _zz_704);
  assign _zz_7873 = _zz_7874;
  assign _zz_7874 = ($signed(_zz_7876) - $signed(_zz_702));
  assign _zz_7875 = ({9'd0,data_mid_4_12_imag} <<< 9);
  assign _zz_7876 = {{9{_zz_7875[26]}}, _zz_7875};
  assign _zz_7877 = fixTo_843_dout;
  assign _zz_7878 = _zz_7879[35 : 0];
  assign _zz_7879 = _zz_7880;
  assign _zz_7880 = ($signed(_zz_7881) >>> _zz_705);
  assign _zz_7881 = _zz_7882;
  assign _zz_7882 = ($signed(_zz_7884) + $signed(_zz_701));
  assign _zz_7883 = ({9'd0,data_mid_4_12_real} <<< 9);
  assign _zz_7884 = {{9{_zz_7883[26]}}, _zz_7883};
  assign _zz_7885 = fixTo_844_dout;
  assign _zz_7886 = _zz_7887[35 : 0];
  assign _zz_7887 = _zz_7888;
  assign _zz_7888 = ($signed(_zz_7889) >>> _zz_705);
  assign _zz_7889 = _zz_7890;
  assign _zz_7890 = ($signed(_zz_7892) + $signed(_zz_702));
  assign _zz_7891 = ({9'd0,data_mid_4_12_imag} <<< 9);
  assign _zz_7892 = {{9{_zz_7891[26]}}, _zz_7891};
  assign _zz_7893 = fixTo_845_dout;
  assign _zz_7894 = ($signed(twiddle_factor_table_28_real) + $signed(twiddle_factor_table_28_imag));
  assign _zz_7895 = ($signed(_zz_708) - $signed(_zz_7896));
  assign _zz_7896 = ($signed(_zz_7897) * $signed(twiddle_factor_table_28_imag));
  assign _zz_7897 = ($signed(data_mid_4_29_real) + $signed(data_mid_4_29_imag));
  assign _zz_7898 = fixTo_846_dout;
  assign _zz_7899 = ($signed(_zz_708) + $signed(_zz_7900));
  assign _zz_7900 = ($signed(_zz_7901) * $signed(twiddle_factor_table_28_real));
  assign _zz_7901 = ($signed(data_mid_4_29_imag) - $signed(data_mid_4_29_real));
  assign _zz_7902 = fixTo_847_dout;
  assign _zz_7903 = _zz_7904[35 : 0];
  assign _zz_7904 = _zz_7905;
  assign _zz_7905 = ($signed(_zz_7906) >>> _zz_709);
  assign _zz_7906 = _zz_7907;
  assign _zz_7907 = ($signed(_zz_7909) - $signed(_zz_706));
  assign _zz_7908 = ({9'd0,data_mid_4_13_real} <<< 9);
  assign _zz_7909 = {{9{_zz_7908[26]}}, _zz_7908};
  assign _zz_7910 = fixTo_848_dout;
  assign _zz_7911 = _zz_7912[35 : 0];
  assign _zz_7912 = _zz_7913;
  assign _zz_7913 = ($signed(_zz_7914) >>> _zz_709);
  assign _zz_7914 = _zz_7915;
  assign _zz_7915 = ($signed(_zz_7917) - $signed(_zz_707));
  assign _zz_7916 = ({9'd0,data_mid_4_13_imag} <<< 9);
  assign _zz_7917 = {{9{_zz_7916[26]}}, _zz_7916};
  assign _zz_7918 = fixTo_849_dout;
  assign _zz_7919 = _zz_7920[35 : 0];
  assign _zz_7920 = _zz_7921;
  assign _zz_7921 = ($signed(_zz_7922) >>> _zz_710);
  assign _zz_7922 = _zz_7923;
  assign _zz_7923 = ($signed(_zz_7925) + $signed(_zz_706));
  assign _zz_7924 = ({9'd0,data_mid_4_13_real} <<< 9);
  assign _zz_7925 = {{9{_zz_7924[26]}}, _zz_7924};
  assign _zz_7926 = fixTo_850_dout;
  assign _zz_7927 = _zz_7928[35 : 0];
  assign _zz_7928 = _zz_7929;
  assign _zz_7929 = ($signed(_zz_7930) >>> _zz_710);
  assign _zz_7930 = _zz_7931;
  assign _zz_7931 = ($signed(_zz_7933) + $signed(_zz_707));
  assign _zz_7932 = ({9'd0,data_mid_4_13_imag} <<< 9);
  assign _zz_7933 = {{9{_zz_7932[26]}}, _zz_7932};
  assign _zz_7934 = fixTo_851_dout;
  assign _zz_7935 = ($signed(twiddle_factor_table_29_real) + $signed(twiddle_factor_table_29_imag));
  assign _zz_7936 = ($signed(_zz_713) - $signed(_zz_7937));
  assign _zz_7937 = ($signed(_zz_7938) * $signed(twiddle_factor_table_29_imag));
  assign _zz_7938 = ($signed(data_mid_4_30_real) + $signed(data_mid_4_30_imag));
  assign _zz_7939 = fixTo_852_dout;
  assign _zz_7940 = ($signed(_zz_713) + $signed(_zz_7941));
  assign _zz_7941 = ($signed(_zz_7942) * $signed(twiddle_factor_table_29_real));
  assign _zz_7942 = ($signed(data_mid_4_30_imag) - $signed(data_mid_4_30_real));
  assign _zz_7943 = fixTo_853_dout;
  assign _zz_7944 = _zz_7945[35 : 0];
  assign _zz_7945 = _zz_7946;
  assign _zz_7946 = ($signed(_zz_7947) >>> _zz_714);
  assign _zz_7947 = _zz_7948;
  assign _zz_7948 = ($signed(_zz_7950) - $signed(_zz_711));
  assign _zz_7949 = ({9'd0,data_mid_4_14_real} <<< 9);
  assign _zz_7950 = {{9{_zz_7949[26]}}, _zz_7949};
  assign _zz_7951 = fixTo_854_dout;
  assign _zz_7952 = _zz_7953[35 : 0];
  assign _zz_7953 = _zz_7954;
  assign _zz_7954 = ($signed(_zz_7955) >>> _zz_714);
  assign _zz_7955 = _zz_7956;
  assign _zz_7956 = ($signed(_zz_7958) - $signed(_zz_712));
  assign _zz_7957 = ({9'd0,data_mid_4_14_imag} <<< 9);
  assign _zz_7958 = {{9{_zz_7957[26]}}, _zz_7957};
  assign _zz_7959 = fixTo_855_dout;
  assign _zz_7960 = _zz_7961[35 : 0];
  assign _zz_7961 = _zz_7962;
  assign _zz_7962 = ($signed(_zz_7963) >>> _zz_715);
  assign _zz_7963 = _zz_7964;
  assign _zz_7964 = ($signed(_zz_7966) + $signed(_zz_711));
  assign _zz_7965 = ({9'd0,data_mid_4_14_real} <<< 9);
  assign _zz_7966 = {{9{_zz_7965[26]}}, _zz_7965};
  assign _zz_7967 = fixTo_856_dout;
  assign _zz_7968 = _zz_7969[35 : 0];
  assign _zz_7969 = _zz_7970;
  assign _zz_7970 = ($signed(_zz_7971) >>> _zz_715);
  assign _zz_7971 = _zz_7972;
  assign _zz_7972 = ($signed(_zz_7974) + $signed(_zz_712));
  assign _zz_7973 = ({9'd0,data_mid_4_14_imag} <<< 9);
  assign _zz_7974 = {{9{_zz_7973[26]}}, _zz_7973};
  assign _zz_7975 = fixTo_857_dout;
  assign _zz_7976 = ($signed(twiddle_factor_table_30_real) + $signed(twiddle_factor_table_30_imag));
  assign _zz_7977 = ($signed(_zz_718) - $signed(_zz_7978));
  assign _zz_7978 = ($signed(_zz_7979) * $signed(twiddle_factor_table_30_imag));
  assign _zz_7979 = ($signed(data_mid_4_31_real) + $signed(data_mid_4_31_imag));
  assign _zz_7980 = fixTo_858_dout;
  assign _zz_7981 = ($signed(_zz_718) + $signed(_zz_7982));
  assign _zz_7982 = ($signed(_zz_7983) * $signed(twiddle_factor_table_30_real));
  assign _zz_7983 = ($signed(data_mid_4_31_imag) - $signed(data_mid_4_31_real));
  assign _zz_7984 = fixTo_859_dout;
  assign _zz_7985 = _zz_7986[35 : 0];
  assign _zz_7986 = _zz_7987;
  assign _zz_7987 = ($signed(_zz_7988) >>> _zz_719);
  assign _zz_7988 = _zz_7989;
  assign _zz_7989 = ($signed(_zz_7991) - $signed(_zz_716));
  assign _zz_7990 = ({9'd0,data_mid_4_15_real} <<< 9);
  assign _zz_7991 = {{9{_zz_7990[26]}}, _zz_7990};
  assign _zz_7992 = fixTo_860_dout;
  assign _zz_7993 = _zz_7994[35 : 0];
  assign _zz_7994 = _zz_7995;
  assign _zz_7995 = ($signed(_zz_7996) >>> _zz_719);
  assign _zz_7996 = _zz_7997;
  assign _zz_7997 = ($signed(_zz_7999) - $signed(_zz_717));
  assign _zz_7998 = ({9'd0,data_mid_4_15_imag} <<< 9);
  assign _zz_7999 = {{9{_zz_7998[26]}}, _zz_7998};
  assign _zz_8000 = fixTo_861_dout;
  assign _zz_8001 = _zz_8002[35 : 0];
  assign _zz_8002 = _zz_8003;
  assign _zz_8003 = ($signed(_zz_8004) >>> _zz_720);
  assign _zz_8004 = _zz_8005;
  assign _zz_8005 = ($signed(_zz_8007) + $signed(_zz_716));
  assign _zz_8006 = ({9'd0,data_mid_4_15_real} <<< 9);
  assign _zz_8007 = {{9{_zz_8006[26]}}, _zz_8006};
  assign _zz_8008 = fixTo_862_dout;
  assign _zz_8009 = _zz_8010[35 : 0];
  assign _zz_8010 = _zz_8011;
  assign _zz_8011 = ($signed(_zz_8012) >>> _zz_720);
  assign _zz_8012 = _zz_8013;
  assign _zz_8013 = ($signed(_zz_8015) + $signed(_zz_717));
  assign _zz_8014 = ({9'd0,data_mid_4_15_imag} <<< 9);
  assign _zz_8015 = {{9{_zz_8014[26]}}, _zz_8014};
  assign _zz_8016 = fixTo_863_dout;
  assign _zz_8017 = ($signed(twiddle_factor_table_15_real) + $signed(twiddle_factor_table_15_imag));
  assign _zz_8018 = ($signed(_zz_723) - $signed(_zz_8019));
  assign _zz_8019 = ($signed(_zz_8020) * $signed(twiddle_factor_table_15_imag));
  assign _zz_8020 = ($signed(data_mid_4_48_real) + $signed(data_mid_4_48_imag));
  assign _zz_8021 = fixTo_864_dout;
  assign _zz_8022 = ($signed(_zz_723) + $signed(_zz_8023));
  assign _zz_8023 = ($signed(_zz_8024) * $signed(twiddle_factor_table_15_real));
  assign _zz_8024 = ($signed(data_mid_4_48_imag) - $signed(data_mid_4_48_real));
  assign _zz_8025 = fixTo_865_dout;
  assign _zz_8026 = _zz_8027[35 : 0];
  assign _zz_8027 = _zz_8028;
  assign _zz_8028 = ($signed(_zz_8029) >>> _zz_724);
  assign _zz_8029 = _zz_8030;
  assign _zz_8030 = ($signed(_zz_8032) - $signed(_zz_721));
  assign _zz_8031 = ({9'd0,data_mid_4_32_real} <<< 9);
  assign _zz_8032 = {{9{_zz_8031[26]}}, _zz_8031};
  assign _zz_8033 = fixTo_866_dout;
  assign _zz_8034 = _zz_8035[35 : 0];
  assign _zz_8035 = _zz_8036;
  assign _zz_8036 = ($signed(_zz_8037) >>> _zz_724);
  assign _zz_8037 = _zz_8038;
  assign _zz_8038 = ($signed(_zz_8040) - $signed(_zz_722));
  assign _zz_8039 = ({9'd0,data_mid_4_32_imag} <<< 9);
  assign _zz_8040 = {{9{_zz_8039[26]}}, _zz_8039};
  assign _zz_8041 = fixTo_867_dout;
  assign _zz_8042 = _zz_8043[35 : 0];
  assign _zz_8043 = _zz_8044;
  assign _zz_8044 = ($signed(_zz_8045) >>> _zz_725);
  assign _zz_8045 = _zz_8046;
  assign _zz_8046 = ($signed(_zz_8048) + $signed(_zz_721));
  assign _zz_8047 = ({9'd0,data_mid_4_32_real} <<< 9);
  assign _zz_8048 = {{9{_zz_8047[26]}}, _zz_8047};
  assign _zz_8049 = fixTo_868_dout;
  assign _zz_8050 = _zz_8051[35 : 0];
  assign _zz_8051 = _zz_8052;
  assign _zz_8052 = ($signed(_zz_8053) >>> _zz_725);
  assign _zz_8053 = _zz_8054;
  assign _zz_8054 = ($signed(_zz_8056) + $signed(_zz_722));
  assign _zz_8055 = ({9'd0,data_mid_4_32_imag} <<< 9);
  assign _zz_8056 = {{9{_zz_8055[26]}}, _zz_8055};
  assign _zz_8057 = fixTo_869_dout;
  assign _zz_8058 = ($signed(twiddle_factor_table_16_real) + $signed(twiddle_factor_table_16_imag));
  assign _zz_8059 = ($signed(_zz_728) - $signed(_zz_8060));
  assign _zz_8060 = ($signed(_zz_8061) * $signed(twiddle_factor_table_16_imag));
  assign _zz_8061 = ($signed(data_mid_4_49_real) + $signed(data_mid_4_49_imag));
  assign _zz_8062 = fixTo_870_dout;
  assign _zz_8063 = ($signed(_zz_728) + $signed(_zz_8064));
  assign _zz_8064 = ($signed(_zz_8065) * $signed(twiddle_factor_table_16_real));
  assign _zz_8065 = ($signed(data_mid_4_49_imag) - $signed(data_mid_4_49_real));
  assign _zz_8066 = fixTo_871_dout;
  assign _zz_8067 = _zz_8068[35 : 0];
  assign _zz_8068 = _zz_8069;
  assign _zz_8069 = ($signed(_zz_8070) >>> _zz_729);
  assign _zz_8070 = _zz_8071;
  assign _zz_8071 = ($signed(_zz_8073) - $signed(_zz_726));
  assign _zz_8072 = ({9'd0,data_mid_4_33_real} <<< 9);
  assign _zz_8073 = {{9{_zz_8072[26]}}, _zz_8072};
  assign _zz_8074 = fixTo_872_dout;
  assign _zz_8075 = _zz_8076[35 : 0];
  assign _zz_8076 = _zz_8077;
  assign _zz_8077 = ($signed(_zz_8078) >>> _zz_729);
  assign _zz_8078 = _zz_8079;
  assign _zz_8079 = ($signed(_zz_8081) - $signed(_zz_727));
  assign _zz_8080 = ({9'd0,data_mid_4_33_imag} <<< 9);
  assign _zz_8081 = {{9{_zz_8080[26]}}, _zz_8080};
  assign _zz_8082 = fixTo_873_dout;
  assign _zz_8083 = _zz_8084[35 : 0];
  assign _zz_8084 = _zz_8085;
  assign _zz_8085 = ($signed(_zz_8086) >>> _zz_730);
  assign _zz_8086 = _zz_8087;
  assign _zz_8087 = ($signed(_zz_8089) + $signed(_zz_726));
  assign _zz_8088 = ({9'd0,data_mid_4_33_real} <<< 9);
  assign _zz_8089 = {{9{_zz_8088[26]}}, _zz_8088};
  assign _zz_8090 = fixTo_874_dout;
  assign _zz_8091 = _zz_8092[35 : 0];
  assign _zz_8092 = _zz_8093;
  assign _zz_8093 = ($signed(_zz_8094) >>> _zz_730);
  assign _zz_8094 = _zz_8095;
  assign _zz_8095 = ($signed(_zz_8097) + $signed(_zz_727));
  assign _zz_8096 = ({9'd0,data_mid_4_33_imag} <<< 9);
  assign _zz_8097 = {{9{_zz_8096[26]}}, _zz_8096};
  assign _zz_8098 = fixTo_875_dout;
  assign _zz_8099 = ($signed(twiddle_factor_table_17_real) + $signed(twiddle_factor_table_17_imag));
  assign _zz_8100 = ($signed(_zz_733) - $signed(_zz_8101));
  assign _zz_8101 = ($signed(_zz_8102) * $signed(twiddle_factor_table_17_imag));
  assign _zz_8102 = ($signed(data_mid_4_50_real) + $signed(data_mid_4_50_imag));
  assign _zz_8103 = fixTo_876_dout;
  assign _zz_8104 = ($signed(_zz_733) + $signed(_zz_8105));
  assign _zz_8105 = ($signed(_zz_8106) * $signed(twiddle_factor_table_17_real));
  assign _zz_8106 = ($signed(data_mid_4_50_imag) - $signed(data_mid_4_50_real));
  assign _zz_8107 = fixTo_877_dout;
  assign _zz_8108 = _zz_8109[35 : 0];
  assign _zz_8109 = _zz_8110;
  assign _zz_8110 = ($signed(_zz_8111) >>> _zz_734);
  assign _zz_8111 = _zz_8112;
  assign _zz_8112 = ($signed(_zz_8114) - $signed(_zz_731));
  assign _zz_8113 = ({9'd0,data_mid_4_34_real} <<< 9);
  assign _zz_8114 = {{9{_zz_8113[26]}}, _zz_8113};
  assign _zz_8115 = fixTo_878_dout;
  assign _zz_8116 = _zz_8117[35 : 0];
  assign _zz_8117 = _zz_8118;
  assign _zz_8118 = ($signed(_zz_8119) >>> _zz_734);
  assign _zz_8119 = _zz_8120;
  assign _zz_8120 = ($signed(_zz_8122) - $signed(_zz_732));
  assign _zz_8121 = ({9'd0,data_mid_4_34_imag} <<< 9);
  assign _zz_8122 = {{9{_zz_8121[26]}}, _zz_8121};
  assign _zz_8123 = fixTo_879_dout;
  assign _zz_8124 = _zz_8125[35 : 0];
  assign _zz_8125 = _zz_8126;
  assign _zz_8126 = ($signed(_zz_8127) >>> _zz_735);
  assign _zz_8127 = _zz_8128;
  assign _zz_8128 = ($signed(_zz_8130) + $signed(_zz_731));
  assign _zz_8129 = ({9'd0,data_mid_4_34_real} <<< 9);
  assign _zz_8130 = {{9{_zz_8129[26]}}, _zz_8129};
  assign _zz_8131 = fixTo_880_dout;
  assign _zz_8132 = _zz_8133[35 : 0];
  assign _zz_8133 = _zz_8134;
  assign _zz_8134 = ($signed(_zz_8135) >>> _zz_735);
  assign _zz_8135 = _zz_8136;
  assign _zz_8136 = ($signed(_zz_8138) + $signed(_zz_732));
  assign _zz_8137 = ({9'd0,data_mid_4_34_imag} <<< 9);
  assign _zz_8138 = {{9{_zz_8137[26]}}, _zz_8137};
  assign _zz_8139 = fixTo_881_dout;
  assign _zz_8140 = ($signed(twiddle_factor_table_18_real) + $signed(twiddle_factor_table_18_imag));
  assign _zz_8141 = ($signed(_zz_738) - $signed(_zz_8142));
  assign _zz_8142 = ($signed(_zz_8143) * $signed(twiddle_factor_table_18_imag));
  assign _zz_8143 = ($signed(data_mid_4_51_real) + $signed(data_mid_4_51_imag));
  assign _zz_8144 = fixTo_882_dout;
  assign _zz_8145 = ($signed(_zz_738) + $signed(_zz_8146));
  assign _zz_8146 = ($signed(_zz_8147) * $signed(twiddle_factor_table_18_real));
  assign _zz_8147 = ($signed(data_mid_4_51_imag) - $signed(data_mid_4_51_real));
  assign _zz_8148 = fixTo_883_dout;
  assign _zz_8149 = _zz_8150[35 : 0];
  assign _zz_8150 = _zz_8151;
  assign _zz_8151 = ($signed(_zz_8152) >>> _zz_739);
  assign _zz_8152 = _zz_8153;
  assign _zz_8153 = ($signed(_zz_8155) - $signed(_zz_736));
  assign _zz_8154 = ({9'd0,data_mid_4_35_real} <<< 9);
  assign _zz_8155 = {{9{_zz_8154[26]}}, _zz_8154};
  assign _zz_8156 = fixTo_884_dout;
  assign _zz_8157 = _zz_8158[35 : 0];
  assign _zz_8158 = _zz_8159;
  assign _zz_8159 = ($signed(_zz_8160) >>> _zz_739);
  assign _zz_8160 = _zz_8161;
  assign _zz_8161 = ($signed(_zz_8163) - $signed(_zz_737));
  assign _zz_8162 = ({9'd0,data_mid_4_35_imag} <<< 9);
  assign _zz_8163 = {{9{_zz_8162[26]}}, _zz_8162};
  assign _zz_8164 = fixTo_885_dout;
  assign _zz_8165 = _zz_8166[35 : 0];
  assign _zz_8166 = _zz_8167;
  assign _zz_8167 = ($signed(_zz_8168) >>> _zz_740);
  assign _zz_8168 = _zz_8169;
  assign _zz_8169 = ($signed(_zz_8171) + $signed(_zz_736));
  assign _zz_8170 = ({9'd0,data_mid_4_35_real} <<< 9);
  assign _zz_8171 = {{9{_zz_8170[26]}}, _zz_8170};
  assign _zz_8172 = fixTo_886_dout;
  assign _zz_8173 = _zz_8174[35 : 0];
  assign _zz_8174 = _zz_8175;
  assign _zz_8175 = ($signed(_zz_8176) >>> _zz_740);
  assign _zz_8176 = _zz_8177;
  assign _zz_8177 = ($signed(_zz_8179) + $signed(_zz_737));
  assign _zz_8178 = ({9'd0,data_mid_4_35_imag} <<< 9);
  assign _zz_8179 = {{9{_zz_8178[26]}}, _zz_8178};
  assign _zz_8180 = fixTo_887_dout;
  assign _zz_8181 = ($signed(twiddle_factor_table_19_real) + $signed(twiddle_factor_table_19_imag));
  assign _zz_8182 = ($signed(_zz_743) - $signed(_zz_8183));
  assign _zz_8183 = ($signed(_zz_8184) * $signed(twiddle_factor_table_19_imag));
  assign _zz_8184 = ($signed(data_mid_4_52_real) + $signed(data_mid_4_52_imag));
  assign _zz_8185 = fixTo_888_dout;
  assign _zz_8186 = ($signed(_zz_743) + $signed(_zz_8187));
  assign _zz_8187 = ($signed(_zz_8188) * $signed(twiddle_factor_table_19_real));
  assign _zz_8188 = ($signed(data_mid_4_52_imag) - $signed(data_mid_4_52_real));
  assign _zz_8189 = fixTo_889_dout;
  assign _zz_8190 = _zz_8191[35 : 0];
  assign _zz_8191 = _zz_8192;
  assign _zz_8192 = ($signed(_zz_8193) >>> _zz_744);
  assign _zz_8193 = _zz_8194;
  assign _zz_8194 = ($signed(_zz_8196) - $signed(_zz_741));
  assign _zz_8195 = ({9'd0,data_mid_4_36_real} <<< 9);
  assign _zz_8196 = {{9{_zz_8195[26]}}, _zz_8195};
  assign _zz_8197 = fixTo_890_dout;
  assign _zz_8198 = _zz_8199[35 : 0];
  assign _zz_8199 = _zz_8200;
  assign _zz_8200 = ($signed(_zz_8201) >>> _zz_744);
  assign _zz_8201 = _zz_8202;
  assign _zz_8202 = ($signed(_zz_8204) - $signed(_zz_742));
  assign _zz_8203 = ({9'd0,data_mid_4_36_imag} <<< 9);
  assign _zz_8204 = {{9{_zz_8203[26]}}, _zz_8203};
  assign _zz_8205 = fixTo_891_dout;
  assign _zz_8206 = _zz_8207[35 : 0];
  assign _zz_8207 = _zz_8208;
  assign _zz_8208 = ($signed(_zz_8209) >>> _zz_745);
  assign _zz_8209 = _zz_8210;
  assign _zz_8210 = ($signed(_zz_8212) + $signed(_zz_741));
  assign _zz_8211 = ({9'd0,data_mid_4_36_real} <<< 9);
  assign _zz_8212 = {{9{_zz_8211[26]}}, _zz_8211};
  assign _zz_8213 = fixTo_892_dout;
  assign _zz_8214 = _zz_8215[35 : 0];
  assign _zz_8215 = _zz_8216;
  assign _zz_8216 = ($signed(_zz_8217) >>> _zz_745);
  assign _zz_8217 = _zz_8218;
  assign _zz_8218 = ($signed(_zz_8220) + $signed(_zz_742));
  assign _zz_8219 = ({9'd0,data_mid_4_36_imag} <<< 9);
  assign _zz_8220 = {{9{_zz_8219[26]}}, _zz_8219};
  assign _zz_8221 = fixTo_893_dout;
  assign _zz_8222 = ($signed(twiddle_factor_table_20_real) + $signed(twiddle_factor_table_20_imag));
  assign _zz_8223 = ($signed(_zz_748) - $signed(_zz_8224));
  assign _zz_8224 = ($signed(_zz_8225) * $signed(twiddle_factor_table_20_imag));
  assign _zz_8225 = ($signed(data_mid_4_53_real) + $signed(data_mid_4_53_imag));
  assign _zz_8226 = fixTo_894_dout;
  assign _zz_8227 = ($signed(_zz_748) + $signed(_zz_8228));
  assign _zz_8228 = ($signed(_zz_8229) * $signed(twiddle_factor_table_20_real));
  assign _zz_8229 = ($signed(data_mid_4_53_imag) - $signed(data_mid_4_53_real));
  assign _zz_8230 = fixTo_895_dout;
  assign _zz_8231 = _zz_8232[35 : 0];
  assign _zz_8232 = _zz_8233;
  assign _zz_8233 = ($signed(_zz_8234) >>> _zz_749);
  assign _zz_8234 = _zz_8235;
  assign _zz_8235 = ($signed(_zz_8237) - $signed(_zz_746));
  assign _zz_8236 = ({9'd0,data_mid_4_37_real} <<< 9);
  assign _zz_8237 = {{9{_zz_8236[26]}}, _zz_8236};
  assign _zz_8238 = fixTo_896_dout;
  assign _zz_8239 = _zz_8240[35 : 0];
  assign _zz_8240 = _zz_8241;
  assign _zz_8241 = ($signed(_zz_8242) >>> _zz_749);
  assign _zz_8242 = _zz_8243;
  assign _zz_8243 = ($signed(_zz_8245) - $signed(_zz_747));
  assign _zz_8244 = ({9'd0,data_mid_4_37_imag} <<< 9);
  assign _zz_8245 = {{9{_zz_8244[26]}}, _zz_8244};
  assign _zz_8246 = fixTo_897_dout;
  assign _zz_8247 = _zz_8248[35 : 0];
  assign _zz_8248 = _zz_8249;
  assign _zz_8249 = ($signed(_zz_8250) >>> _zz_750);
  assign _zz_8250 = _zz_8251;
  assign _zz_8251 = ($signed(_zz_8253) + $signed(_zz_746));
  assign _zz_8252 = ({9'd0,data_mid_4_37_real} <<< 9);
  assign _zz_8253 = {{9{_zz_8252[26]}}, _zz_8252};
  assign _zz_8254 = fixTo_898_dout;
  assign _zz_8255 = _zz_8256[35 : 0];
  assign _zz_8256 = _zz_8257;
  assign _zz_8257 = ($signed(_zz_8258) >>> _zz_750);
  assign _zz_8258 = _zz_8259;
  assign _zz_8259 = ($signed(_zz_8261) + $signed(_zz_747));
  assign _zz_8260 = ({9'd0,data_mid_4_37_imag} <<< 9);
  assign _zz_8261 = {{9{_zz_8260[26]}}, _zz_8260};
  assign _zz_8262 = fixTo_899_dout;
  assign _zz_8263 = ($signed(twiddle_factor_table_21_real) + $signed(twiddle_factor_table_21_imag));
  assign _zz_8264 = ($signed(_zz_753) - $signed(_zz_8265));
  assign _zz_8265 = ($signed(_zz_8266) * $signed(twiddle_factor_table_21_imag));
  assign _zz_8266 = ($signed(data_mid_4_54_real) + $signed(data_mid_4_54_imag));
  assign _zz_8267 = fixTo_900_dout;
  assign _zz_8268 = ($signed(_zz_753) + $signed(_zz_8269));
  assign _zz_8269 = ($signed(_zz_8270) * $signed(twiddle_factor_table_21_real));
  assign _zz_8270 = ($signed(data_mid_4_54_imag) - $signed(data_mid_4_54_real));
  assign _zz_8271 = fixTo_901_dout;
  assign _zz_8272 = _zz_8273[35 : 0];
  assign _zz_8273 = _zz_8274;
  assign _zz_8274 = ($signed(_zz_8275) >>> _zz_754);
  assign _zz_8275 = _zz_8276;
  assign _zz_8276 = ($signed(_zz_8278) - $signed(_zz_751));
  assign _zz_8277 = ({9'd0,data_mid_4_38_real} <<< 9);
  assign _zz_8278 = {{9{_zz_8277[26]}}, _zz_8277};
  assign _zz_8279 = fixTo_902_dout;
  assign _zz_8280 = _zz_8281[35 : 0];
  assign _zz_8281 = _zz_8282;
  assign _zz_8282 = ($signed(_zz_8283) >>> _zz_754);
  assign _zz_8283 = _zz_8284;
  assign _zz_8284 = ($signed(_zz_8286) - $signed(_zz_752));
  assign _zz_8285 = ({9'd0,data_mid_4_38_imag} <<< 9);
  assign _zz_8286 = {{9{_zz_8285[26]}}, _zz_8285};
  assign _zz_8287 = fixTo_903_dout;
  assign _zz_8288 = _zz_8289[35 : 0];
  assign _zz_8289 = _zz_8290;
  assign _zz_8290 = ($signed(_zz_8291) >>> _zz_755);
  assign _zz_8291 = _zz_8292;
  assign _zz_8292 = ($signed(_zz_8294) + $signed(_zz_751));
  assign _zz_8293 = ({9'd0,data_mid_4_38_real} <<< 9);
  assign _zz_8294 = {{9{_zz_8293[26]}}, _zz_8293};
  assign _zz_8295 = fixTo_904_dout;
  assign _zz_8296 = _zz_8297[35 : 0];
  assign _zz_8297 = _zz_8298;
  assign _zz_8298 = ($signed(_zz_8299) >>> _zz_755);
  assign _zz_8299 = _zz_8300;
  assign _zz_8300 = ($signed(_zz_8302) + $signed(_zz_752));
  assign _zz_8301 = ({9'd0,data_mid_4_38_imag} <<< 9);
  assign _zz_8302 = {{9{_zz_8301[26]}}, _zz_8301};
  assign _zz_8303 = fixTo_905_dout;
  assign _zz_8304 = ($signed(twiddle_factor_table_22_real) + $signed(twiddle_factor_table_22_imag));
  assign _zz_8305 = ($signed(_zz_758) - $signed(_zz_8306));
  assign _zz_8306 = ($signed(_zz_8307) * $signed(twiddle_factor_table_22_imag));
  assign _zz_8307 = ($signed(data_mid_4_55_real) + $signed(data_mid_4_55_imag));
  assign _zz_8308 = fixTo_906_dout;
  assign _zz_8309 = ($signed(_zz_758) + $signed(_zz_8310));
  assign _zz_8310 = ($signed(_zz_8311) * $signed(twiddle_factor_table_22_real));
  assign _zz_8311 = ($signed(data_mid_4_55_imag) - $signed(data_mid_4_55_real));
  assign _zz_8312 = fixTo_907_dout;
  assign _zz_8313 = _zz_8314[35 : 0];
  assign _zz_8314 = _zz_8315;
  assign _zz_8315 = ($signed(_zz_8316) >>> _zz_759);
  assign _zz_8316 = _zz_8317;
  assign _zz_8317 = ($signed(_zz_8319) - $signed(_zz_756));
  assign _zz_8318 = ({9'd0,data_mid_4_39_real} <<< 9);
  assign _zz_8319 = {{9{_zz_8318[26]}}, _zz_8318};
  assign _zz_8320 = fixTo_908_dout;
  assign _zz_8321 = _zz_8322[35 : 0];
  assign _zz_8322 = _zz_8323;
  assign _zz_8323 = ($signed(_zz_8324) >>> _zz_759);
  assign _zz_8324 = _zz_8325;
  assign _zz_8325 = ($signed(_zz_8327) - $signed(_zz_757));
  assign _zz_8326 = ({9'd0,data_mid_4_39_imag} <<< 9);
  assign _zz_8327 = {{9{_zz_8326[26]}}, _zz_8326};
  assign _zz_8328 = fixTo_909_dout;
  assign _zz_8329 = _zz_8330[35 : 0];
  assign _zz_8330 = _zz_8331;
  assign _zz_8331 = ($signed(_zz_8332) >>> _zz_760);
  assign _zz_8332 = _zz_8333;
  assign _zz_8333 = ($signed(_zz_8335) + $signed(_zz_756));
  assign _zz_8334 = ({9'd0,data_mid_4_39_real} <<< 9);
  assign _zz_8335 = {{9{_zz_8334[26]}}, _zz_8334};
  assign _zz_8336 = fixTo_910_dout;
  assign _zz_8337 = _zz_8338[35 : 0];
  assign _zz_8338 = _zz_8339;
  assign _zz_8339 = ($signed(_zz_8340) >>> _zz_760);
  assign _zz_8340 = _zz_8341;
  assign _zz_8341 = ($signed(_zz_8343) + $signed(_zz_757));
  assign _zz_8342 = ({9'd0,data_mid_4_39_imag} <<< 9);
  assign _zz_8343 = {{9{_zz_8342[26]}}, _zz_8342};
  assign _zz_8344 = fixTo_911_dout;
  assign _zz_8345 = ($signed(twiddle_factor_table_23_real) + $signed(twiddle_factor_table_23_imag));
  assign _zz_8346 = ($signed(_zz_763) - $signed(_zz_8347));
  assign _zz_8347 = ($signed(_zz_8348) * $signed(twiddle_factor_table_23_imag));
  assign _zz_8348 = ($signed(data_mid_4_56_real) + $signed(data_mid_4_56_imag));
  assign _zz_8349 = fixTo_912_dout;
  assign _zz_8350 = ($signed(_zz_763) + $signed(_zz_8351));
  assign _zz_8351 = ($signed(_zz_8352) * $signed(twiddle_factor_table_23_real));
  assign _zz_8352 = ($signed(data_mid_4_56_imag) - $signed(data_mid_4_56_real));
  assign _zz_8353 = fixTo_913_dout;
  assign _zz_8354 = _zz_8355[35 : 0];
  assign _zz_8355 = _zz_8356;
  assign _zz_8356 = ($signed(_zz_8357) >>> _zz_764);
  assign _zz_8357 = _zz_8358;
  assign _zz_8358 = ($signed(_zz_8360) - $signed(_zz_761));
  assign _zz_8359 = ({9'd0,data_mid_4_40_real} <<< 9);
  assign _zz_8360 = {{9{_zz_8359[26]}}, _zz_8359};
  assign _zz_8361 = fixTo_914_dout;
  assign _zz_8362 = _zz_8363[35 : 0];
  assign _zz_8363 = _zz_8364;
  assign _zz_8364 = ($signed(_zz_8365) >>> _zz_764);
  assign _zz_8365 = _zz_8366;
  assign _zz_8366 = ($signed(_zz_8368) - $signed(_zz_762));
  assign _zz_8367 = ({9'd0,data_mid_4_40_imag} <<< 9);
  assign _zz_8368 = {{9{_zz_8367[26]}}, _zz_8367};
  assign _zz_8369 = fixTo_915_dout;
  assign _zz_8370 = _zz_8371[35 : 0];
  assign _zz_8371 = _zz_8372;
  assign _zz_8372 = ($signed(_zz_8373) >>> _zz_765);
  assign _zz_8373 = _zz_8374;
  assign _zz_8374 = ($signed(_zz_8376) + $signed(_zz_761));
  assign _zz_8375 = ({9'd0,data_mid_4_40_real} <<< 9);
  assign _zz_8376 = {{9{_zz_8375[26]}}, _zz_8375};
  assign _zz_8377 = fixTo_916_dout;
  assign _zz_8378 = _zz_8379[35 : 0];
  assign _zz_8379 = _zz_8380;
  assign _zz_8380 = ($signed(_zz_8381) >>> _zz_765);
  assign _zz_8381 = _zz_8382;
  assign _zz_8382 = ($signed(_zz_8384) + $signed(_zz_762));
  assign _zz_8383 = ({9'd0,data_mid_4_40_imag} <<< 9);
  assign _zz_8384 = {{9{_zz_8383[26]}}, _zz_8383};
  assign _zz_8385 = fixTo_917_dout;
  assign _zz_8386 = ($signed(twiddle_factor_table_24_real) + $signed(twiddle_factor_table_24_imag));
  assign _zz_8387 = ($signed(_zz_768) - $signed(_zz_8388));
  assign _zz_8388 = ($signed(_zz_8389) * $signed(twiddle_factor_table_24_imag));
  assign _zz_8389 = ($signed(data_mid_4_57_real) + $signed(data_mid_4_57_imag));
  assign _zz_8390 = fixTo_918_dout;
  assign _zz_8391 = ($signed(_zz_768) + $signed(_zz_8392));
  assign _zz_8392 = ($signed(_zz_8393) * $signed(twiddle_factor_table_24_real));
  assign _zz_8393 = ($signed(data_mid_4_57_imag) - $signed(data_mid_4_57_real));
  assign _zz_8394 = fixTo_919_dout;
  assign _zz_8395 = _zz_8396[35 : 0];
  assign _zz_8396 = _zz_8397;
  assign _zz_8397 = ($signed(_zz_8398) >>> _zz_769);
  assign _zz_8398 = _zz_8399;
  assign _zz_8399 = ($signed(_zz_8401) - $signed(_zz_766));
  assign _zz_8400 = ({9'd0,data_mid_4_41_real} <<< 9);
  assign _zz_8401 = {{9{_zz_8400[26]}}, _zz_8400};
  assign _zz_8402 = fixTo_920_dout;
  assign _zz_8403 = _zz_8404[35 : 0];
  assign _zz_8404 = _zz_8405;
  assign _zz_8405 = ($signed(_zz_8406) >>> _zz_769);
  assign _zz_8406 = _zz_8407;
  assign _zz_8407 = ($signed(_zz_8409) - $signed(_zz_767));
  assign _zz_8408 = ({9'd0,data_mid_4_41_imag} <<< 9);
  assign _zz_8409 = {{9{_zz_8408[26]}}, _zz_8408};
  assign _zz_8410 = fixTo_921_dout;
  assign _zz_8411 = _zz_8412[35 : 0];
  assign _zz_8412 = _zz_8413;
  assign _zz_8413 = ($signed(_zz_8414) >>> _zz_770);
  assign _zz_8414 = _zz_8415;
  assign _zz_8415 = ($signed(_zz_8417) + $signed(_zz_766));
  assign _zz_8416 = ({9'd0,data_mid_4_41_real} <<< 9);
  assign _zz_8417 = {{9{_zz_8416[26]}}, _zz_8416};
  assign _zz_8418 = fixTo_922_dout;
  assign _zz_8419 = _zz_8420[35 : 0];
  assign _zz_8420 = _zz_8421;
  assign _zz_8421 = ($signed(_zz_8422) >>> _zz_770);
  assign _zz_8422 = _zz_8423;
  assign _zz_8423 = ($signed(_zz_8425) + $signed(_zz_767));
  assign _zz_8424 = ({9'd0,data_mid_4_41_imag} <<< 9);
  assign _zz_8425 = {{9{_zz_8424[26]}}, _zz_8424};
  assign _zz_8426 = fixTo_923_dout;
  assign _zz_8427 = ($signed(twiddle_factor_table_25_real) + $signed(twiddle_factor_table_25_imag));
  assign _zz_8428 = ($signed(_zz_773) - $signed(_zz_8429));
  assign _zz_8429 = ($signed(_zz_8430) * $signed(twiddle_factor_table_25_imag));
  assign _zz_8430 = ($signed(data_mid_4_58_real) + $signed(data_mid_4_58_imag));
  assign _zz_8431 = fixTo_924_dout;
  assign _zz_8432 = ($signed(_zz_773) + $signed(_zz_8433));
  assign _zz_8433 = ($signed(_zz_8434) * $signed(twiddle_factor_table_25_real));
  assign _zz_8434 = ($signed(data_mid_4_58_imag) - $signed(data_mid_4_58_real));
  assign _zz_8435 = fixTo_925_dout;
  assign _zz_8436 = _zz_8437[35 : 0];
  assign _zz_8437 = _zz_8438;
  assign _zz_8438 = ($signed(_zz_8439) >>> _zz_774);
  assign _zz_8439 = _zz_8440;
  assign _zz_8440 = ($signed(_zz_8442) - $signed(_zz_771));
  assign _zz_8441 = ({9'd0,data_mid_4_42_real} <<< 9);
  assign _zz_8442 = {{9{_zz_8441[26]}}, _zz_8441};
  assign _zz_8443 = fixTo_926_dout;
  assign _zz_8444 = _zz_8445[35 : 0];
  assign _zz_8445 = _zz_8446;
  assign _zz_8446 = ($signed(_zz_8447) >>> _zz_774);
  assign _zz_8447 = _zz_8448;
  assign _zz_8448 = ($signed(_zz_8450) - $signed(_zz_772));
  assign _zz_8449 = ({9'd0,data_mid_4_42_imag} <<< 9);
  assign _zz_8450 = {{9{_zz_8449[26]}}, _zz_8449};
  assign _zz_8451 = fixTo_927_dout;
  assign _zz_8452 = _zz_8453[35 : 0];
  assign _zz_8453 = _zz_8454;
  assign _zz_8454 = ($signed(_zz_8455) >>> _zz_775);
  assign _zz_8455 = _zz_8456;
  assign _zz_8456 = ($signed(_zz_8458) + $signed(_zz_771));
  assign _zz_8457 = ({9'd0,data_mid_4_42_real} <<< 9);
  assign _zz_8458 = {{9{_zz_8457[26]}}, _zz_8457};
  assign _zz_8459 = fixTo_928_dout;
  assign _zz_8460 = _zz_8461[35 : 0];
  assign _zz_8461 = _zz_8462;
  assign _zz_8462 = ($signed(_zz_8463) >>> _zz_775);
  assign _zz_8463 = _zz_8464;
  assign _zz_8464 = ($signed(_zz_8466) + $signed(_zz_772));
  assign _zz_8465 = ({9'd0,data_mid_4_42_imag} <<< 9);
  assign _zz_8466 = {{9{_zz_8465[26]}}, _zz_8465};
  assign _zz_8467 = fixTo_929_dout;
  assign _zz_8468 = ($signed(twiddle_factor_table_26_real) + $signed(twiddle_factor_table_26_imag));
  assign _zz_8469 = ($signed(_zz_778) - $signed(_zz_8470));
  assign _zz_8470 = ($signed(_zz_8471) * $signed(twiddle_factor_table_26_imag));
  assign _zz_8471 = ($signed(data_mid_4_59_real) + $signed(data_mid_4_59_imag));
  assign _zz_8472 = fixTo_930_dout;
  assign _zz_8473 = ($signed(_zz_778) + $signed(_zz_8474));
  assign _zz_8474 = ($signed(_zz_8475) * $signed(twiddle_factor_table_26_real));
  assign _zz_8475 = ($signed(data_mid_4_59_imag) - $signed(data_mid_4_59_real));
  assign _zz_8476 = fixTo_931_dout;
  assign _zz_8477 = _zz_8478[35 : 0];
  assign _zz_8478 = _zz_8479;
  assign _zz_8479 = ($signed(_zz_8480) >>> _zz_779);
  assign _zz_8480 = _zz_8481;
  assign _zz_8481 = ($signed(_zz_8483) - $signed(_zz_776));
  assign _zz_8482 = ({9'd0,data_mid_4_43_real} <<< 9);
  assign _zz_8483 = {{9{_zz_8482[26]}}, _zz_8482};
  assign _zz_8484 = fixTo_932_dout;
  assign _zz_8485 = _zz_8486[35 : 0];
  assign _zz_8486 = _zz_8487;
  assign _zz_8487 = ($signed(_zz_8488) >>> _zz_779);
  assign _zz_8488 = _zz_8489;
  assign _zz_8489 = ($signed(_zz_8491) - $signed(_zz_777));
  assign _zz_8490 = ({9'd0,data_mid_4_43_imag} <<< 9);
  assign _zz_8491 = {{9{_zz_8490[26]}}, _zz_8490};
  assign _zz_8492 = fixTo_933_dout;
  assign _zz_8493 = _zz_8494[35 : 0];
  assign _zz_8494 = _zz_8495;
  assign _zz_8495 = ($signed(_zz_8496) >>> _zz_780);
  assign _zz_8496 = _zz_8497;
  assign _zz_8497 = ($signed(_zz_8499) + $signed(_zz_776));
  assign _zz_8498 = ({9'd0,data_mid_4_43_real} <<< 9);
  assign _zz_8499 = {{9{_zz_8498[26]}}, _zz_8498};
  assign _zz_8500 = fixTo_934_dout;
  assign _zz_8501 = _zz_8502[35 : 0];
  assign _zz_8502 = _zz_8503;
  assign _zz_8503 = ($signed(_zz_8504) >>> _zz_780);
  assign _zz_8504 = _zz_8505;
  assign _zz_8505 = ($signed(_zz_8507) + $signed(_zz_777));
  assign _zz_8506 = ({9'd0,data_mid_4_43_imag} <<< 9);
  assign _zz_8507 = {{9{_zz_8506[26]}}, _zz_8506};
  assign _zz_8508 = fixTo_935_dout;
  assign _zz_8509 = ($signed(twiddle_factor_table_27_real) + $signed(twiddle_factor_table_27_imag));
  assign _zz_8510 = ($signed(_zz_783) - $signed(_zz_8511));
  assign _zz_8511 = ($signed(_zz_8512) * $signed(twiddle_factor_table_27_imag));
  assign _zz_8512 = ($signed(data_mid_4_60_real) + $signed(data_mid_4_60_imag));
  assign _zz_8513 = fixTo_936_dout;
  assign _zz_8514 = ($signed(_zz_783) + $signed(_zz_8515));
  assign _zz_8515 = ($signed(_zz_8516) * $signed(twiddle_factor_table_27_real));
  assign _zz_8516 = ($signed(data_mid_4_60_imag) - $signed(data_mid_4_60_real));
  assign _zz_8517 = fixTo_937_dout;
  assign _zz_8518 = _zz_8519[35 : 0];
  assign _zz_8519 = _zz_8520;
  assign _zz_8520 = ($signed(_zz_8521) >>> _zz_784);
  assign _zz_8521 = _zz_8522;
  assign _zz_8522 = ($signed(_zz_8524) - $signed(_zz_781));
  assign _zz_8523 = ({9'd0,data_mid_4_44_real} <<< 9);
  assign _zz_8524 = {{9{_zz_8523[26]}}, _zz_8523};
  assign _zz_8525 = fixTo_938_dout;
  assign _zz_8526 = _zz_8527[35 : 0];
  assign _zz_8527 = _zz_8528;
  assign _zz_8528 = ($signed(_zz_8529) >>> _zz_784);
  assign _zz_8529 = _zz_8530;
  assign _zz_8530 = ($signed(_zz_8532) - $signed(_zz_782));
  assign _zz_8531 = ({9'd0,data_mid_4_44_imag} <<< 9);
  assign _zz_8532 = {{9{_zz_8531[26]}}, _zz_8531};
  assign _zz_8533 = fixTo_939_dout;
  assign _zz_8534 = _zz_8535[35 : 0];
  assign _zz_8535 = _zz_8536;
  assign _zz_8536 = ($signed(_zz_8537) >>> _zz_785);
  assign _zz_8537 = _zz_8538;
  assign _zz_8538 = ($signed(_zz_8540) + $signed(_zz_781));
  assign _zz_8539 = ({9'd0,data_mid_4_44_real} <<< 9);
  assign _zz_8540 = {{9{_zz_8539[26]}}, _zz_8539};
  assign _zz_8541 = fixTo_940_dout;
  assign _zz_8542 = _zz_8543[35 : 0];
  assign _zz_8543 = _zz_8544;
  assign _zz_8544 = ($signed(_zz_8545) >>> _zz_785);
  assign _zz_8545 = _zz_8546;
  assign _zz_8546 = ($signed(_zz_8548) + $signed(_zz_782));
  assign _zz_8547 = ({9'd0,data_mid_4_44_imag} <<< 9);
  assign _zz_8548 = {{9{_zz_8547[26]}}, _zz_8547};
  assign _zz_8549 = fixTo_941_dout;
  assign _zz_8550 = ($signed(twiddle_factor_table_28_real) + $signed(twiddle_factor_table_28_imag));
  assign _zz_8551 = ($signed(_zz_788) - $signed(_zz_8552));
  assign _zz_8552 = ($signed(_zz_8553) * $signed(twiddle_factor_table_28_imag));
  assign _zz_8553 = ($signed(data_mid_4_61_real) + $signed(data_mid_4_61_imag));
  assign _zz_8554 = fixTo_942_dout;
  assign _zz_8555 = ($signed(_zz_788) + $signed(_zz_8556));
  assign _zz_8556 = ($signed(_zz_8557) * $signed(twiddle_factor_table_28_real));
  assign _zz_8557 = ($signed(data_mid_4_61_imag) - $signed(data_mid_4_61_real));
  assign _zz_8558 = fixTo_943_dout;
  assign _zz_8559 = _zz_8560[35 : 0];
  assign _zz_8560 = _zz_8561;
  assign _zz_8561 = ($signed(_zz_8562) >>> _zz_789);
  assign _zz_8562 = _zz_8563;
  assign _zz_8563 = ($signed(_zz_8565) - $signed(_zz_786));
  assign _zz_8564 = ({9'd0,data_mid_4_45_real} <<< 9);
  assign _zz_8565 = {{9{_zz_8564[26]}}, _zz_8564};
  assign _zz_8566 = fixTo_944_dout;
  assign _zz_8567 = _zz_8568[35 : 0];
  assign _zz_8568 = _zz_8569;
  assign _zz_8569 = ($signed(_zz_8570) >>> _zz_789);
  assign _zz_8570 = _zz_8571;
  assign _zz_8571 = ($signed(_zz_8573) - $signed(_zz_787));
  assign _zz_8572 = ({9'd0,data_mid_4_45_imag} <<< 9);
  assign _zz_8573 = {{9{_zz_8572[26]}}, _zz_8572};
  assign _zz_8574 = fixTo_945_dout;
  assign _zz_8575 = _zz_8576[35 : 0];
  assign _zz_8576 = _zz_8577;
  assign _zz_8577 = ($signed(_zz_8578) >>> _zz_790);
  assign _zz_8578 = _zz_8579;
  assign _zz_8579 = ($signed(_zz_8581) + $signed(_zz_786));
  assign _zz_8580 = ({9'd0,data_mid_4_45_real} <<< 9);
  assign _zz_8581 = {{9{_zz_8580[26]}}, _zz_8580};
  assign _zz_8582 = fixTo_946_dout;
  assign _zz_8583 = _zz_8584[35 : 0];
  assign _zz_8584 = _zz_8585;
  assign _zz_8585 = ($signed(_zz_8586) >>> _zz_790);
  assign _zz_8586 = _zz_8587;
  assign _zz_8587 = ($signed(_zz_8589) + $signed(_zz_787));
  assign _zz_8588 = ({9'd0,data_mid_4_45_imag} <<< 9);
  assign _zz_8589 = {{9{_zz_8588[26]}}, _zz_8588};
  assign _zz_8590 = fixTo_947_dout;
  assign _zz_8591 = ($signed(twiddle_factor_table_29_real) + $signed(twiddle_factor_table_29_imag));
  assign _zz_8592 = ($signed(_zz_793) - $signed(_zz_8593));
  assign _zz_8593 = ($signed(_zz_8594) * $signed(twiddle_factor_table_29_imag));
  assign _zz_8594 = ($signed(data_mid_4_62_real) + $signed(data_mid_4_62_imag));
  assign _zz_8595 = fixTo_948_dout;
  assign _zz_8596 = ($signed(_zz_793) + $signed(_zz_8597));
  assign _zz_8597 = ($signed(_zz_8598) * $signed(twiddle_factor_table_29_real));
  assign _zz_8598 = ($signed(data_mid_4_62_imag) - $signed(data_mid_4_62_real));
  assign _zz_8599 = fixTo_949_dout;
  assign _zz_8600 = _zz_8601[35 : 0];
  assign _zz_8601 = _zz_8602;
  assign _zz_8602 = ($signed(_zz_8603) >>> _zz_794);
  assign _zz_8603 = _zz_8604;
  assign _zz_8604 = ($signed(_zz_8606) - $signed(_zz_791));
  assign _zz_8605 = ({9'd0,data_mid_4_46_real} <<< 9);
  assign _zz_8606 = {{9{_zz_8605[26]}}, _zz_8605};
  assign _zz_8607 = fixTo_950_dout;
  assign _zz_8608 = _zz_8609[35 : 0];
  assign _zz_8609 = _zz_8610;
  assign _zz_8610 = ($signed(_zz_8611) >>> _zz_794);
  assign _zz_8611 = _zz_8612;
  assign _zz_8612 = ($signed(_zz_8614) - $signed(_zz_792));
  assign _zz_8613 = ({9'd0,data_mid_4_46_imag} <<< 9);
  assign _zz_8614 = {{9{_zz_8613[26]}}, _zz_8613};
  assign _zz_8615 = fixTo_951_dout;
  assign _zz_8616 = _zz_8617[35 : 0];
  assign _zz_8617 = _zz_8618;
  assign _zz_8618 = ($signed(_zz_8619) >>> _zz_795);
  assign _zz_8619 = _zz_8620;
  assign _zz_8620 = ($signed(_zz_8622) + $signed(_zz_791));
  assign _zz_8621 = ({9'd0,data_mid_4_46_real} <<< 9);
  assign _zz_8622 = {{9{_zz_8621[26]}}, _zz_8621};
  assign _zz_8623 = fixTo_952_dout;
  assign _zz_8624 = _zz_8625[35 : 0];
  assign _zz_8625 = _zz_8626;
  assign _zz_8626 = ($signed(_zz_8627) >>> _zz_795);
  assign _zz_8627 = _zz_8628;
  assign _zz_8628 = ($signed(_zz_8630) + $signed(_zz_792));
  assign _zz_8629 = ({9'd0,data_mid_4_46_imag} <<< 9);
  assign _zz_8630 = {{9{_zz_8629[26]}}, _zz_8629};
  assign _zz_8631 = fixTo_953_dout;
  assign _zz_8632 = ($signed(twiddle_factor_table_30_real) + $signed(twiddle_factor_table_30_imag));
  assign _zz_8633 = ($signed(_zz_798) - $signed(_zz_8634));
  assign _zz_8634 = ($signed(_zz_8635) * $signed(twiddle_factor_table_30_imag));
  assign _zz_8635 = ($signed(data_mid_4_63_real) + $signed(data_mid_4_63_imag));
  assign _zz_8636 = fixTo_954_dout;
  assign _zz_8637 = ($signed(_zz_798) + $signed(_zz_8638));
  assign _zz_8638 = ($signed(_zz_8639) * $signed(twiddle_factor_table_30_real));
  assign _zz_8639 = ($signed(data_mid_4_63_imag) - $signed(data_mid_4_63_real));
  assign _zz_8640 = fixTo_955_dout;
  assign _zz_8641 = _zz_8642[35 : 0];
  assign _zz_8642 = _zz_8643;
  assign _zz_8643 = ($signed(_zz_8644) >>> _zz_799);
  assign _zz_8644 = _zz_8645;
  assign _zz_8645 = ($signed(_zz_8647) - $signed(_zz_796));
  assign _zz_8646 = ({9'd0,data_mid_4_47_real} <<< 9);
  assign _zz_8647 = {{9{_zz_8646[26]}}, _zz_8646};
  assign _zz_8648 = fixTo_956_dout;
  assign _zz_8649 = _zz_8650[35 : 0];
  assign _zz_8650 = _zz_8651;
  assign _zz_8651 = ($signed(_zz_8652) >>> _zz_799);
  assign _zz_8652 = _zz_8653;
  assign _zz_8653 = ($signed(_zz_8655) - $signed(_zz_797));
  assign _zz_8654 = ({9'd0,data_mid_4_47_imag} <<< 9);
  assign _zz_8655 = {{9{_zz_8654[26]}}, _zz_8654};
  assign _zz_8656 = fixTo_957_dout;
  assign _zz_8657 = _zz_8658[35 : 0];
  assign _zz_8658 = _zz_8659;
  assign _zz_8659 = ($signed(_zz_8660) >>> _zz_800);
  assign _zz_8660 = _zz_8661;
  assign _zz_8661 = ($signed(_zz_8663) + $signed(_zz_796));
  assign _zz_8662 = ({9'd0,data_mid_4_47_real} <<< 9);
  assign _zz_8663 = {{9{_zz_8662[26]}}, _zz_8662};
  assign _zz_8664 = fixTo_958_dout;
  assign _zz_8665 = _zz_8666[35 : 0];
  assign _zz_8666 = _zz_8667;
  assign _zz_8667 = ($signed(_zz_8668) >>> _zz_800);
  assign _zz_8668 = _zz_8669;
  assign _zz_8669 = ($signed(_zz_8671) + $signed(_zz_797));
  assign _zz_8670 = ({9'd0,data_mid_4_47_imag} <<< 9);
  assign _zz_8671 = {{9{_zz_8670[26]}}, _zz_8670};
  assign _zz_8672 = fixTo_959_dout;
  assign _zz_8673 = ($signed(twiddle_factor_table_31_real) + $signed(twiddle_factor_table_31_imag));
  assign _zz_8674 = ($signed(_zz_803) - $signed(_zz_8675));
  assign _zz_8675 = ($signed(_zz_8676) * $signed(twiddle_factor_table_31_imag));
  assign _zz_8676 = ($signed(data_mid_5_32_real) + $signed(data_mid_5_32_imag));
  assign _zz_8677 = fixTo_960_dout;
  assign _zz_8678 = ($signed(_zz_803) + $signed(_zz_8679));
  assign _zz_8679 = ($signed(_zz_8680) * $signed(twiddle_factor_table_31_real));
  assign _zz_8680 = ($signed(data_mid_5_32_imag) - $signed(data_mid_5_32_real));
  assign _zz_8681 = fixTo_961_dout;
  assign _zz_8682 = _zz_8683[35 : 0];
  assign _zz_8683 = _zz_8684;
  assign _zz_8684 = ($signed(_zz_8685) >>> _zz_804);
  assign _zz_8685 = _zz_8686;
  assign _zz_8686 = ($signed(_zz_8688) - $signed(_zz_801));
  assign _zz_8687 = ({9'd0,data_mid_5_0_real} <<< 9);
  assign _zz_8688 = {{9{_zz_8687[26]}}, _zz_8687};
  assign _zz_8689 = fixTo_962_dout;
  assign _zz_8690 = _zz_8691[35 : 0];
  assign _zz_8691 = _zz_8692;
  assign _zz_8692 = ($signed(_zz_8693) >>> _zz_804);
  assign _zz_8693 = _zz_8694;
  assign _zz_8694 = ($signed(_zz_8696) - $signed(_zz_802));
  assign _zz_8695 = ({9'd0,data_mid_5_0_imag} <<< 9);
  assign _zz_8696 = {{9{_zz_8695[26]}}, _zz_8695};
  assign _zz_8697 = fixTo_963_dout;
  assign _zz_8698 = _zz_8699[35 : 0];
  assign _zz_8699 = _zz_8700;
  assign _zz_8700 = ($signed(_zz_8701) >>> _zz_805);
  assign _zz_8701 = _zz_8702;
  assign _zz_8702 = ($signed(_zz_8704) + $signed(_zz_801));
  assign _zz_8703 = ({9'd0,data_mid_5_0_real} <<< 9);
  assign _zz_8704 = {{9{_zz_8703[26]}}, _zz_8703};
  assign _zz_8705 = fixTo_964_dout;
  assign _zz_8706 = _zz_8707[35 : 0];
  assign _zz_8707 = _zz_8708;
  assign _zz_8708 = ($signed(_zz_8709) >>> _zz_805);
  assign _zz_8709 = _zz_8710;
  assign _zz_8710 = ($signed(_zz_8712) + $signed(_zz_802));
  assign _zz_8711 = ({9'd0,data_mid_5_0_imag} <<< 9);
  assign _zz_8712 = {{9{_zz_8711[26]}}, _zz_8711};
  assign _zz_8713 = fixTo_965_dout;
  assign _zz_8714 = ($signed(twiddle_factor_table_32_real) + $signed(twiddle_factor_table_32_imag));
  assign _zz_8715 = ($signed(_zz_808) - $signed(_zz_8716));
  assign _zz_8716 = ($signed(_zz_8717) * $signed(twiddle_factor_table_32_imag));
  assign _zz_8717 = ($signed(data_mid_5_33_real) + $signed(data_mid_5_33_imag));
  assign _zz_8718 = fixTo_966_dout;
  assign _zz_8719 = ($signed(_zz_808) + $signed(_zz_8720));
  assign _zz_8720 = ($signed(_zz_8721) * $signed(twiddle_factor_table_32_real));
  assign _zz_8721 = ($signed(data_mid_5_33_imag) - $signed(data_mid_5_33_real));
  assign _zz_8722 = fixTo_967_dout;
  assign _zz_8723 = _zz_8724[35 : 0];
  assign _zz_8724 = _zz_8725;
  assign _zz_8725 = ($signed(_zz_8726) >>> _zz_809);
  assign _zz_8726 = _zz_8727;
  assign _zz_8727 = ($signed(_zz_8729) - $signed(_zz_806));
  assign _zz_8728 = ({9'd0,data_mid_5_1_real} <<< 9);
  assign _zz_8729 = {{9{_zz_8728[26]}}, _zz_8728};
  assign _zz_8730 = fixTo_968_dout;
  assign _zz_8731 = _zz_8732[35 : 0];
  assign _zz_8732 = _zz_8733;
  assign _zz_8733 = ($signed(_zz_8734) >>> _zz_809);
  assign _zz_8734 = _zz_8735;
  assign _zz_8735 = ($signed(_zz_8737) - $signed(_zz_807));
  assign _zz_8736 = ({9'd0,data_mid_5_1_imag} <<< 9);
  assign _zz_8737 = {{9{_zz_8736[26]}}, _zz_8736};
  assign _zz_8738 = fixTo_969_dout;
  assign _zz_8739 = _zz_8740[35 : 0];
  assign _zz_8740 = _zz_8741;
  assign _zz_8741 = ($signed(_zz_8742) >>> _zz_810);
  assign _zz_8742 = _zz_8743;
  assign _zz_8743 = ($signed(_zz_8745) + $signed(_zz_806));
  assign _zz_8744 = ({9'd0,data_mid_5_1_real} <<< 9);
  assign _zz_8745 = {{9{_zz_8744[26]}}, _zz_8744};
  assign _zz_8746 = fixTo_970_dout;
  assign _zz_8747 = _zz_8748[35 : 0];
  assign _zz_8748 = _zz_8749;
  assign _zz_8749 = ($signed(_zz_8750) >>> _zz_810);
  assign _zz_8750 = _zz_8751;
  assign _zz_8751 = ($signed(_zz_8753) + $signed(_zz_807));
  assign _zz_8752 = ({9'd0,data_mid_5_1_imag} <<< 9);
  assign _zz_8753 = {{9{_zz_8752[26]}}, _zz_8752};
  assign _zz_8754 = fixTo_971_dout;
  assign _zz_8755 = ($signed(twiddle_factor_table_33_real) + $signed(twiddle_factor_table_33_imag));
  assign _zz_8756 = ($signed(_zz_813) - $signed(_zz_8757));
  assign _zz_8757 = ($signed(_zz_8758) * $signed(twiddle_factor_table_33_imag));
  assign _zz_8758 = ($signed(data_mid_5_34_real) + $signed(data_mid_5_34_imag));
  assign _zz_8759 = fixTo_972_dout;
  assign _zz_8760 = ($signed(_zz_813) + $signed(_zz_8761));
  assign _zz_8761 = ($signed(_zz_8762) * $signed(twiddle_factor_table_33_real));
  assign _zz_8762 = ($signed(data_mid_5_34_imag) - $signed(data_mid_5_34_real));
  assign _zz_8763 = fixTo_973_dout;
  assign _zz_8764 = _zz_8765[35 : 0];
  assign _zz_8765 = _zz_8766;
  assign _zz_8766 = ($signed(_zz_8767) >>> _zz_814);
  assign _zz_8767 = _zz_8768;
  assign _zz_8768 = ($signed(_zz_8770) - $signed(_zz_811));
  assign _zz_8769 = ({9'd0,data_mid_5_2_real} <<< 9);
  assign _zz_8770 = {{9{_zz_8769[26]}}, _zz_8769};
  assign _zz_8771 = fixTo_974_dout;
  assign _zz_8772 = _zz_8773[35 : 0];
  assign _zz_8773 = _zz_8774;
  assign _zz_8774 = ($signed(_zz_8775) >>> _zz_814);
  assign _zz_8775 = _zz_8776;
  assign _zz_8776 = ($signed(_zz_8778) - $signed(_zz_812));
  assign _zz_8777 = ({9'd0,data_mid_5_2_imag} <<< 9);
  assign _zz_8778 = {{9{_zz_8777[26]}}, _zz_8777};
  assign _zz_8779 = fixTo_975_dout;
  assign _zz_8780 = _zz_8781[35 : 0];
  assign _zz_8781 = _zz_8782;
  assign _zz_8782 = ($signed(_zz_8783) >>> _zz_815);
  assign _zz_8783 = _zz_8784;
  assign _zz_8784 = ($signed(_zz_8786) + $signed(_zz_811));
  assign _zz_8785 = ({9'd0,data_mid_5_2_real} <<< 9);
  assign _zz_8786 = {{9{_zz_8785[26]}}, _zz_8785};
  assign _zz_8787 = fixTo_976_dout;
  assign _zz_8788 = _zz_8789[35 : 0];
  assign _zz_8789 = _zz_8790;
  assign _zz_8790 = ($signed(_zz_8791) >>> _zz_815);
  assign _zz_8791 = _zz_8792;
  assign _zz_8792 = ($signed(_zz_8794) + $signed(_zz_812));
  assign _zz_8793 = ({9'd0,data_mid_5_2_imag} <<< 9);
  assign _zz_8794 = {{9{_zz_8793[26]}}, _zz_8793};
  assign _zz_8795 = fixTo_977_dout;
  assign _zz_8796 = ($signed(twiddle_factor_table_34_real) + $signed(twiddle_factor_table_34_imag));
  assign _zz_8797 = ($signed(_zz_818) - $signed(_zz_8798));
  assign _zz_8798 = ($signed(_zz_8799) * $signed(twiddle_factor_table_34_imag));
  assign _zz_8799 = ($signed(data_mid_5_35_real) + $signed(data_mid_5_35_imag));
  assign _zz_8800 = fixTo_978_dout;
  assign _zz_8801 = ($signed(_zz_818) + $signed(_zz_8802));
  assign _zz_8802 = ($signed(_zz_8803) * $signed(twiddle_factor_table_34_real));
  assign _zz_8803 = ($signed(data_mid_5_35_imag) - $signed(data_mid_5_35_real));
  assign _zz_8804 = fixTo_979_dout;
  assign _zz_8805 = _zz_8806[35 : 0];
  assign _zz_8806 = _zz_8807;
  assign _zz_8807 = ($signed(_zz_8808) >>> _zz_819);
  assign _zz_8808 = _zz_8809;
  assign _zz_8809 = ($signed(_zz_8811) - $signed(_zz_816));
  assign _zz_8810 = ({9'd0,data_mid_5_3_real} <<< 9);
  assign _zz_8811 = {{9{_zz_8810[26]}}, _zz_8810};
  assign _zz_8812 = fixTo_980_dout;
  assign _zz_8813 = _zz_8814[35 : 0];
  assign _zz_8814 = _zz_8815;
  assign _zz_8815 = ($signed(_zz_8816) >>> _zz_819);
  assign _zz_8816 = _zz_8817;
  assign _zz_8817 = ($signed(_zz_8819) - $signed(_zz_817));
  assign _zz_8818 = ({9'd0,data_mid_5_3_imag} <<< 9);
  assign _zz_8819 = {{9{_zz_8818[26]}}, _zz_8818};
  assign _zz_8820 = fixTo_981_dout;
  assign _zz_8821 = _zz_8822[35 : 0];
  assign _zz_8822 = _zz_8823;
  assign _zz_8823 = ($signed(_zz_8824) >>> _zz_820);
  assign _zz_8824 = _zz_8825;
  assign _zz_8825 = ($signed(_zz_8827) + $signed(_zz_816));
  assign _zz_8826 = ({9'd0,data_mid_5_3_real} <<< 9);
  assign _zz_8827 = {{9{_zz_8826[26]}}, _zz_8826};
  assign _zz_8828 = fixTo_982_dout;
  assign _zz_8829 = _zz_8830[35 : 0];
  assign _zz_8830 = _zz_8831;
  assign _zz_8831 = ($signed(_zz_8832) >>> _zz_820);
  assign _zz_8832 = _zz_8833;
  assign _zz_8833 = ($signed(_zz_8835) + $signed(_zz_817));
  assign _zz_8834 = ({9'd0,data_mid_5_3_imag} <<< 9);
  assign _zz_8835 = {{9{_zz_8834[26]}}, _zz_8834};
  assign _zz_8836 = fixTo_983_dout;
  assign _zz_8837 = ($signed(twiddle_factor_table_35_real) + $signed(twiddle_factor_table_35_imag));
  assign _zz_8838 = ($signed(_zz_823) - $signed(_zz_8839));
  assign _zz_8839 = ($signed(_zz_8840) * $signed(twiddle_factor_table_35_imag));
  assign _zz_8840 = ($signed(data_mid_5_36_real) + $signed(data_mid_5_36_imag));
  assign _zz_8841 = fixTo_984_dout;
  assign _zz_8842 = ($signed(_zz_823) + $signed(_zz_8843));
  assign _zz_8843 = ($signed(_zz_8844) * $signed(twiddle_factor_table_35_real));
  assign _zz_8844 = ($signed(data_mid_5_36_imag) - $signed(data_mid_5_36_real));
  assign _zz_8845 = fixTo_985_dout;
  assign _zz_8846 = _zz_8847[35 : 0];
  assign _zz_8847 = _zz_8848;
  assign _zz_8848 = ($signed(_zz_8849) >>> _zz_824);
  assign _zz_8849 = _zz_8850;
  assign _zz_8850 = ($signed(_zz_8852) - $signed(_zz_821));
  assign _zz_8851 = ({9'd0,data_mid_5_4_real} <<< 9);
  assign _zz_8852 = {{9{_zz_8851[26]}}, _zz_8851};
  assign _zz_8853 = fixTo_986_dout;
  assign _zz_8854 = _zz_8855[35 : 0];
  assign _zz_8855 = _zz_8856;
  assign _zz_8856 = ($signed(_zz_8857) >>> _zz_824);
  assign _zz_8857 = _zz_8858;
  assign _zz_8858 = ($signed(_zz_8860) - $signed(_zz_822));
  assign _zz_8859 = ({9'd0,data_mid_5_4_imag} <<< 9);
  assign _zz_8860 = {{9{_zz_8859[26]}}, _zz_8859};
  assign _zz_8861 = fixTo_987_dout;
  assign _zz_8862 = _zz_8863[35 : 0];
  assign _zz_8863 = _zz_8864;
  assign _zz_8864 = ($signed(_zz_8865) >>> _zz_825);
  assign _zz_8865 = _zz_8866;
  assign _zz_8866 = ($signed(_zz_8868) + $signed(_zz_821));
  assign _zz_8867 = ({9'd0,data_mid_5_4_real} <<< 9);
  assign _zz_8868 = {{9{_zz_8867[26]}}, _zz_8867};
  assign _zz_8869 = fixTo_988_dout;
  assign _zz_8870 = _zz_8871[35 : 0];
  assign _zz_8871 = _zz_8872;
  assign _zz_8872 = ($signed(_zz_8873) >>> _zz_825);
  assign _zz_8873 = _zz_8874;
  assign _zz_8874 = ($signed(_zz_8876) + $signed(_zz_822));
  assign _zz_8875 = ({9'd0,data_mid_5_4_imag} <<< 9);
  assign _zz_8876 = {{9{_zz_8875[26]}}, _zz_8875};
  assign _zz_8877 = fixTo_989_dout;
  assign _zz_8878 = ($signed(twiddle_factor_table_36_real) + $signed(twiddle_factor_table_36_imag));
  assign _zz_8879 = ($signed(_zz_828) - $signed(_zz_8880));
  assign _zz_8880 = ($signed(_zz_8881) * $signed(twiddle_factor_table_36_imag));
  assign _zz_8881 = ($signed(data_mid_5_37_real) + $signed(data_mid_5_37_imag));
  assign _zz_8882 = fixTo_990_dout;
  assign _zz_8883 = ($signed(_zz_828) + $signed(_zz_8884));
  assign _zz_8884 = ($signed(_zz_8885) * $signed(twiddle_factor_table_36_real));
  assign _zz_8885 = ($signed(data_mid_5_37_imag) - $signed(data_mid_5_37_real));
  assign _zz_8886 = fixTo_991_dout;
  assign _zz_8887 = _zz_8888[35 : 0];
  assign _zz_8888 = _zz_8889;
  assign _zz_8889 = ($signed(_zz_8890) >>> _zz_829);
  assign _zz_8890 = _zz_8891;
  assign _zz_8891 = ($signed(_zz_8893) - $signed(_zz_826));
  assign _zz_8892 = ({9'd0,data_mid_5_5_real} <<< 9);
  assign _zz_8893 = {{9{_zz_8892[26]}}, _zz_8892};
  assign _zz_8894 = fixTo_992_dout;
  assign _zz_8895 = _zz_8896[35 : 0];
  assign _zz_8896 = _zz_8897;
  assign _zz_8897 = ($signed(_zz_8898) >>> _zz_829);
  assign _zz_8898 = _zz_8899;
  assign _zz_8899 = ($signed(_zz_8901) - $signed(_zz_827));
  assign _zz_8900 = ({9'd0,data_mid_5_5_imag} <<< 9);
  assign _zz_8901 = {{9{_zz_8900[26]}}, _zz_8900};
  assign _zz_8902 = fixTo_993_dout;
  assign _zz_8903 = _zz_8904[35 : 0];
  assign _zz_8904 = _zz_8905;
  assign _zz_8905 = ($signed(_zz_8906) >>> _zz_830);
  assign _zz_8906 = _zz_8907;
  assign _zz_8907 = ($signed(_zz_8909) + $signed(_zz_826));
  assign _zz_8908 = ({9'd0,data_mid_5_5_real} <<< 9);
  assign _zz_8909 = {{9{_zz_8908[26]}}, _zz_8908};
  assign _zz_8910 = fixTo_994_dout;
  assign _zz_8911 = _zz_8912[35 : 0];
  assign _zz_8912 = _zz_8913;
  assign _zz_8913 = ($signed(_zz_8914) >>> _zz_830);
  assign _zz_8914 = _zz_8915;
  assign _zz_8915 = ($signed(_zz_8917) + $signed(_zz_827));
  assign _zz_8916 = ({9'd0,data_mid_5_5_imag} <<< 9);
  assign _zz_8917 = {{9{_zz_8916[26]}}, _zz_8916};
  assign _zz_8918 = fixTo_995_dout;
  assign _zz_8919 = ($signed(twiddle_factor_table_37_real) + $signed(twiddle_factor_table_37_imag));
  assign _zz_8920 = ($signed(_zz_833) - $signed(_zz_8921));
  assign _zz_8921 = ($signed(_zz_8922) * $signed(twiddle_factor_table_37_imag));
  assign _zz_8922 = ($signed(data_mid_5_38_real) + $signed(data_mid_5_38_imag));
  assign _zz_8923 = fixTo_996_dout;
  assign _zz_8924 = ($signed(_zz_833) + $signed(_zz_8925));
  assign _zz_8925 = ($signed(_zz_8926) * $signed(twiddle_factor_table_37_real));
  assign _zz_8926 = ($signed(data_mid_5_38_imag) - $signed(data_mid_5_38_real));
  assign _zz_8927 = fixTo_997_dout;
  assign _zz_8928 = _zz_8929[35 : 0];
  assign _zz_8929 = _zz_8930;
  assign _zz_8930 = ($signed(_zz_8931) >>> _zz_834);
  assign _zz_8931 = _zz_8932;
  assign _zz_8932 = ($signed(_zz_8934) - $signed(_zz_831));
  assign _zz_8933 = ({9'd0,data_mid_5_6_real} <<< 9);
  assign _zz_8934 = {{9{_zz_8933[26]}}, _zz_8933};
  assign _zz_8935 = fixTo_998_dout;
  assign _zz_8936 = _zz_8937[35 : 0];
  assign _zz_8937 = _zz_8938;
  assign _zz_8938 = ($signed(_zz_8939) >>> _zz_834);
  assign _zz_8939 = _zz_8940;
  assign _zz_8940 = ($signed(_zz_8942) - $signed(_zz_832));
  assign _zz_8941 = ({9'd0,data_mid_5_6_imag} <<< 9);
  assign _zz_8942 = {{9{_zz_8941[26]}}, _zz_8941};
  assign _zz_8943 = fixTo_999_dout;
  assign _zz_8944 = _zz_8945[35 : 0];
  assign _zz_8945 = _zz_8946;
  assign _zz_8946 = ($signed(_zz_8947) >>> _zz_835);
  assign _zz_8947 = _zz_8948;
  assign _zz_8948 = ($signed(_zz_8950) + $signed(_zz_831));
  assign _zz_8949 = ({9'd0,data_mid_5_6_real} <<< 9);
  assign _zz_8950 = {{9{_zz_8949[26]}}, _zz_8949};
  assign _zz_8951 = fixTo_1000_dout;
  assign _zz_8952 = _zz_8953[35 : 0];
  assign _zz_8953 = _zz_8954;
  assign _zz_8954 = ($signed(_zz_8955) >>> _zz_835);
  assign _zz_8955 = _zz_8956;
  assign _zz_8956 = ($signed(_zz_8958) + $signed(_zz_832));
  assign _zz_8957 = ({9'd0,data_mid_5_6_imag} <<< 9);
  assign _zz_8958 = {{9{_zz_8957[26]}}, _zz_8957};
  assign _zz_8959 = fixTo_1001_dout;
  assign _zz_8960 = ($signed(twiddle_factor_table_38_real) + $signed(twiddle_factor_table_38_imag));
  assign _zz_8961 = ($signed(_zz_838) - $signed(_zz_8962));
  assign _zz_8962 = ($signed(_zz_8963) * $signed(twiddle_factor_table_38_imag));
  assign _zz_8963 = ($signed(data_mid_5_39_real) + $signed(data_mid_5_39_imag));
  assign _zz_8964 = fixTo_1002_dout;
  assign _zz_8965 = ($signed(_zz_838) + $signed(_zz_8966));
  assign _zz_8966 = ($signed(_zz_8967) * $signed(twiddle_factor_table_38_real));
  assign _zz_8967 = ($signed(data_mid_5_39_imag) - $signed(data_mid_5_39_real));
  assign _zz_8968 = fixTo_1003_dout;
  assign _zz_8969 = _zz_8970[35 : 0];
  assign _zz_8970 = _zz_8971;
  assign _zz_8971 = ($signed(_zz_8972) >>> _zz_839);
  assign _zz_8972 = _zz_8973;
  assign _zz_8973 = ($signed(_zz_8975) - $signed(_zz_836));
  assign _zz_8974 = ({9'd0,data_mid_5_7_real} <<< 9);
  assign _zz_8975 = {{9{_zz_8974[26]}}, _zz_8974};
  assign _zz_8976 = fixTo_1004_dout;
  assign _zz_8977 = _zz_8978[35 : 0];
  assign _zz_8978 = _zz_8979;
  assign _zz_8979 = ($signed(_zz_8980) >>> _zz_839);
  assign _zz_8980 = _zz_8981;
  assign _zz_8981 = ($signed(_zz_8983) - $signed(_zz_837));
  assign _zz_8982 = ({9'd0,data_mid_5_7_imag} <<< 9);
  assign _zz_8983 = {{9{_zz_8982[26]}}, _zz_8982};
  assign _zz_8984 = fixTo_1005_dout;
  assign _zz_8985 = _zz_8986[35 : 0];
  assign _zz_8986 = _zz_8987;
  assign _zz_8987 = ($signed(_zz_8988) >>> _zz_840);
  assign _zz_8988 = _zz_8989;
  assign _zz_8989 = ($signed(_zz_8991) + $signed(_zz_836));
  assign _zz_8990 = ({9'd0,data_mid_5_7_real} <<< 9);
  assign _zz_8991 = {{9{_zz_8990[26]}}, _zz_8990};
  assign _zz_8992 = fixTo_1006_dout;
  assign _zz_8993 = _zz_8994[35 : 0];
  assign _zz_8994 = _zz_8995;
  assign _zz_8995 = ($signed(_zz_8996) >>> _zz_840);
  assign _zz_8996 = _zz_8997;
  assign _zz_8997 = ($signed(_zz_8999) + $signed(_zz_837));
  assign _zz_8998 = ({9'd0,data_mid_5_7_imag} <<< 9);
  assign _zz_8999 = {{9{_zz_8998[26]}}, _zz_8998};
  assign _zz_9000 = fixTo_1007_dout;
  assign _zz_9001 = ($signed(twiddle_factor_table_39_real) + $signed(twiddle_factor_table_39_imag));
  assign _zz_9002 = ($signed(_zz_843) - $signed(_zz_9003));
  assign _zz_9003 = ($signed(_zz_9004) * $signed(twiddle_factor_table_39_imag));
  assign _zz_9004 = ($signed(data_mid_5_40_real) + $signed(data_mid_5_40_imag));
  assign _zz_9005 = fixTo_1008_dout;
  assign _zz_9006 = ($signed(_zz_843) + $signed(_zz_9007));
  assign _zz_9007 = ($signed(_zz_9008) * $signed(twiddle_factor_table_39_real));
  assign _zz_9008 = ($signed(data_mid_5_40_imag) - $signed(data_mid_5_40_real));
  assign _zz_9009 = fixTo_1009_dout;
  assign _zz_9010 = _zz_9011[35 : 0];
  assign _zz_9011 = _zz_9012;
  assign _zz_9012 = ($signed(_zz_9013) >>> _zz_844);
  assign _zz_9013 = _zz_9014;
  assign _zz_9014 = ($signed(_zz_9016) - $signed(_zz_841));
  assign _zz_9015 = ({9'd0,data_mid_5_8_real} <<< 9);
  assign _zz_9016 = {{9{_zz_9015[26]}}, _zz_9015};
  assign _zz_9017 = fixTo_1010_dout;
  assign _zz_9018 = _zz_9019[35 : 0];
  assign _zz_9019 = _zz_9020;
  assign _zz_9020 = ($signed(_zz_9021) >>> _zz_844);
  assign _zz_9021 = _zz_9022;
  assign _zz_9022 = ($signed(_zz_9024) - $signed(_zz_842));
  assign _zz_9023 = ({9'd0,data_mid_5_8_imag} <<< 9);
  assign _zz_9024 = {{9{_zz_9023[26]}}, _zz_9023};
  assign _zz_9025 = fixTo_1011_dout;
  assign _zz_9026 = _zz_9027[35 : 0];
  assign _zz_9027 = _zz_9028;
  assign _zz_9028 = ($signed(_zz_9029) >>> _zz_845);
  assign _zz_9029 = _zz_9030;
  assign _zz_9030 = ($signed(_zz_9032) + $signed(_zz_841));
  assign _zz_9031 = ({9'd0,data_mid_5_8_real} <<< 9);
  assign _zz_9032 = {{9{_zz_9031[26]}}, _zz_9031};
  assign _zz_9033 = fixTo_1012_dout;
  assign _zz_9034 = _zz_9035[35 : 0];
  assign _zz_9035 = _zz_9036;
  assign _zz_9036 = ($signed(_zz_9037) >>> _zz_845);
  assign _zz_9037 = _zz_9038;
  assign _zz_9038 = ($signed(_zz_9040) + $signed(_zz_842));
  assign _zz_9039 = ({9'd0,data_mid_5_8_imag} <<< 9);
  assign _zz_9040 = {{9{_zz_9039[26]}}, _zz_9039};
  assign _zz_9041 = fixTo_1013_dout;
  assign _zz_9042 = ($signed(twiddle_factor_table_40_real) + $signed(twiddle_factor_table_40_imag));
  assign _zz_9043 = ($signed(_zz_848) - $signed(_zz_9044));
  assign _zz_9044 = ($signed(_zz_9045) * $signed(twiddle_factor_table_40_imag));
  assign _zz_9045 = ($signed(data_mid_5_41_real) + $signed(data_mid_5_41_imag));
  assign _zz_9046 = fixTo_1014_dout;
  assign _zz_9047 = ($signed(_zz_848) + $signed(_zz_9048));
  assign _zz_9048 = ($signed(_zz_9049) * $signed(twiddle_factor_table_40_real));
  assign _zz_9049 = ($signed(data_mid_5_41_imag) - $signed(data_mid_5_41_real));
  assign _zz_9050 = fixTo_1015_dout;
  assign _zz_9051 = _zz_9052[35 : 0];
  assign _zz_9052 = _zz_9053;
  assign _zz_9053 = ($signed(_zz_9054) >>> _zz_849);
  assign _zz_9054 = _zz_9055;
  assign _zz_9055 = ($signed(_zz_9057) - $signed(_zz_846));
  assign _zz_9056 = ({9'd0,data_mid_5_9_real} <<< 9);
  assign _zz_9057 = {{9{_zz_9056[26]}}, _zz_9056};
  assign _zz_9058 = fixTo_1016_dout;
  assign _zz_9059 = _zz_9060[35 : 0];
  assign _zz_9060 = _zz_9061;
  assign _zz_9061 = ($signed(_zz_9062) >>> _zz_849);
  assign _zz_9062 = _zz_9063;
  assign _zz_9063 = ($signed(_zz_9065) - $signed(_zz_847));
  assign _zz_9064 = ({9'd0,data_mid_5_9_imag} <<< 9);
  assign _zz_9065 = {{9{_zz_9064[26]}}, _zz_9064};
  assign _zz_9066 = fixTo_1017_dout;
  assign _zz_9067 = _zz_9068[35 : 0];
  assign _zz_9068 = _zz_9069;
  assign _zz_9069 = ($signed(_zz_9070) >>> _zz_850);
  assign _zz_9070 = _zz_9071;
  assign _zz_9071 = ($signed(_zz_9073) + $signed(_zz_846));
  assign _zz_9072 = ({9'd0,data_mid_5_9_real} <<< 9);
  assign _zz_9073 = {{9{_zz_9072[26]}}, _zz_9072};
  assign _zz_9074 = fixTo_1018_dout;
  assign _zz_9075 = _zz_9076[35 : 0];
  assign _zz_9076 = _zz_9077;
  assign _zz_9077 = ($signed(_zz_9078) >>> _zz_850);
  assign _zz_9078 = _zz_9079;
  assign _zz_9079 = ($signed(_zz_9081) + $signed(_zz_847));
  assign _zz_9080 = ({9'd0,data_mid_5_9_imag} <<< 9);
  assign _zz_9081 = {{9{_zz_9080[26]}}, _zz_9080};
  assign _zz_9082 = fixTo_1019_dout;
  assign _zz_9083 = ($signed(twiddle_factor_table_41_real) + $signed(twiddle_factor_table_41_imag));
  assign _zz_9084 = ($signed(_zz_853) - $signed(_zz_9085));
  assign _zz_9085 = ($signed(_zz_9086) * $signed(twiddle_factor_table_41_imag));
  assign _zz_9086 = ($signed(data_mid_5_42_real) + $signed(data_mid_5_42_imag));
  assign _zz_9087 = fixTo_1020_dout;
  assign _zz_9088 = ($signed(_zz_853) + $signed(_zz_9089));
  assign _zz_9089 = ($signed(_zz_9090) * $signed(twiddle_factor_table_41_real));
  assign _zz_9090 = ($signed(data_mid_5_42_imag) - $signed(data_mid_5_42_real));
  assign _zz_9091 = fixTo_1021_dout;
  assign _zz_9092 = _zz_9093[35 : 0];
  assign _zz_9093 = _zz_9094;
  assign _zz_9094 = ($signed(_zz_9095) >>> _zz_854);
  assign _zz_9095 = _zz_9096;
  assign _zz_9096 = ($signed(_zz_9098) - $signed(_zz_851));
  assign _zz_9097 = ({9'd0,data_mid_5_10_real} <<< 9);
  assign _zz_9098 = {{9{_zz_9097[26]}}, _zz_9097};
  assign _zz_9099 = fixTo_1022_dout;
  assign _zz_9100 = _zz_9101[35 : 0];
  assign _zz_9101 = _zz_9102;
  assign _zz_9102 = ($signed(_zz_9103) >>> _zz_854);
  assign _zz_9103 = _zz_9104;
  assign _zz_9104 = ($signed(_zz_9106) - $signed(_zz_852));
  assign _zz_9105 = ({9'd0,data_mid_5_10_imag} <<< 9);
  assign _zz_9106 = {{9{_zz_9105[26]}}, _zz_9105};
  assign _zz_9107 = fixTo_1023_dout;
  assign _zz_9108 = _zz_9109[35 : 0];
  assign _zz_9109 = _zz_9110;
  assign _zz_9110 = ($signed(_zz_9111) >>> _zz_855);
  assign _zz_9111 = _zz_9112;
  assign _zz_9112 = ($signed(_zz_9114) + $signed(_zz_851));
  assign _zz_9113 = ({9'd0,data_mid_5_10_real} <<< 9);
  assign _zz_9114 = {{9{_zz_9113[26]}}, _zz_9113};
  assign _zz_9115 = fixTo_1024_dout;
  assign _zz_9116 = _zz_9117[35 : 0];
  assign _zz_9117 = _zz_9118;
  assign _zz_9118 = ($signed(_zz_9119) >>> _zz_855);
  assign _zz_9119 = _zz_9120;
  assign _zz_9120 = ($signed(_zz_9122) + $signed(_zz_852));
  assign _zz_9121 = ({9'd0,data_mid_5_10_imag} <<< 9);
  assign _zz_9122 = {{9{_zz_9121[26]}}, _zz_9121};
  assign _zz_9123 = fixTo_1025_dout;
  assign _zz_9124 = ($signed(twiddle_factor_table_42_real) + $signed(twiddle_factor_table_42_imag));
  assign _zz_9125 = ($signed(_zz_858) - $signed(_zz_9126));
  assign _zz_9126 = ($signed(_zz_9127) * $signed(twiddle_factor_table_42_imag));
  assign _zz_9127 = ($signed(data_mid_5_43_real) + $signed(data_mid_5_43_imag));
  assign _zz_9128 = fixTo_1026_dout;
  assign _zz_9129 = ($signed(_zz_858) + $signed(_zz_9130));
  assign _zz_9130 = ($signed(_zz_9131) * $signed(twiddle_factor_table_42_real));
  assign _zz_9131 = ($signed(data_mid_5_43_imag) - $signed(data_mid_5_43_real));
  assign _zz_9132 = fixTo_1027_dout;
  assign _zz_9133 = _zz_9134[35 : 0];
  assign _zz_9134 = _zz_9135;
  assign _zz_9135 = ($signed(_zz_9136) >>> _zz_859);
  assign _zz_9136 = _zz_9137;
  assign _zz_9137 = ($signed(_zz_9139) - $signed(_zz_856));
  assign _zz_9138 = ({9'd0,data_mid_5_11_real} <<< 9);
  assign _zz_9139 = {{9{_zz_9138[26]}}, _zz_9138};
  assign _zz_9140 = fixTo_1028_dout;
  assign _zz_9141 = _zz_9142[35 : 0];
  assign _zz_9142 = _zz_9143;
  assign _zz_9143 = ($signed(_zz_9144) >>> _zz_859);
  assign _zz_9144 = _zz_9145;
  assign _zz_9145 = ($signed(_zz_9147) - $signed(_zz_857));
  assign _zz_9146 = ({9'd0,data_mid_5_11_imag} <<< 9);
  assign _zz_9147 = {{9{_zz_9146[26]}}, _zz_9146};
  assign _zz_9148 = fixTo_1029_dout;
  assign _zz_9149 = _zz_9150[35 : 0];
  assign _zz_9150 = _zz_9151;
  assign _zz_9151 = ($signed(_zz_9152) >>> _zz_860);
  assign _zz_9152 = _zz_9153;
  assign _zz_9153 = ($signed(_zz_9155) + $signed(_zz_856));
  assign _zz_9154 = ({9'd0,data_mid_5_11_real} <<< 9);
  assign _zz_9155 = {{9{_zz_9154[26]}}, _zz_9154};
  assign _zz_9156 = fixTo_1030_dout;
  assign _zz_9157 = _zz_9158[35 : 0];
  assign _zz_9158 = _zz_9159;
  assign _zz_9159 = ($signed(_zz_9160) >>> _zz_860);
  assign _zz_9160 = _zz_9161;
  assign _zz_9161 = ($signed(_zz_9163) + $signed(_zz_857));
  assign _zz_9162 = ({9'd0,data_mid_5_11_imag} <<< 9);
  assign _zz_9163 = {{9{_zz_9162[26]}}, _zz_9162};
  assign _zz_9164 = fixTo_1031_dout;
  assign _zz_9165 = ($signed(twiddle_factor_table_43_real) + $signed(twiddle_factor_table_43_imag));
  assign _zz_9166 = ($signed(_zz_863) - $signed(_zz_9167));
  assign _zz_9167 = ($signed(_zz_9168) * $signed(twiddle_factor_table_43_imag));
  assign _zz_9168 = ($signed(data_mid_5_44_real) + $signed(data_mid_5_44_imag));
  assign _zz_9169 = fixTo_1032_dout;
  assign _zz_9170 = ($signed(_zz_863) + $signed(_zz_9171));
  assign _zz_9171 = ($signed(_zz_9172) * $signed(twiddle_factor_table_43_real));
  assign _zz_9172 = ($signed(data_mid_5_44_imag) - $signed(data_mid_5_44_real));
  assign _zz_9173 = fixTo_1033_dout;
  assign _zz_9174 = _zz_9175[35 : 0];
  assign _zz_9175 = _zz_9176;
  assign _zz_9176 = ($signed(_zz_9177) >>> _zz_864);
  assign _zz_9177 = _zz_9178;
  assign _zz_9178 = ($signed(_zz_9180) - $signed(_zz_861));
  assign _zz_9179 = ({9'd0,data_mid_5_12_real} <<< 9);
  assign _zz_9180 = {{9{_zz_9179[26]}}, _zz_9179};
  assign _zz_9181 = fixTo_1034_dout;
  assign _zz_9182 = _zz_9183[35 : 0];
  assign _zz_9183 = _zz_9184;
  assign _zz_9184 = ($signed(_zz_9185) >>> _zz_864);
  assign _zz_9185 = _zz_9186;
  assign _zz_9186 = ($signed(_zz_9188) - $signed(_zz_862));
  assign _zz_9187 = ({9'd0,data_mid_5_12_imag} <<< 9);
  assign _zz_9188 = {{9{_zz_9187[26]}}, _zz_9187};
  assign _zz_9189 = fixTo_1035_dout;
  assign _zz_9190 = _zz_9191[35 : 0];
  assign _zz_9191 = _zz_9192;
  assign _zz_9192 = ($signed(_zz_9193) >>> _zz_865);
  assign _zz_9193 = _zz_9194;
  assign _zz_9194 = ($signed(_zz_9196) + $signed(_zz_861));
  assign _zz_9195 = ({9'd0,data_mid_5_12_real} <<< 9);
  assign _zz_9196 = {{9{_zz_9195[26]}}, _zz_9195};
  assign _zz_9197 = fixTo_1036_dout;
  assign _zz_9198 = _zz_9199[35 : 0];
  assign _zz_9199 = _zz_9200;
  assign _zz_9200 = ($signed(_zz_9201) >>> _zz_865);
  assign _zz_9201 = _zz_9202;
  assign _zz_9202 = ($signed(_zz_9204) + $signed(_zz_862));
  assign _zz_9203 = ({9'd0,data_mid_5_12_imag} <<< 9);
  assign _zz_9204 = {{9{_zz_9203[26]}}, _zz_9203};
  assign _zz_9205 = fixTo_1037_dout;
  assign _zz_9206 = ($signed(twiddle_factor_table_44_real) + $signed(twiddle_factor_table_44_imag));
  assign _zz_9207 = ($signed(_zz_868) - $signed(_zz_9208));
  assign _zz_9208 = ($signed(_zz_9209) * $signed(twiddle_factor_table_44_imag));
  assign _zz_9209 = ($signed(data_mid_5_45_real) + $signed(data_mid_5_45_imag));
  assign _zz_9210 = fixTo_1038_dout;
  assign _zz_9211 = ($signed(_zz_868) + $signed(_zz_9212));
  assign _zz_9212 = ($signed(_zz_9213) * $signed(twiddle_factor_table_44_real));
  assign _zz_9213 = ($signed(data_mid_5_45_imag) - $signed(data_mid_5_45_real));
  assign _zz_9214 = fixTo_1039_dout;
  assign _zz_9215 = _zz_9216[35 : 0];
  assign _zz_9216 = _zz_9217;
  assign _zz_9217 = ($signed(_zz_9218) >>> _zz_869);
  assign _zz_9218 = _zz_9219;
  assign _zz_9219 = ($signed(_zz_9221) - $signed(_zz_866));
  assign _zz_9220 = ({9'd0,data_mid_5_13_real} <<< 9);
  assign _zz_9221 = {{9{_zz_9220[26]}}, _zz_9220};
  assign _zz_9222 = fixTo_1040_dout;
  assign _zz_9223 = _zz_9224[35 : 0];
  assign _zz_9224 = _zz_9225;
  assign _zz_9225 = ($signed(_zz_9226) >>> _zz_869);
  assign _zz_9226 = _zz_9227;
  assign _zz_9227 = ($signed(_zz_9229) - $signed(_zz_867));
  assign _zz_9228 = ({9'd0,data_mid_5_13_imag} <<< 9);
  assign _zz_9229 = {{9{_zz_9228[26]}}, _zz_9228};
  assign _zz_9230 = fixTo_1041_dout;
  assign _zz_9231 = _zz_9232[35 : 0];
  assign _zz_9232 = _zz_9233;
  assign _zz_9233 = ($signed(_zz_9234) >>> _zz_870);
  assign _zz_9234 = _zz_9235;
  assign _zz_9235 = ($signed(_zz_9237) + $signed(_zz_866));
  assign _zz_9236 = ({9'd0,data_mid_5_13_real} <<< 9);
  assign _zz_9237 = {{9{_zz_9236[26]}}, _zz_9236};
  assign _zz_9238 = fixTo_1042_dout;
  assign _zz_9239 = _zz_9240[35 : 0];
  assign _zz_9240 = _zz_9241;
  assign _zz_9241 = ($signed(_zz_9242) >>> _zz_870);
  assign _zz_9242 = _zz_9243;
  assign _zz_9243 = ($signed(_zz_9245) + $signed(_zz_867));
  assign _zz_9244 = ({9'd0,data_mid_5_13_imag} <<< 9);
  assign _zz_9245 = {{9{_zz_9244[26]}}, _zz_9244};
  assign _zz_9246 = fixTo_1043_dout;
  assign _zz_9247 = ($signed(twiddle_factor_table_45_real) + $signed(twiddle_factor_table_45_imag));
  assign _zz_9248 = ($signed(_zz_873) - $signed(_zz_9249));
  assign _zz_9249 = ($signed(_zz_9250) * $signed(twiddle_factor_table_45_imag));
  assign _zz_9250 = ($signed(data_mid_5_46_real) + $signed(data_mid_5_46_imag));
  assign _zz_9251 = fixTo_1044_dout;
  assign _zz_9252 = ($signed(_zz_873) + $signed(_zz_9253));
  assign _zz_9253 = ($signed(_zz_9254) * $signed(twiddle_factor_table_45_real));
  assign _zz_9254 = ($signed(data_mid_5_46_imag) - $signed(data_mid_5_46_real));
  assign _zz_9255 = fixTo_1045_dout;
  assign _zz_9256 = _zz_9257[35 : 0];
  assign _zz_9257 = _zz_9258;
  assign _zz_9258 = ($signed(_zz_9259) >>> _zz_874);
  assign _zz_9259 = _zz_9260;
  assign _zz_9260 = ($signed(_zz_9262) - $signed(_zz_871));
  assign _zz_9261 = ({9'd0,data_mid_5_14_real} <<< 9);
  assign _zz_9262 = {{9{_zz_9261[26]}}, _zz_9261};
  assign _zz_9263 = fixTo_1046_dout;
  assign _zz_9264 = _zz_9265[35 : 0];
  assign _zz_9265 = _zz_9266;
  assign _zz_9266 = ($signed(_zz_9267) >>> _zz_874);
  assign _zz_9267 = _zz_9268;
  assign _zz_9268 = ($signed(_zz_9270) - $signed(_zz_872));
  assign _zz_9269 = ({9'd0,data_mid_5_14_imag} <<< 9);
  assign _zz_9270 = {{9{_zz_9269[26]}}, _zz_9269};
  assign _zz_9271 = fixTo_1047_dout;
  assign _zz_9272 = _zz_9273[35 : 0];
  assign _zz_9273 = _zz_9274;
  assign _zz_9274 = ($signed(_zz_9275) >>> _zz_875);
  assign _zz_9275 = _zz_9276;
  assign _zz_9276 = ($signed(_zz_9278) + $signed(_zz_871));
  assign _zz_9277 = ({9'd0,data_mid_5_14_real} <<< 9);
  assign _zz_9278 = {{9{_zz_9277[26]}}, _zz_9277};
  assign _zz_9279 = fixTo_1048_dout;
  assign _zz_9280 = _zz_9281[35 : 0];
  assign _zz_9281 = _zz_9282;
  assign _zz_9282 = ($signed(_zz_9283) >>> _zz_875);
  assign _zz_9283 = _zz_9284;
  assign _zz_9284 = ($signed(_zz_9286) + $signed(_zz_872));
  assign _zz_9285 = ({9'd0,data_mid_5_14_imag} <<< 9);
  assign _zz_9286 = {{9{_zz_9285[26]}}, _zz_9285};
  assign _zz_9287 = fixTo_1049_dout;
  assign _zz_9288 = ($signed(twiddle_factor_table_46_real) + $signed(twiddle_factor_table_46_imag));
  assign _zz_9289 = ($signed(_zz_878) - $signed(_zz_9290));
  assign _zz_9290 = ($signed(_zz_9291) * $signed(twiddle_factor_table_46_imag));
  assign _zz_9291 = ($signed(data_mid_5_47_real) + $signed(data_mid_5_47_imag));
  assign _zz_9292 = fixTo_1050_dout;
  assign _zz_9293 = ($signed(_zz_878) + $signed(_zz_9294));
  assign _zz_9294 = ($signed(_zz_9295) * $signed(twiddle_factor_table_46_real));
  assign _zz_9295 = ($signed(data_mid_5_47_imag) - $signed(data_mid_5_47_real));
  assign _zz_9296 = fixTo_1051_dout;
  assign _zz_9297 = _zz_9298[35 : 0];
  assign _zz_9298 = _zz_9299;
  assign _zz_9299 = ($signed(_zz_9300) >>> _zz_879);
  assign _zz_9300 = _zz_9301;
  assign _zz_9301 = ($signed(_zz_9303) - $signed(_zz_876));
  assign _zz_9302 = ({9'd0,data_mid_5_15_real} <<< 9);
  assign _zz_9303 = {{9{_zz_9302[26]}}, _zz_9302};
  assign _zz_9304 = fixTo_1052_dout;
  assign _zz_9305 = _zz_9306[35 : 0];
  assign _zz_9306 = _zz_9307;
  assign _zz_9307 = ($signed(_zz_9308) >>> _zz_879);
  assign _zz_9308 = _zz_9309;
  assign _zz_9309 = ($signed(_zz_9311) - $signed(_zz_877));
  assign _zz_9310 = ({9'd0,data_mid_5_15_imag} <<< 9);
  assign _zz_9311 = {{9{_zz_9310[26]}}, _zz_9310};
  assign _zz_9312 = fixTo_1053_dout;
  assign _zz_9313 = _zz_9314[35 : 0];
  assign _zz_9314 = _zz_9315;
  assign _zz_9315 = ($signed(_zz_9316) >>> _zz_880);
  assign _zz_9316 = _zz_9317;
  assign _zz_9317 = ($signed(_zz_9319) + $signed(_zz_876));
  assign _zz_9318 = ({9'd0,data_mid_5_15_real} <<< 9);
  assign _zz_9319 = {{9{_zz_9318[26]}}, _zz_9318};
  assign _zz_9320 = fixTo_1054_dout;
  assign _zz_9321 = _zz_9322[35 : 0];
  assign _zz_9322 = _zz_9323;
  assign _zz_9323 = ($signed(_zz_9324) >>> _zz_880);
  assign _zz_9324 = _zz_9325;
  assign _zz_9325 = ($signed(_zz_9327) + $signed(_zz_877));
  assign _zz_9326 = ({9'd0,data_mid_5_15_imag} <<< 9);
  assign _zz_9327 = {{9{_zz_9326[26]}}, _zz_9326};
  assign _zz_9328 = fixTo_1055_dout;
  assign _zz_9329 = ($signed(twiddle_factor_table_47_real) + $signed(twiddle_factor_table_47_imag));
  assign _zz_9330 = ($signed(_zz_883) - $signed(_zz_9331));
  assign _zz_9331 = ($signed(_zz_9332) * $signed(twiddle_factor_table_47_imag));
  assign _zz_9332 = ($signed(data_mid_5_48_real) + $signed(data_mid_5_48_imag));
  assign _zz_9333 = fixTo_1056_dout;
  assign _zz_9334 = ($signed(_zz_883) + $signed(_zz_9335));
  assign _zz_9335 = ($signed(_zz_9336) * $signed(twiddle_factor_table_47_real));
  assign _zz_9336 = ($signed(data_mid_5_48_imag) - $signed(data_mid_5_48_real));
  assign _zz_9337 = fixTo_1057_dout;
  assign _zz_9338 = _zz_9339[35 : 0];
  assign _zz_9339 = _zz_9340;
  assign _zz_9340 = ($signed(_zz_9341) >>> _zz_884);
  assign _zz_9341 = _zz_9342;
  assign _zz_9342 = ($signed(_zz_9344) - $signed(_zz_881));
  assign _zz_9343 = ({9'd0,data_mid_5_16_real} <<< 9);
  assign _zz_9344 = {{9{_zz_9343[26]}}, _zz_9343};
  assign _zz_9345 = fixTo_1058_dout;
  assign _zz_9346 = _zz_9347[35 : 0];
  assign _zz_9347 = _zz_9348;
  assign _zz_9348 = ($signed(_zz_9349) >>> _zz_884);
  assign _zz_9349 = _zz_9350;
  assign _zz_9350 = ($signed(_zz_9352) - $signed(_zz_882));
  assign _zz_9351 = ({9'd0,data_mid_5_16_imag} <<< 9);
  assign _zz_9352 = {{9{_zz_9351[26]}}, _zz_9351};
  assign _zz_9353 = fixTo_1059_dout;
  assign _zz_9354 = _zz_9355[35 : 0];
  assign _zz_9355 = _zz_9356;
  assign _zz_9356 = ($signed(_zz_9357) >>> _zz_885);
  assign _zz_9357 = _zz_9358;
  assign _zz_9358 = ($signed(_zz_9360) + $signed(_zz_881));
  assign _zz_9359 = ({9'd0,data_mid_5_16_real} <<< 9);
  assign _zz_9360 = {{9{_zz_9359[26]}}, _zz_9359};
  assign _zz_9361 = fixTo_1060_dout;
  assign _zz_9362 = _zz_9363[35 : 0];
  assign _zz_9363 = _zz_9364;
  assign _zz_9364 = ($signed(_zz_9365) >>> _zz_885);
  assign _zz_9365 = _zz_9366;
  assign _zz_9366 = ($signed(_zz_9368) + $signed(_zz_882));
  assign _zz_9367 = ({9'd0,data_mid_5_16_imag} <<< 9);
  assign _zz_9368 = {{9{_zz_9367[26]}}, _zz_9367};
  assign _zz_9369 = fixTo_1061_dout;
  assign _zz_9370 = ($signed(twiddle_factor_table_48_real) + $signed(twiddle_factor_table_48_imag));
  assign _zz_9371 = ($signed(_zz_888) - $signed(_zz_9372));
  assign _zz_9372 = ($signed(_zz_9373) * $signed(twiddle_factor_table_48_imag));
  assign _zz_9373 = ($signed(data_mid_5_49_real) + $signed(data_mid_5_49_imag));
  assign _zz_9374 = fixTo_1062_dout;
  assign _zz_9375 = ($signed(_zz_888) + $signed(_zz_9376));
  assign _zz_9376 = ($signed(_zz_9377) * $signed(twiddle_factor_table_48_real));
  assign _zz_9377 = ($signed(data_mid_5_49_imag) - $signed(data_mid_5_49_real));
  assign _zz_9378 = fixTo_1063_dout;
  assign _zz_9379 = _zz_9380[35 : 0];
  assign _zz_9380 = _zz_9381;
  assign _zz_9381 = ($signed(_zz_9382) >>> _zz_889);
  assign _zz_9382 = _zz_9383;
  assign _zz_9383 = ($signed(_zz_9385) - $signed(_zz_886));
  assign _zz_9384 = ({9'd0,data_mid_5_17_real} <<< 9);
  assign _zz_9385 = {{9{_zz_9384[26]}}, _zz_9384};
  assign _zz_9386 = fixTo_1064_dout;
  assign _zz_9387 = _zz_9388[35 : 0];
  assign _zz_9388 = _zz_9389;
  assign _zz_9389 = ($signed(_zz_9390) >>> _zz_889);
  assign _zz_9390 = _zz_9391;
  assign _zz_9391 = ($signed(_zz_9393) - $signed(_zz_887));
  assign _zz_9392 = ({9'd0,data_mid_5_17_imag} <<< 9);
  assign _zz_9393 = {{9{_zz_9392[26]}}, _zz_9392};
  assign _zz_9394 = fixTo_1065_dout;
  assign _zz_9395 = _zz_9396[35 : 0];
  assign _zz_9396 = _zz_9397;
  assign _zz_9397 = ($signed(_zz_9398) >>> _zz_890);
  assign _zz_9398 = _zz_9399;
  assign _zz_9399 = ($signed(_zz_9401) + $signed(_zz_886));
  assign _zz_9400 = ({9'd0,data_mid_5_17_real} <<< 9);
  assign _zz_9401 = {{9{_zz_9400[26]}}, _zz_9400};
  assign _zz_9402 = fixTo_1066_dout;
  assign _zz_9403 = _zz_9404[35 : 0];
  assign _zz_9404 = _zz_9405;
  assign _zz_9405 = ($signed(_zz_9406) >>> _zz_890);
  assign _zz_9406 = _zz_9407;
  assign _zz_9407 = ($signed(_zz_9409) + $signed(_zz_887));
  assign _zz_9408 = ({9'd0,data_mid_5_17_imag} <<< 9);
  assign _zz_9409 = {{9{_zz_9408[26]}}, _zz_9408};
  assign _zz_9410 = fixTo_1067_dout;
  assign _zz_9411 = ($signed(twiddle_factor_table_49_real) + $signed(twiddle_factor_table_49_imag));
  assign _zz_9412 = ($signed(_zz_893) - $signed(_zz_9413));
  assign _zz_9413 = ($signed(_zz_9414) * $signed(twiddle_factor_table_49_imag));
  assign _zz_9414 = ($signed(data_mid_5_50_real) + $signed(data_mid_5_50_imag));
  assign _zz_9415 = fixTo_1068_dout;
  assign _zz_9416 = ($signed(_zz_893) + $signed(_zz_9417));
  assign _zz_9417 = ($signed(_zz_9418) * $signed(twiddle_factor_table_49_real));
  assign _zz_9418 = ($signed(data_mid_5_50_imag) - $signed(data_mid_5_50_real));
  assign _zz_9419 = fixTo_1069_dout;
  assign _zz_9420 = _zz_9421[35 : 0];
  assign _zz_9421 = _zz_9422;
  assign _zz_9422 = ($signed(_zz_9423) >>> _zz_894);
  assign _zz_9423 = _zz_9424;
  assign _zz_9424 = ($signed(_zz_9426) - $signed(_zz_891));
  assign _zz_9425 = ({9'd0,data_mid_5_18_real} <<< 9);
  assign _zz_9426 = {{9{_zz_9425[26]}}, _zz_9425};
  assign _zz_9427 = fixTo_1070_dout;
  assign _zz_9428 = _zz_9429[35 : 0];
  assign _zz_9429 = _zz_9430;
  assign _zz_9430 = ($signed(_zz_9431) >>> _zz_894);
  assign _zz_9431 = _zz_9432;
  assign _zz_9432 = ($signed(_zz_9434) - $signed(_zz_892));
  assign _zz_9433 = ({9'd0,data_mid_5_18_imag} <<< 9);
  assign _zz_9434 = {{9{_zz_9433[26]}}, _zz_9433};
  assign _zz_9435 = fixTo_1071_dout;
  assign _zz_9436 = _zz_9437[35 : 0];
  assign _zz_9437 = _zz_9438;
  assign _zz_9438 = ($signed(_zz_9439) >>> _zz_895);
  assign _zz_9439 = _zz_9440;
  assign _zz_9440 = ($signed(_zz_9442) + $signed(_zz_891));
  assign _zz_9441 = ({9'd0,data_mid_5_18_real} <<< 9);
  assign _zz_9442 = {{9{_zz_9441[26]}}, _zz_9441};
  assign _zz_9443 = fixTo_1072_dout;
  assign _zz_9444 = _zz_9445[35 : 0];
  assign _zz_9445 = _zz_9446;
  assign _zz_9446 = ($signed(_zz_9447) >>> _zz_895);
  assign _zz_9447 = _zz_9448;
  assign _zz_9448 = ($signed(_zz_9450) + $signed(_zz_892));
  assign _zz_9449 = ({9'd0,data_mid_5_18_imag} <<< 9);
  assign _zz_9450 = {{9{_zz_9449[26]}}, _zz_9449};
  assign _zz_9451 = fixTo_1073_dout;
  assign _zz_9452 = ($signed(twiddle_factor_table_50_real) + $signed(twiddle_factor_table_50_imag));
  assign _zz_9453 = ($signed(_zz_898) - $signed(_zz_9454));
  assign _zz_9454 = ($signed(_zz_9455) * $signed(twiddle_factor_table_50_imag));
  assign _zz_9455 = ($signed(data_mid_5_51_real) + $signed(data_mid_5_51_imag));
  assign _zz_9456 = fixTo_1074_dout;
  assign _zz_9457 = ($signed(_zz_898) + $signed(_zz_9458));
  assign _zz_9458 = ($signed(_zz_9459) * $signed(twiddle_factor_table_50_real));
  assign _zz_9459 = ($signed(data_mid_5_51_imag) - $signed(data_mid_5_51_real));
  assign _zz_9460 = fixTo_1075_dout;
  assign _zz_9461 = _zz_9462[35 : 0];
  assign _zz_9462 = _zz_9463;
  assign _zz_9463 = ($signed(_zz_9464) >>> _zz_899);
  assign _zz_9464 = _zz_9465;
  assign _zz_9465 = ($signed(_zz_9467) - $signed(_zz_896));
  assign _zz_9466 = ({9'd0,data_mid_5_19_real} <<< 9);
  assign _zz_9467 = {{9{_zz_9466[26]}}, _zz_9466};
  assign _zz_9468 = fixTo_1076_dout;
  assign _zz_9469 = _zz_9470[35 : 0];
  assign _zz_9470 = _zz_9471;
  assign _zz_9471 = ($signed(_zz_9472) >>> _zz_899);
  assign _zz_9472 = _zz_9473;
  assign _zz_9473 = ($signed(_zz_9475) - $signed(_zz_897));
  assign _zz_9474 = ({9'd0,data_mid_5_19_imag} <<< 9);
  assign _zz_9475 = {{9{_zz_9474[26]}}, _zz_9474};
  assign _zz_9476 = fixTo_1077_dout;
  assign _zz_9477 = _zz_9478[35 : 0];
  assign _zz_9478 = _zz_9479;
  assign _zz_9479 = ($signed(_zz_9480) >>> _zz_900);
  assign _zz_9480 = _zz_9481;
  assign _zz_9481 = ($signed(_zz_9483) + $signed(_zz_896));
  assign _zz_9482 = ({9'd0,data_mid_5_19_real} <<< 9);
  assign _zz_9483 = {{9{_zz_9482[26]}}, _zz_9482};
  assign _zz_9484 = fixTo_1078_dout;
  assign _zz_9485 = _zz_9486[35 : 0];
  assign _zz_9486 = _zz_9487;
  assign _zz_9487 = ($signed(_zz_9488) >>> _zz_900);
  assign _zz_9488 = _zz_9489;
  assign _zz_9489 = ($signed(_zz_9491) + $signed(_zz_897));
  assign _zz_9490 = ({9'd0,data_mid_5_19_imag} <<< 9);
  assign _zz_9491 = {{9{_zz_9490[26]}}, _zz_9490};
  assign _zz_9492 = fixTo_1079_dout;
  assign _zz_9493 = ($signed(twiddle_factor_table_51_real) + $signed(twiddle_factor_table_51_imag));
  assign _zz_9494 = ($signed(_zz_903) - $signed(_zz_9495));
  assign _zz_9495 = ($signed(_zz_9496) * $signed(twiddle_factor_table_51_imag));
  assign _zz_9496 = ($signed(data_mid_5_52_real) + $signed(data_mid_5_52_imag));
  assign _zz_9497 = fixTo_1080_dout;
  assign _zz_9498 = ($signed(_zz_903) + $signed(_zz_9499));
  assign _zz_9499 = ($signed(_zz_9500) * $signed(twiddle_factor_table_51_real));
  assign _zz_9500 = ($signed(data_mid_5_52_imag) - $signed(data_mid_5_52_real));
  assign _zz_9501 = fixTo_1081_dout;
  assign _zz_9502 = _zz_9503[35 : 0];
  assign _zz_9503 = _zz_9504;
  assign _zz_9504 = ($signed(_zz_9505) >>> _zz_904);
  assign _zz_9505 = _zz_9506;
  assign _zz_9506 = ($signed(_zz_9508) - $signed(_zz_901));
  assign _zz_9507 = ({9'd0,data_mid_5_20_real} <<< 9);
  assign _zz_9508 = {{9{_zz_9507[26]}}, _zz_9507};
  assign _zz_9509 = fixTo_1082_dout;
  assign _zz_9510 = _zz_9511[35 : 0];
  assign _zz_9511 = _zz_9512;
  assign _zz_9512 = ($signed(_zz_9513) >>> _zz_904);
  assign _zz_9513 = _zz_9514;
  assign _zz_9514 = ($signed(_zz_9516) - $signed(_zz_902));
  assign _zz_9515 = ({9'd0,data_mid_5_20_imag} <<< 9);
  assign _zz_9516 = {{9{_zz_9515[26]}}, _zz_9515};
  assign _zz_9517 = fixTo_1083_dout;
  assign _zz_9518 = _zz_9519[35 : 0];
  assign _zz_9519 = _zz_9520;
  assign _zz_9520 = ($signed(_zz_9521) >>> _zz_905);
  assign _zz_9521 = _zz_9522;
  assign _zz_9522 = ($signed(_zz_9524) + $signed(_zz_901));
  assign _zz_9523 = ({9'd0,data_mid_5_20_real} <<< 9);
  assign _zz_9524 = {{9{_zz_9523[26]}}, _zz_9523};
  assign _zz_9525 = fixTo_1084_dout;
  assign _zz_9526 = _zz_9527[35 : 0];
  assign _zz_9527 = _zz_9528;
  assign _zz_9528 = ($signed(_zz_9529) >>> _zz_905);
  assign _zz_9529 = _zz_9530;
  assign _zz_9530 = ($signed(_zz_9532) + $signed(_zz_902));
  assign _zz_9531 = ({9'd0,data_mid_5_20_imag} <<< 9);
  assign _zz_9532 = {{9{_zz_9531[26]}}, _zz_9531};
  assign _zz_9533 = fixTo_1085_dout;
  assign _zz_9534 = ($signed(twiddle_factor_table_52_real) + $signed(twiddle_factor_table_52_imag));
  assign _zz_9535 = ($signed(_zz_908) - $signed(_zz_9536));
  assign _zz_9536 = ($signed(_zz_9537) * $signed(twiddle_factor_table_52_imag));
  assign _zz_9537 = ($signed(data_mid_5_53_real) + $signed(data_mid_5_53_imag));
  assign _zz_9538 = fixTo_1086_dout;
  assign _zz_9539 = ($signed(_zz_908) + $signed(_zz_9540));
  assign _zz_9540 = ($signed(_zz_9541) * $signed(twiddle_factor_table_52_real));
  assign _zz_9541 = ($signed(data_mid_5_53_imag) - $signed(data_mid_5_53_real));
  assign _zz_9542 = fixTo_1087_dout;
  assign _zz_9543 = _zz_9544[35 : 0];
  assign _zz_9544 = _zz_9545;
  assign _zz_9545 = ($signed(_zz_9546) >>> _zz_909);
  assign _zz_9546 = _zz_9547;
  assign _zz_9547 = ($signed(_zz_9549) - $signed(_zz_906));
  assign _zz_9548 = ({9'd0,data_mid_5_21_real} <<< 9);
  assign _zz_9549 = {{9{_zz_9548[26]}}, _zz_9548};
  assign _zz_9550 = fixTo_1088_dout;
  assign _zz_9551 = _zz_9552[35 : 0];
  assign _zz_9552 = _zz_9553;
  assign _zz_9553 = ($signed(_zz_9554) >>> _zz_909);
  assign _zz_9554 = _zz_9555;
  assign _zz_9555 = ($signed(_zz_9557) - $signed(_zz_907));
  assign _zz_9556 = ({9'd0,data_mid_5_21_imag} <<< 9);
  assign _zz_9557 = {{9{_zz_9556[26]}}, _zz_9556};
  assign _zz_9558 = fixTo_1089_dout;
  assign _zz_9559 = _zz_9560[35 : 0];
  assign _zz_9560 = _zz_9561;
  assign _zz_9561 = ($signed(_zz_9562) >>> _zz_910);
  assign _zz_9562 = _zz_9563;
  assign _zz_9563 = ($signed(_zz_9565) + $signed(_zz_906));
  assign _zz_9564 = ({9'd0,data_mid_5_21_real} <<< 9);
  assign _zz_9565 = {{9{_zz_9564[26]}}, _zz_9564};
  assign _zz_9566 = fixTo_1090_dout;
  assign _zz_9567 = _zz_9568[35 : 0];
  assign _zz_9568 = _zz_9569;
  assign _zz_9569 = ($signed(_zz_9570) >>> _zz_910);
  assign _zz_9570 = _zz_9571;
  assign _zz_9571 = ($signed(_zz_9573) + $signed(_zz_907));
  assign _zz_9572 = ({9'd0,data_mid_5_21_imag} <<< 9);
  assign _zz_9573 = {{9{_zz_9572[26]}}, _zz_9572};
  assign _zz_9574 = fixTo_1091_dout;
  assign _zz_9575 = ($signed(twiddle_factor_table_53_real) + $signed(twiddle_factor_table_53_imag));
  assign _zz_9576 = ($signed(_zz_913) - $signed(_zz_9577));
  assign _zz_9577 = ($signed(_zz_9578) * $signed(twiddle_factor_table_53_imag));
  assign _zz_9578 = ($signed(data_mid_5_54_real) + $signed(data_mid_5_54_imag));
  assign _zz_9579 = fixTo_1092_dout;
  assign _zz_9580 = ($signed(_zz_913) + $signed(_zz_9581));
  assign _zz_9581 = ($signed(_zz_9582) * $signed(twiddle_factor_table_53_real));
  assign _zz_9582 = ($signed(data_mid_5_54_imag) - $signed(data_mid_5_54_real));
  assign _zz_9583 = fixTo_1093_dout;
  assign _zz_9584 = _zz_9585[35 : 0];
  assign _zz_9585 = _zz_9586;
  assign _zz_9586 = ($signed(_zz_9587) >>> _zz_914);
  assign _zz_9587 = _zz_9588;
  assign _zz_9588 = ($signed(_zz_9590) - $signed(_zz_911));
  assign _zz_9589 = ({9'd0,data_mid_5_22_real} <<< 9);
  assign _zz_9590 = {{9{_zz_9589[26]}}, _zz_9589};
  assign _zz_9591 = fixTo_1094_dout;
  assign _zz_9592 = _zz_9593[35 : 0];
  assign _zz_9593 = _zz_9594;
  assign _zz_9594 = ($signed(_zz_9595) >>> _zz_914);
  assign _zz_9595 = _zz_9596;
  assign _zz_9596 = ($signed(_zz_9598) - $signed(_zz_912));
  assign _zz_9597 = ({9'd0,data_mid_5_22_imag} <<< 9);
  assign _zz_9598 = {{9{_zz_9597[26]}}, _zz_9597};
  assign _zz_9599 = fixTo_1095_dout;
  assign _zz_9600 = _zz_9601[35 : 0];
  assign _zz_9601 = _zz_9602;
  assign _zz_9602 = ($signed(_zz_9603) >>> _zz_915);
  assign _zz_9603 = _zz_9604;
  assign _zz_9604 = ($signed(_zz_9606) + $signed(_zz_911));
  assign _zz_9605 = ({9'd0,data_mid_5_22_real} <<< 9);
  assign _zz_9606 = {{9{_zz_9605[26]}}, _zz_9605};
  assign _zz_9607 = fixTo_1096_dout;
  assign _zz_9608 = _zz_9609[35 : 0];
  assign _zz_9609 = _zz_9610;
  assign _zz_9610 = ($signed(_zz_9611) >>> _zz_915);
  assign _zz_9611 = _zz_9612;
  assign _zz_9612 = ($signed(_zz_9614) + $signed(_zz_912));
  assign _zz_9613 = ({9'd0,data_mid_5_22_imag} <<< 9);
  assign _zz_9614 = {{9{_zz_9613[26]}}, _zz_9613};
  assign _zz_9615 = fixTo_1097_dout;
  assign _zz_9616 = ($signed(twiddle_factor_table_54_real) + $signed(twiddle_factor_table_54_imag));
  assign _zz_9617 = ($signed(_zz_918) - $signed(_zz_9618));
  assign _zz_9618 = ($signed(_zz_9619) * $signed(twiddle_factor_table_54_imag));
  assign _zz_9619 = ($signed(data_mid_5_55_real) + $signed(data_mid_5_55_imag));
  assign _zz_9620 = fixTo_1098_dout;
  assign _zz_9621 = ($signed(_zz_918) + $signed(_zz_9622));
  assign _zz_9622 = ($signed(_zz_9623) * $signed(twiddle_factor_table_54_real));
  assign _zz_9623 = ($signed(data_mid_5_55_imag) - $signed(data_mid_5_55_real));
  assign _zz_9624 = fixTo_1099_dout;
  assign _zz_9625 = _zz_9626[35 : 0];
  assign _zz_9626 = _zz_9627;
  assign _zz_9627 = ($signed(_zz_9628) >>> _zz_919);
  assign _zz_9628 = _zz_9629;
  assign _zz_9629 = ($signed(_zz_9631) - $signed(_zz_916));
  assign _zz_9630 = ({9'd0,data_mid_5_23_real} <<< 9);
  assign _zz_9631 = {{9{_zz_9630[26]}}, _zz_9630};
  assign _zz_9632 = fixTo_1100_dout;
  assign _zz_9633 = _zz_9634[35 : 0];
  assign _zz_9634 = _zz_9635;
  assign _zz_9635 = ($signed(_zz_9636) >>> _zz_919);
  assign _zz_9636 = _zz_9637;
  assign _zz_9637 = ($signed(_zz_9639) - $signed(_zz_917));
  assign _zz_9638 = ({9'd0,data_mid_5_23_imag} <<< 9);
  assign _zz_9639 = {{9{_zz_9638[26]}}, _zz_9638};
  assign _zz_9640 = fixTo_1101_dout;
  assign _zz_9641 = _zz_9642[35 : 0];
  assign _zz_9642 = _zz_9643;
  assign _zz_9643 = ($signed(_zz_9644) >>> _zz_920);
  assign _zz_9644 = _zz_9645;
  assign _zz_9645 = ($signed(_zz_9647) + $signed(_zz_916));
  assign _zz_9646 = ({9'd0,data_mid_5_23_real} <<< 9);
  assign _zz_9647 = {{9{_zz_9646[26]}}, _zz_9646};
  assign _zz_9648 = fixTo_1102_dout;
  assign _zz_9649 = _zz_9650[35 : 0];
  assign _zz_9650 = _zz_9651;
  assign _zz_9651 = ($signed(_zz_9652) >>> _zz_920);
  assign _zz_9652 = _zz_9653;
  assign _zz_9653 = ($signed(_zz_9655) + $signed(_zz_917));
  assign _zz_9654 = ({9'd0,data_mid_5_23_imag} <<< 9);
  assign _zz_9655 = {{9{_zz_9654[26]}}, _zz_9654};
  assign _zz_9656 = fixTo_1103_dout;
  assign _zz_9657 = ($signed(twiddle_factor_table_55_real) + $signed(twiddle_factor_table_55_imag));
  assign _zz_9658 = ($signed(_zz_923) - $signed(_zz_9659));
  assign _zz_9659 = ($signed(_zz_9660) * $signed(twiddle_factor_table_55_imag));
  assign _zz_9660 = ($signed(data_mid_5_56_real) + $signed(data_mid_5_56_imag));
  assign _zz_9661 = fixTo_1104_dout;
  assign _zz_9662 = ($signed(_zz_923) + $signed(_zz_9663));
  assign _zz_9663 = ($signed(_zz_9664) * $signed(twiddle_factor_table_55_real));
  assign _zz_9664 = ($signed(data_mid_5_56_imag) - $signed(data_mid_5_56_real));
  assign _zz_9665 = fixTo_1105_dout;
  assign _zz_9666 = _zz_9667[35 : 0];
  assign _zz_9667 = _zz_9668;
  assign _zz_9668 = ($signed(_zz_9669) >>> _zz_924);
  assign _zz_9669 = _zz_9670;
  assign _zz_9670 = ($signed(_zz_9672) - $signed(_zz_921));
  assign _zz_9671 = ({9'd0,data_mid_5_24_real} <<< 9);
  assign _zz_9672 = {{9{_zz_9671[26]}}, _zz_9671};
  assign _zz_9673 = fixTo_1106_dout;
  assign _zz_9674 = _zz_9675[35 : 0];
  assign _zz_9675 = _zz_9676;
  assign _zz_9676 = ($signed(_zz_9677) >>> _zz_924);
  assign _zz_9677 = _zz_9678;
  assign _zz_9678 = ($signed(_zz_9680) - $signed(_zz_922));
  assign _zz_9679 = ({9'd0,data_mid_5_24_imag} <<< 9);
  assign _zz_9680 = {{9{_zz_9679[26]}}, _zz_9679};
  assign _zz_9681 = fixTo_1107_dout;
  assign _zz_9682 = _zz_9683[35 : 0];
  assign _zz_9683 = _zz_9684;
  assign _zz_9684 = ($signed(_zz_9685) >>> _zz_925);
  assign _zz_9685 = _zz_9686;
  assign _zz_9686 = ($signed(_zz_9688) + $signed(_zz_921));
  assign _zz_9687 = ({9'd0,data_mid_5_24_real} <<< 9);
  assign _zz_9688 = {{9{_zz_9687[26]}}, _zz_9687};
  assign _zz_9689 = fixTo_1108_dout;
  assign _zz_9690 = _zz_9691[35 : 0];
  assign _zz_9691 = _zz_9692;
  assign _zz_9692 = ($signed(_zz_9693) >>> _zz_925);
  assign _zz_9693 = _zz_9694;
  assign _zz_9694 = ($signed(_zz_9696) + $signed(_zz_922));
  assign _zz_9695 = ({9'd0,data_mid_5_24_imag} <<< 9);
  assign _zz_9696 = {{9{_zz_9695[26]}}, _zz_9695};
  assign _zz_9697 = fixTo_1109_dout;
  assign _zz_9698 = ($signed(twiddle_factor_table_56_real) + $signed(twiddle_factor_table_56_imag));
  assign _zz_9699 = ($signed(_zz_928) - $signed(_zz_9700));
  assign _zz_9700 = ($signed(_zz_9701) * $signed(twiddle_factor_table_56_imag));
  assign _zz_9701 = ($signed(data_mid_5_57_real) + $signed(data_mid_5_57_imag));
  assign _zz_9702 = fixTo_1110_dout;
  assign _zz_9703 = ($signed(_zz_928) + $signed(_zz_9704));
  assign _zz_9704 = ($signed(_zz_9705) * $signed(twiddle_factor_table_56_real));
  assign _zz_9705 = ($signed(data_mid_5_57_imag) - $signed(data_mid_5_57_real));
  assign _zz_9706 = fixTo_1111_dout;
  assign _zz_9707 = _zz_9708[35 : 0];
  assign _zz_9708 = _zz_9709;
  assign _zz_9709 = ($signed(_zz_9710) >>> _zz_929);
  assign _zz_9710 = _zz_9711;
  assign _zz_9711 = ($signed(_zz_9713) - $signed(_zz_926));
  assign _zz_9712 = ({9'd0,data_mid_5_25_real} <<< 9);
  assign _zz_9713 = {{9{_zz_9712[26]}}, _zz_9712};
  assign _zz_9714 = fixTo_1112_dout;
  assign _zz_9715 = _zz_9716[35 : 0];
  assign _zz_9716 = _zz_9717;
  assign _zz_9717 = ($signed(_zz_9718) >>> _zz_929);
  assign _zz_9718 = _zz_9719;
  assign _zz_9719 = ($signed(_zz_9721) - $signed(_zz_927));
  assign _zz_9720 = ({9'd0,data_mid_5_25_imag} <<< 9);
  assign _zz_9721 = {{9{_zz_9720[26]}}, _zz_9720};
  assign _zz_9722 = fixTo_1113_dout;
  assign _zz_9723 = _zz_9724[35 : 0];
  assign _zz_9724 = _zz_9725;
  assign _zz_9725 = ($signed(_zz_9726) >>> _zz_930);
  assign _zz_9726 = _zz_9727;
  assign _zz_9727 = ($signed(_zz_9729) + $signed(_zz_926));
  assign _zz_9728 = ({9'd0,data_mid_5_25_real} <<< 9);
  assign _zz_9729 = {{9{_zz_9728[26]}}, _zz_9728};
  assign _zz_9730 = fixTo_1114_dout;
  assign _zz_9731 = _zz_9732[35 : 0];
  assign _zz_9732 = _zz_9733;
  assign _zz_9733 = ($signed(_zz_9734) >>> _zz_930);
  assign _zz_9734 = _zz_9735;
  assign _zz_9735 = ($signed(_zz_9737) + $signed(_zz_927));
  assign _zz_9736 = ({9'd0,data_mid_5_25_imag} <<< 9);
  assign _zz_9737 = {{9{_zz_9736[26]}}, _zz_9736};
  assign _zz_9738 = fixTo_1115_dout;
  assign _zz_9739 = ($signed(twiddle_factor_table_57_real) + $signed(twiddle_factor_table_57_imag));
  assign _zz_9740 = ($signed(_zz_933) - $signed(_zz_9741));
  assign _zz_9741 = ($signed(_zz_9742) * $signed(twiddle_factor_table_57_imag));
  assign _zz_9742 = ($signed(data_mid_5_58_real) + $signed(data_mid_5_58_imag));
  assign _zz_9743 = fixTo_1116_dout;
  assign _zz_9744 = ($signed(_zz_933) + $signed(_zz_9745));
  assign _zz_9745 = ($signed(_zz_9746) * $signed(twiddle_factor_table_57_real));
  assign _zz_9746 = ($signed(data_mid_5_58_imag) - $signed(data_mid_5_58_real));
  assign _zz_9747 = fixTo_1117_dout;
  assign _zz_9748 = _zz_9749[35 : 0];
  assign _zz_9749 = _zz_9750;
  assign _zz_9750 = ($signed(_zz_9751) >>> _zz_934);
  assign _zz_9751 = _zz_9752;
  assign _zz_9752 = ($signed(_zz_9754) - $signed(_zz_931));
  assign _zz_9753 = ({9'd0,data_mid_5_26_real} <<< 9);
  assign _zz_9754 = {{9{_zz_9753[26]}}, _zz_9753};
  assign _zz_9755 = fixTo_1118_dout;
  assign _zz_9756 = _zz_9757[35 : 0];
  assign _zz_9757 = _zz_9758;
  assign _zz_9758 = ($signed(_zz_9759) >>> _zz_934);
  assign _zz_9759 = _zz_9760;
  assign _zz_9760 = ($signed(_zz_9762) - $signed(_zz_932));
  assign _zz_9761 = ({9'd0,data_mid_5_26_imag} <<< 9);
  assign _zz_9762 = {{9{_zz_9761[26]}}, _zz_9761};
  assign _zz_9763 = fixTo_1119_dout;
  assign _zz_9764 = _zz_9765[35 : 0];
  assign _zz_9765 = _zz_9766;
  assign _zz_9766 = ($signed(_zz_9767) >>> _zz_935);
  assign _zz_9767 = _zz_9768;
  assign _zz_9768 = ($signed(_zz_9770) + $signed(_zz_931));
  assign _zz_9769 = ({9'd0,data_mid_5_26_real} <<< 9);
  assign _zz_9770 = {{9{_zz_9769[26]}}, _zz_9769};
  assign _zz_9771 = fixTo_1120_dout;
  assign _zz_9772 = _zz_9773[35 : 0];
  assign _zz_9773 = _zz_9774;
  assign _zz_9774 = ($signed(_zz_9775) >>> _zz_935);
  assign _zz_9775 = _zz_9776;
  assign _zz_9776 = ($signed(_zz_9778) + $signed(_zz_932));
  assign _zz_9777 = ({9'd0,data_mid_5_26_imag} <<< 9);
  assign _zz_9778 = {{9{_zz_9777[26]}}, _zz_9777};
  assign _zz_9779 = fixTo_1121_dout;
  assign _zz_9780 = ($signed(twiddle_factor_table_58_real) + $signed(twiddle_factor_table_58_imag));
  assign _zz_9781 = ($signed(_zz_938) - $signed(_zz_9782));
  assign _zz_9782 = ($signed(_zz_9783) * $signed(twiddle_factor_table_58_imag));
  assign _zz_9783 = ($signed(data_mid_5_59_real) + $signed(data_mid_5_59_imag));
  assign _zz_9784 = fixTo_1122_dout;
  assign _zz_9785 = ($signed(_zz_938) + $signed(_zz_9786));
  assign _zz_9786 = ($signed(_zz_9787) * $signed(twiddle_factor_table_58_real));
  assign _zz_9787 = ($signed(data_mid_5_59_imag) - $signed(data_mid_5_59_real));
  assign _zz_9788 = fixTo_1123_dout;
  assign _zz_9789 = _zz_9790[35 : 0];
  assign _zz_9790 = _zz_9791;
  assign _zz_9791 = ($signed(_zz_9792) >>> _zz_939);
  assign _zz_9792 = _zz_9793;
  assign _zz_9793 = ($signed(_zz_9795) - $signed(_zz_936));
  assign _zz_9794 = ({9'd0,data_mid_5_27_real} <<< 9);
  assign _zz_9795 = {{9{_zz_9794[26]}}, _zz_9794};
  assign _zz_9796 = fixTo_1124_dout;
  assign _zz_9797 = _zz_9798[35 : 0];
  assign _zz_9798 = _zz_9799;
  assign _zz_9799 = ($signed(_zz_9800) >>> _zz_939);
  assign _zz_9800 = _zz_9801;
  assign _zz_9801 = ($signed(_zz_9803) - $signed(_zz_937));
  assign _zz_9802 = ({9'd0,data_mid_5_27_imag} <<< 9);
  assign _zz_9803 = {{9{_zz_9802[26]}}, _zz_9802};
  assign _zz_9804 = fixTo_1125_dout;
  assign _zz_9805 = _zz_9806[35 : 0];
  assign _zz_9806 = _zz_9807;
  assign _zz_9807 = ($signed(_zz_9808) >>> _zz_940);
  assign _zz_9808 = _zz_9809;
  assign _zz_9809 = ($signed(_zz_9811) + $signed(_zz_936));
  assign _zz_9810 = ({9'd0,data_mid_5_27_real} <<< 9);
  assign _zz_9811 = {{9{_zz_9810[26]}}, _zz_9810};
  assign _zz_9812 = fixTo_1126_dout;
  assign _zz_9813 = _zz_9814[35 : 0];
  assign _zz_9814 = _zz_9815;
  assign _zz_9815 = ($signed(_zz_9816) >>> _zz_940);
  assign _zz_9816 = _zz_9817;
  assign _zz_9817 = ($signed(_zz_9819) + $signed(_zz_937));
  assign _zz_9818 = ({9'd0,data_mid_5_27_imag} <<< 9);
  assign _zz_9819 = {{9{_zz_9818[26]}}, _zz_9818};
  assign _zz_9820 = fixTo_1127_dout;
  assign _zz_9821 = ($signed(twiddle_factor_table_59_real) + $signed(twiddle_factor_table_59_imag));
  assign _zz_9822 = ($signed(_zz_943) - $signed(_zz_9823));
  assign _zz_9823 = ($signed(_zz_9824) * $signed(twiddle_factor_table_59_imag));
  assign _zz_9824 = ($signed(data_mid_5_60_real) + $signed(data_mid_5_60_imag));
  assign _zz_9825 = fixTo_1128_dout;
  assign _zz_9826 = ($signed(_zz_943) + $signed(_zz_9827));
  assign _zz_9827 = ($signed(_zz_9828) * $signed(twiddle_factor_table_59_real));
  assign _zz_9828 = ($signed(data_mid_5_60_imag) - $signed(data_mid_5_60_real));
  assign _zz_9829 = fixTo_1129_dout;
  assign _zz_9830 = _zz_9831[35 : 0];
  assign _zz_9831 = _zz_9832;
  assign _zz_9832 = ($signed(_zz_9833) >>> _zz_944);
  assign _zz_9833 = _zz_9834;
  assign _zz_9834 = ($signed(_zz_9836) - $signed(_zz_941));
  assign _zz_9835 = ({9'd0,data_mid_5_28_real} <<< 9);
  assign _zz_9836 = {{9{_zz_9835[26]}}, _zz_9835};
  assign _zz_9837 = fixTo_1130_dout;
  assign _zz_9838 = _zz_9839[35 : 0];
  assign _zz_9839 = _zz_9840;
  assign _zz_9840 = ($signed(_zz_9841) >>> _zz_944);
  assign _zz_9841 = _zz_9842;
  assign _zz_9842 = ($signed(_zz_9844) - $signed(_zz_942));
  assign _zz_9843 = ({9'd0,data_mid_5_28_imag} <<< 9);
  assign _zz_9844 = {{9{_zz_9843[26]}}, _zz_9843};
  assign _zz_9845 = fixTo_1131_dout;
  assign _zz_9846 = _zz_9847[35 : 0];
  assign _zz_9847 = _zz_9848;
  assign _zz_9848 = ($signed(_zz_9849) >>> _zz_945);
  assign _zz_9849 = _zz_9850;
  assign _zz_9850 = ($signed(_zz_9852) + $signed(_zz_941));
  assign _zz_9851 = ({9'd0,data_mid_5_28_real} <<< 9);
  assign _zz_9852 = {{9{_zz_9851[26]}}, _zz_9851};
  assign _zz_9853 = fixTo_1132_dout;
  assign _zz_9854 = _zz_9855[35 : 0];
  assign _zz_9855 = _zz_9856;
  assign _zz_9856 = ($signed(_zz_9857) >>> _zz_945);
  assign _zz_9857 = _zz_9858;
  assign _zz_9858 = ($signed(_zz_9860) + $signed(_zz_942));
  assign _zz_9859 = ({9'd0,data_mid_5_28_imag} <<< 9);
  assign _zz_9860 = {{9{_zz_9859[26]}}, _zz_9859};
  assign _zz_9861 = fixTo_1133_dout;
  assign _zz_9862 = ($signed(twiddle_factor_table_60_real) + $signed(twiddle_factor_table_60_imag));
  assign _zz_9863 = ($signed(_zz_948) - $signed(_zz_9864));
  assign _zz_9864 = ($signed(_zz_9865) * $signed(twiddle_factor_table_60_imag));
  assign _zz_9865 = ($signed(data_mid_5_61_real) + $signed(data_mid_5_61_imag));
  assign _zz_9866 = fixTo_1134_dout;
  assign _zz_9867 = ($signed(_zz_948) + $signed(_zz_9868));
  assign _zz_9868 = ($signed(_zz_9869) * $signed(twiddle_factor_table_60_real));
  assign _zz_9869 = ($signed(data_mid_5_61_imag) - $signed(data_mid_5_61_real));
  assign _zz_9870 = fixTo_1135_dout;
  assign _zz_9871 = _zz_9872[35 : 0];
  assign _zz_9872 = _zz_9873;
  assign _zz_9873 = ($signed(_zz_9874) >>> _zz_949);
  assign _zz_9874 = _zz_9875;
  assign _zz_9875 = ($signed(_zz_9877) - $signed(_zz_946));
  assign _zz_9876 = ({9'd0,data_mid_5_29_real} <<< 9);
  assign _zz_9877 = {{9{_zz_9876[26]}}, _zz_9876};
  assign _zz_9878 = fixTo_1136_dout;
  assign _zz_9879 = _zz_9880[35 : 0];
  assign _zz_9880 = _zz_9881;
  assign _zz_9881 = ($signed(_zz_9882) >>> _zz_949);
  assign _zz_9882 = _zz_9883;
  assign _zz_9883 = ($signed(_zz_9885) - $signed(_zz_947));
  assign _zz_9884 = ({9'd0,data_mid_5_29_imag} <<< 9);
  assign _zz_9885 = {{9{_zz_9884[26]}}, _zz_9884};
  assign _zz_9886 = fixTo_1137_dout;
  assign _zz_9887 = _zz_9888[35 : 0];
  assign _zz_9888 = _zz_9889;
  assign _zz_9889 = ($signed(_zz_9890) >>> _zz_950);
  assign _zz_9890 = _zz_9891;
  assign _zz_9891 = ($signed(_zz_9893) + $signed(_zz_946));
  assign _zz_9892 = ({9'd0,data_mid_5_29_real} <<< 9);
  assign _zz_9893 = {{9{_zz_9892[26]}}, _zz_9892};
  assign _zz_9894 = fixTo_1138_dout;
  assign _zz_9895 = _zz_9896[35 : 0];
  assign _zz_9896 = _zz_9897;
  assign _zz_9897 = ($signed(_zz_9898) >>> _zz_950);
  assign _zz_9898 = _zz_9899;
  assign _zz_9899 = ($signed(_zz_9901) + $signed(_zz_947));
  assign _zz_9900 = ({9'd0,data_mid_5_29_imag} <<< 9);
  assign _zz_9901 = {{9{_zz_9900[26]}}, _zz_9900};
  assign _zz_9902 = fixTo_1139_dout;
  assign _zz_9903 = ($signed(twiddle_factor_table_61_real) + $signed(twiddle_factor_table_61_imag));
  assign _zz_9904 = ($signed(_zz_953) - $signed(_zz_9905));
  assign _zz_9905 = ($signed(_zz_9906) * $signed(twiddle_factor_table_61_imag));
  assign _zz_9906 = ($signed(data_mid_5_62_real) + $signed(data_mid_5_62_imag));
  assign _zz_9907 = fixTo_1140_dout;
  assign _zz_9908 = ($signed(_zz_953) + $signed(_zz_9909));
  assign _zz_9909 = ($signed(_zz_9910) * $signed(twiddle_factor_table_61_real));
  assign _zz_9910 = ($signed(data_mid_5_62_imag) - $signed(data_mid_5_62_real));
  assign _zz_9911 = fixTo_1141_dout;
  assign _zz_9912 = _zz_9913[35 : 0];
  assign _zz_9913 = _zz_9914;
  assign _zz_9914 = ($signed(_zz_9915) >>> _zz_954);
  assign _zz_9915 = _zz_9916;
  assign _zz_9916 = ($signed(_zz_9918) - $signed(_zz_951));
  assign _zz_9917 = ({9'd0,data_mid_5_30_real} <<< 9);
  assign _zz_9918 = {{9{_zz_9917[26]}}, _zz_9917};
  assign _zz_9919 = fixTo_1142_dout;
  assign _zz_9920 = _zz_9921[35 : 0];
  assign _zz_9921 = _zz_9922;
  assign _zz_9922 = ($signed(_zz_9923) >>> _zz_954);
  assign _zz_9923 = _zz_9924;
  assign _zz_9924 = ($signed(_zz_9926) - $signed(_zz_952));
  assign _zz_9925 = ({9'd0,data_mid_5_30_imag} <<< 9);
  assign _zz_9926 = {{9{_zz_9925[26]}}, _zz_9925};
  assign _zz_9927 = fixTo_1143_dout;
  assign _zz_9928 = _zz_9929[35 : 0];
  assign _zz_9929 = _zz_9930;
  assign _zz_9930 = ($signed(_zz_9931) >>> _zz_955);
  assign _zz_9931 = _zz_9932;
  assign _zz_9932 = ($signed(_zz_9934) + $signed(_zz_951));
  assign _zz_9933 = ({9'd0,data_mid_5_30_real} <<< 9);
  assign _zz_9934 = {{9{_zz_9933[26]}}, _zz_9933};
  assign _zz_9935 = fixTo_1144_dout;
  assign _zz_9936 = _zz_9937[35 : 0];
  assign _zz_9937 = _zz_9938;
  assign _zz_9938 = ($signed(_zz_9939) >>> _zz_955);
  assign _zz_9939 = _zz_9940;
  assign _zz_9940 = ($signed(_zz_9942) + $signed(_zz_952));
  assign _zz_9941 = ({9'd0,data_mid_5_30_imag} <<< 9);
  assign _zz_9942 = {{9{_zz_9941[26]}}, _zz_9941};
  assign _zz_9943 = fixTo_1145_dout;
  assign _zz_9944 = ($signed(twiddle_factor_table_62_real) + $signed(twiddle_factor_table_62_imag));
  assign _zz_9945 = ($signed(_zz_958) - $signed(_zz_9946));
  assign _zz_9946 = ($signed(_zz_9947) * $signed(twiddle_factor_table_62_imag));
  assign _zz_9947 = ($signed(data_mid_5_63_real) + $signed(data_mid_5_63_imag));
  assign _zz_9948 = fixTo_1146_dout;
  assign _zz_9949 = ($signed(_zz_958) + $signed(_zz_9950));
  assign _zz_9950 = ($signed(_zz_9951) * $signed(twiddle_factor_table_62_real));
  assign _zz_9951 = ($signed(data_mid_5_63_imag) - $signed(data_mid_5_63_real));
  assign _zz_9952 = fixTo_1147_dout;
  assign _zz_9953 = _zz_9954[35 : 0];
  assign _zz_9954 = _zz_9955;
  assign _zz_9955 = ($signed(_zz_9956) >>> _zz_959);
  assign _zz_9956 = _zz_9957;
  assign _zz_9957 = ($signed(_zz_9959) - $signed(_zz_956));
  assign _zz_9958 = ({9'd0,data_mid_5_31_real} <<< 9);
  assign _zz_9959 = {{9{_zz_9958[26]}}, _zz_9958};
  assign _zz_9960 = fixTo_1148_dout;
  assign _zz_9961 = _zz_9962[35 : 0];
  assign _zz_9962 = _zz_9963;
  assign _zz_9963 = ($signed(_zz_9964) >>> _zz_959);
  assign _zz_9964 = _zz_9965;
  assign _zz_9965 = ($signed(_zz_9967) - $signed(_zz_957));
  assign _zz_9966 = ({9'd0,data_mid_5_31_imag} <<< 9);
  assign _zz_9967 = {{9{_zz_9966[26]}}, _zz_9966};
  assign _zz_9968 = fixTo_1149_dout;
  assign _zz_9969 = _zz_9970[35 : 0];
  assign _zz_9970 = _zz_9971;
  assign _zz_9971 = ($signed(_zz_9972) >>> _zz_960);
  assign _zz_9972 = _zz_9973;
  assign _zz_9973 = ($signed(_zz_9975) + $signed(_zz_956));
  assign _zz_9974 = ({9'd0,data_mid_5_31_real} <<< 9);
  assign _zz_9975 = {{9{_zz_9974[26]}}, _zz_9974};
  assign _zz_9976 = fixTo_1150_dout;
  assign _zz_9977 = _zz_9978[35 : 0];
  assign _zz_9978 = _zz_9979;
  assign _zz_9979 = ($signed(_zz_9980) >>> _zz_960);
  assign _zz_9980 = _zz_9981;
  assign _zz_9981 = ($signed(_zz_9983) + $signed(_zz_957));
  assign _zz_9982 = ({9'd0,data_mid_5_31_imag} <<< 9);
  assign _zz_9983 = {{9{_zz_9982[26]}}, _zz_9982};
  assign _zz_9984 = fixTo_1151_dout;
  SInt36fixTo35_0_ROUNDTOINF fixTo (
    .din     (_zz_961[35:0]     ), //i
    .dout    (fixTo_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1 (
    .din     (_zz_962[35:0]       ), //i
    .dout    (fixTo_1_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_2 (
    .din     (_zz_963[35:0]       ), //i
    .dout    (fixTo_2_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_3 (
    .din     (_zz_964[35:0]       ), //i
    .dout    (fixTo_3_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_4 (
    .din     (_zz_965[35:0]       ), //i
    .dout    (fixTo_4_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_5 (
    .din     (_zz_966[35:0]       ), //i
    .dout    (fixTo_5_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_6 (
    .din     (_zz_967[35:0]       ), //i
    .dout    (fixTo_6_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_7 (
    .din     (_zz_968[35:0]       ), //i
    .dout    (fixTo_7_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_8 (
    .din     (_zz_969[35:0]       ), //i
    .dout    (fixTo_8_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_9 (
    .din     (_zz_970[35:0]       ), //i
    .dout    (fixTo_9_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_10 (
    .din     (_zz_971[35:0]        ), //i
    .dout    (fixTo_10_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_11 (
    .din     (_zz_972[35:0]        ), //i
    .dout    (fixTo_11_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_12 (
    .din     (_zz_973[35:0]        ), //i
    .dout    (fixTo_12_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_13 (
    .din     (_zz_974[35:0]        ), //i
    .dout    (fixTo_13_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_14 (
    .din     (_zz_975[35:0]        ), //i
    .dout    (fixTo_14_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_15 (
    .din     (_zz_976[35:0]        ), //i
    .dout    (fixTo_15_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_16 (
    .din     (_zz_977[35:0]        ), //i
    .dout    (fixTo_16_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_17 (
    .din     (_zz_978[35:0]        ), //i
    .dout    (fixTo_17_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_18 (
    .din     (_zz_979[35:0]        ), //i
    .dout    (fixTo_18_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_19 (
    .din     (_zz_980[35:0]        ), //i
    .dout    (fixTo_19_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_20 (
    .din     (_zz_981[35:0]        ), //i
    .dout    (fixTo_20_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_21 (
    .din     (_zz_982[35:0]        ), //i
    .dout    (fixTo_21_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_22 (
    .din     (_zz_983[35:0]        ), //i
    .dout    (fixTo_22_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_23 (
    .din     (_zz_984[35:0]        ), //i
    .dout    (fixTo_23_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_24 (
    .din     (_zz_985[35:0]        ), //i
    .dout    (fixTo_24_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_25 (
    .din     (_zz_986[35:0]        ), //i
    .dout    (fixTo_25_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_26 (
    .din     (_zz_987[35:0]        ), //i
    .dout    (fixTo_26_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_27 (
    .din     (_zz_988[35:0]        ), //i
    .dout    (fixTo_27_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_28 (
    .din     (_zz_989[35:0]        ), //i
    .dout    (fixTo_28_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_29 (
    .din     (_zz_990[35:0]        ), //i
    .dout    (fixTo_29_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_30 (
    .din     (_zz_991[35:0]        ), //i
    .dout    (fixTo_30_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_31 (
    .din     (_zz_992[35:0]        ), //i
    .dout    (fixTo_31_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_32 (
    .din     (_zz_993[35:0]        ), //i
    .dout    (fixTo_32_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_33 (
    .din     (_zz_994[35:0]        ), //i
    .dout    (fixTo_33_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_34 (
    .din     (_zz_995[35:0]        ), //i
    .dout    (fixTo_34_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_35 (
    .din     (_zz_996[35:0]        ), //i
    .dout    (fixTo_35_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_36 (
    .din     (_zz_997[35:0]        ), //i
    .dout    (fixTo_36_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_37 (
    .din     (_zz_998[35:0]        ), //i
    .dout    (fixTo_37_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_38 (
    .din     (_zz_999[35:0]        ), //i
    .dout    (fixTo_38_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_39 (
    .din     (_zz_1000[35:0]       ), //i
    .dout    (fixTo_39_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_40 (
    .din     (_zz_1001[35:0]       ), //i
    .dout    (fixTo_40_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_41 (
    .din     (_zz_1002[35:0]       ), //i
    .dout    (fixTo_41_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_42 (
    .din     (_zz_1003[35:0]       ), //i
    .dout    (fixTo_42_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_43 (
    .din     (_zz_1004[35:0]       ), //i
    .dout    (fixTo_43_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_44 (
    .din     (_zz_1005[35:0]       ), //i
    .dout    (fixTo_44_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_45 (
    .din     (_zz_1006[35:0]       ), //i
    .dout    (fixTo_45_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_46 (
    .din     (_zz_1007[35:0]       ), //i
    .dout    (fixTo_46_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_47 (
    .din     (_zz_1008[35:0]       ), //i
    .dout    (fixTo_47_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_48 (
    .din     (_zz_1009[35:0]       ), //i
    .dout    (fixTo_48_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_49 (
    .din     (_zz_1010[35:0]       ), //i
    .dout    (fixTo_49_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_50 (
    .din     (_zz_1011[35:0]       ), //i
    .dout    (fixTo_50_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_51 (
    .din     (_zz_1012[35:0]       ), //i
    .dout    (fixTo_51_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_52 (
    .din     (_zz_1013[35:0]       ), //i
    .dout    (fixTo_52_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_53 (
    .din     (_zz_1014[35:0]       ), //i
    .dout    (fixTo_53_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_54 (
    .din     (_zz_1015[35:0]       ), //i
    .dout    (fixTo_54_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_55 (
    .din     (_zz_1016[35:0]       ), //i
    .dout    (fixTo_55_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_56 (
    .din     (_zz_1017[35:0]       ), //i
    .dout    (fixTo_56_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_57 (
    .din     (_zz_1018[35:0]       ), //i
    .dout    (fixTo_57_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_58 (
    .din     (_zz_1019[35:0]       ), //i
    .dout    (fixTo_58_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_59 (
    .din     (_zz_1020[35:0]       ), //i
    .dout    (fixTo_59_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_60 (
    .din     (_zz_1021[35:0]       ), //i
    .dout    (fixTo_60_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_61 (
    .din     (_zz_1022[35:0]       ), //i
    .dout    (fixTo_61_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_62 (
    .din     (_zz_1023[35:0]       ), //i
    .dout    (fixTo_62_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_63 (
    .din     (_zz_1024[35:0]       ), //i
    .dout    (fixTo_63_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_64 (
    .din     (_zz_1025[35:0]       ), //i
    .dout    (fixTo_64_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_65 (
    .din     (_zz_1026[35:0]       ), //i
    .dout    (fixTo_65_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_66 (
    .din     (_zz_1027[35:0]       ), //i
    .dout    (fixTo_66_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_67 (
    .din     (_zz_1028[35:0]       ), //i
    .dout    (fixTo_67_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_68 (
    .din     (_zz_1029[35:0]       ), //i
    .dout    (fixTo_68_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_69 (
    .din     (_zz_1030[35:0]       ), //i
    .dout    (fixTo_69_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_70 (
    .din     (_zz_1031[35:0]       ), //i
    .dout    (fixTo_70_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_71 (
    .din     (_zz_1032[35:0]       ), //i
    .dout    (fixTo_71_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_72 (
    .din     (_zz_1033[35:0]       ), //i
    .dout    (fixTo_72_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_73 (
    .din     (_zz_1034[35:0]       ), //i
    .dout    (fixTo_73_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_74 (
    .din     (_zz_1035[35:0]       ), //i
    .dout    (fixTo_74_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_75 (
    .din     (_zz_1036[35:0]       ), //i
    .dout    (fixTo_75_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_76 (
    .din     (_zz_1037[35:0]       ), //i
    .dout    (fixTo_76_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_77 (
    .din     (_zz_1038[35:0]       ), //i
    .dout    (fixTo_77_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_78 (
    .din     (_zz_1039[35:0]       ), //i
    .dout    (fixTo_78_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_79 (
    .din     (_zz_1040[35:0]       ), //i
    .dout    (fixTo_79_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_80 (
    .din     (_zz_1041[35:0]       ), //i
    .dout    (fixTo_80_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_81 (
    .din     (_zz_1042[35:0]       ), //i
    .dout    (fixTo_81_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_82 (
    .din     (_zz_1043[35:0]       ), //i
    .dout    (fixTo_82_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_83 (
    .din     (_zz_1044[35:0]       ), //i
    .dout    (fixTo_83_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_84 (
    .din     (_zz_1045[35:0]       ), //i
    .dout    (fixTo_84_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_85 (
    .din     (_zz_1046[35:0]       ), //i
    .dout    (fixTo_85_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_86 (
    .din     (_zz_1047[35:0]       ), //i
    .dout    (fixTo_86_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_87 (
    .din     (_zz_1048[35:0]       ), //i
    .dout    (fixTo_87_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_88 (
    .din     (_zz_1049[35:0]       ), //i
    .dout    (fixTo_88_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_89 (
    .din     (_zz_1050[35:0]       ), //i
    .dout    (fixTo_89_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_90 (
    .din     (_zz_1051[35:0]       ), //i
    .dout    (fixTo_90_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_91 (
    .din     (_zz_1052[35:0]       ), //i
    .dout    (fixTo_91_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_92 (
    .din     (_zz_1053[35:0]       ), //i
    .dout    (fixTo_92_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_93 (
    .din     (_zz_1054[35:0]       ), //i
    .dout    (fixTo_93_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_94 (
    .din     (_zz_1055[35:0]       ), //i
    .dout    (fixTo_94_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_95 (
    .din     (_zz_1056[35:0]       ), //i
    .dout    (fixTo_95_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_96 (
    .din     (_zz_1057[35:0]       ), //i
    .dout    (fixTo_96_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_97 (
    .din     (_zz_1058[35:0]       ), //i
    .dout    (fixTo_97_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_98 (
    .din     (_zz_1059[35:0]       ), //i
    .dout    (fixTo_98_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_99 (
    .din     (_zz_1060[35:0]       ), //i
    .dout    (fixTo_99_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_100 (
    .din     (_zz_1061[35:0]        ), //i
    .dout    (fixTo_100_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_101 (
    .din     (_zz_1062[35:0]        ), //i
    .dout    (fixTo_101_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_102 (
    .din     (_zz_1063[35:0]        ), //i
    .dout    (fixTo_102_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_103 (
    .din     (_zz_1064[35:0]        ), //i
    .dout    (fixTo_103_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_104 (
    .din     (_zz_1065[35:0]        ), //i
    .dout    (fixTo_104_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_105 (
    .din     (_zz_1066[35:0]        ), //i
    .dout    (fixTo_105_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_106 (
    .din     (_zz_1067[35:0]        ), //i
    .dout    (fixTo_106_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_107 (
    .din     (_zz_1068[35:0]        ), //i
    .dout    (fixTo_107_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_108 (
    .din     (_zz_1069[35:0]        ), //i
    .dout    (fixTo_108_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_109 (
    .din     (_zz_1070[35:0]        ), //i
    .dout    (fixTo_109_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_110 (
    .din     (_zz_1071[35:0]        ), //i
    .dout    (fixTo_110_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_111 (
    .din     (_zz_1072[35:0]        ), //i
    .dout    (fixTo_111_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_112 (
    .din     (_zz_1073[35:0]        ), //i
    .dout    (fixTo_112_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_113 (
    .din     (_zz_1074[35:0]        ), //i
    .dout    (fixTo_113_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_114 (
    .din     (_zz_1075[35:0]        ), //i
    .dout    (fixTo_114_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_115 (
    .din     (_zz_1076[35:0]        ), //i
    .dout    (fixTo_115_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_116 (
    .din     (_zz_1077[35:0]        ), //i
    .dout    (fixTo_116_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_117 (
    .din     (_zz_1078[35:0]        ), //i
    .dout    (fixTo_117_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_118 (
    .din     (_zz_1079[35:0]        ), //i
    .dout    (fixTo_118_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_119 (
    .din     (_zz_1080[35:0]        ), //i
    .dout    (fixTo_119_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_120 (
    .din     (_zz_1081[35:0]        ), //i
    .dout    (fixTo_120_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_121 (
    .din     (_zz_1082[35:0]        ), //i
    .dout    (fixTo_121_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_122 (
    .din     (_zz_1083[35:0]        ), //i
    .dout    (fixTo_122_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_123 (
    .din     (_zz_1084[35:0]        ), //i
    .dout    (fixTo_123_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_124 (
    .din     (_zz_1085[35:0]        ), //i
    .dout    (fixTo_124_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_125 (
    .din     (_zz_1086[35:0]        ), //i
    .dout    (fixTo_125_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_126 (
    .din     (_zz_1087[35:0]        ), //i
    .dout    (fixTo_126_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_127 (
    .din     (_zz_1088[35:0]        ), //i
    .dout    (fixTo_127_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_128 (
    .din     (_zz_1089[35:0]        ), //i
    .dout    (fixTo_128_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_129 (
    .din     (_zz_1090[35:0]        ), //i
    .dout    (fixTo_129_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_130 (
    .din     (_zz_1091[35:0]        ), //i
    .dout    (fixTo_130_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_131 (
    .din     (_zz_1092[35:0]        ), //i
    .dout    (fixTo_131_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_132 (
    .din     (_zz_1093[35:0]        ), //i
    .dout    (fixTo_132_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_133 (
    .din     (_zz_1094[35:0]        ), //i
    .dout    (fixTo_133_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_134 (
    .din     (_zz_1095[35:0]        ), //i
    .dout    (fixTo_134_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_135 (
    .din     (_zz_1096[35:0]        ), //i
    .dout    (fixTo_135_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_136 (
    .din     (_zz_1097[35:0]        ), //i
    .dout    (fixTo_136_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_137 (
    .din     (_zz_1098[35:0]        ), //i
    .dout    (fixTo_137_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_138 (
    .din     (_zz_1099[35:0]        ), //i
    .dout    (fixTo_138_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_139 (
    .din     (_zz_1100[35:0]        ), //i
    .dout    (fixTo_139_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_140 (
    .din     (_zz_1101[35:0]        ), //i
    .dout    (fixTo_140_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_141 (
    .din     (_zz_1102[35:0]        ), //i
    .dout    (fixTo_141_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_142 (
    .din     (_zz_1103[35:0]        ), //i
    .dout    (fixTo_142_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_143 (
    .din     (_zz_1104[35:0]        ), //i
    .dout    (fixTo_143_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_144 (
    .din     (_zz_1105[35:0]        ), //i
    .dout    (fixTo_144_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_145 (
    .din     (_zz_1106[35:0]        ), //i
    .dout    (fixTo_145_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_146 (
    .din     (_zz_1107[35:0]        ), //i
    .dout    (fixTo_146_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_147 (
    .din     (_zz_1108[35:0]        ), //i
    .dout    (fixTo_147_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_148 (
    .din     (_zz_1109[35:0]        ), //i
    .dout    (fixTo_148_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_149 (
    .din     (_zz_1110[35:0]        ), //i
    .dout    (fixTo_149_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_150 (
    .din     (_zz_1111[35:0]        ), //i
    .dout    (fixTo_150_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_151 (
    .din     (_zz_1112[35:0]        ), //i
    .dout    (fixTo_151_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_152 (
    .din     (_zz_1113[35:0]        ), //i
    .dout    (fixTo_152_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_153 (
    .din     (_zz_1114[35:0]        ), //i
    .dout    (fixTo_153_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_154 (
    .din     (_zz_1115[35:0]        ), //i
    .dout    (fixTo_154_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_155 (
    .din     (_zz_1116[35:0]        ), //i
    .dout    (fixTo_155_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_156 (
    .din     (_zz_1117[35:0]        ), //i
    .dout    (fixTo_156_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_157 (
    .din     (_zz_1118[35:0]        ), //i
    .dout    (fixTo_157_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_158 (
    .din     (_zz_1119[35:0]        ), //i
    .dout    (fixTo_158_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_159 (
    .din     (_zz_1120[35:0]        ), //i
    .dout    (fixTo_159_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_160 (
    .din     (_zz_1121[35:0]        ), //i
    .dout    (fixTo_160_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_161 (
    .din     (_zz_1122[35:0]        ), //i
    .dout    (fixTo_161_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_162 (
    .din     (_zz_1123[35:0]        ), //i
    .dout    (fixTo_162_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_163 (
    .din     (_zz_1124[35:0]        ), //i
    .dout    (fixTo_163_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_164 (
    .din     (_zz_1125[35:0]        ), //i
    .dout    (fixTo_164_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_165 (
    .din     (_zz_1126[35:0]        ), //i
    .dout    (fixTo_165_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_166 (
    .din     (_zz_1127[35:0]        ), //i
    .dout    (fixTo_166_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_167 (
    .din     (_zz_1128[35:0]        ), //i
    .dout    (fixTo_167_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_168 (
    .din     (_zz_1129[35:0]        ), //i
    .dout    (fixTo_168_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_169 (
    .din     (_zz_1130[35:0]        ), //i
    .dout    (fixTo_169_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_170 (
    .din     (_zz_1131[35:0]        ), //i
    .dout    (fixTo_170_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_171 (
    .din     (_zz_1132[35:0]        ), //i
    .dout    (fixTo_171_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_172 (
    .din     (_zz_1133[35:0]        ), //i
    .dout    (fixTo_172_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_173 (
    .din     (_zz_1134[35:0]        ), //i
    .dout    (fixTo_173_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_174 (
    .din     (_zz_1135[35:0]        ), //i
    .dout    (fixTo_174_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_175 (
    .din     (_zz_1136[35:0]        ), //i
    .dout    (fixTo_175_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_176 (
    .din     (_zz_1137[35:0]        ), //i
    .dout    (fixTo_176_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_177 (
    .din     (_zz_1138[35:0]        ), //i
    .dout    (fixTo_177_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_178 (
    .din     (_zz_1139[35:0]        ), //i
    .dout    (fixTo_178_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_179 (
    .din     (_zz_1140[35:0]        ), //i
    .dout    (fixTo_179_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_180 (
    .din     (_zz_1141[35:0]        ), //i
    .dout    (fixTo_180_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_181 (
    .din     (_zz_1142[35:0]        ), //i
    .dout    (fixTo_181_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_182 (
    .din     (_zz_1143[35:0]        ), //i
    .dout    (fixTo_182_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_183 (
    .din     (_zz_1144[35:0]        ), //i
    .dout    (fixTo_183_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_184 (
    .din     (_zz_1145[35:0]        ), //i
    .dout    (fixTo_184_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_185 (
    .din     (_zz_1146[35:0]        ), //i
    .dout    (fixTo_185_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_186 (
    .din     (_zz_1147[35:0]        ), //i
    .dout    (fixTo_186_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_187 (
    .din     (_zz_1148[35:0]        ), //i
    .dout    (fixTo_187_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_188 (
    .din     (_zz_1149[35:0]        ), //i
    .dout    (fixTo_188_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_189 (
    .din     (_zz_1150[35:0]        ), //i
    .dout    (fixTo_189_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_190 (
    .din     (_zz_1151[35:0]        ), //i
    .dout    (fixTo_190_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_191 (
    .din     (_zz_1152[35:0]        ), //i
    .dout    (fixTo_191_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_192 (
    .din     (_zz_1153[35:0]        ), //i
    .dout    (fixTo_192_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_193 (
    .din     (_zz_1154[35:0]        ), //i
    .dout    (fixTo_193_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_194 (
    .din     (_zz_1155[35:0]        ), //i
    .dout    (fixTo_194_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_195 (
    .din     (_zz_1156[35:0]        ), //i
    .dout    (fixTo_195_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_196 (
    .din     (_zz_1157[35:0]        ), //i
    .dout    (fixTo_196_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_197 (
    .din     (_zz_1158[35:0]        ), //i
    .dout    (fixTo_197_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_198 (
    .din     (_zz_1159[35:0]        ), //i
    .dout    (fixTo_198_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_199 (
    .din     (_zz_1160[35:0]        ), //i
    .dout    (fixTo_199_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_200 (
    .din     (_zz_1161[35:0]        ), //i
    .dout    (fixTo_200_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_201 (
    .din     (_zz_1162[35:0]        ), //i
    .dout    (fixTo_201_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_202 (
    .din     (_zz_1163[35:0]        ), //i
    .dout    (fixTo_202_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_203 (
    .din     (_zz_1164[35:0]        ), //i
    .dout    (fixTo_203_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_204 (
    .din     (_zz_1165[35:0]        ), //i
    .dout    (fixTo_204_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_205 (
    .din     (_zz_1166[35:0]        ), //i
    .dout    (fixTo_205_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_206 (
    .din     (_zz_1167[35:0]        ), //i
    .dout    (fixTo_206_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_207 (
    .din     (_zz_1168[35:0]        ), //i
    .dout    (fixTo_207_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_208 (
    .din     (_zz_1169[35:0]        ), //i
    .dout    (fixTo_208_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_209 (
    .din     (_zz_1170[35:0]        ), //i
    .dout    (fixTo_209_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_210 (
    .din     (_zz_1171[35:0]        ), //i
    .dout    (fixTo_210_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_211 (
    .din     (_zz_1172[35:0]        ), //i
    .dout    (fixTo_211_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_212 (
    .din     (_zz_1173[35:0]        ), //i
    .dout    (fixTo_212_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_213 (
    .din     (_zz_1174[35:0]        ), //i
    .dout    (fixTo_213_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_214 (
    .din     (_zz_1175[35:0]        ), //i
    .dout    (fixTo_214_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_215 (
    .din     (_zz_1176[35:0]        ), //i
    .dout    (fixTo_215_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_216 (
    .din     (_zz_1177[35:0]        ), //i
    .dout    (fixTo_216_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_217 (
    .din     (_zz_1178[35:0]        ), //i
    .dout    (fixTo_217_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_218 (
    .din     (_zz_1179[35:0]        ), //i
    .dout    (fixTo_218_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_219 (
    .din     (_zz_1180[35:0]        ), //i
    .dout    (fixTo_219_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_220 (
    .din     (_zz_1181[35:0]        ), //i
    .dout    (fixTo_220_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_221 (
    .din     (_zz_1182[35:0]        ), //i
    .dout    (fixTo_221_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_222 (
    .din     (_zz_1183[35:0]        ), //i
    .dout    (fixTo_222_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_223 (
    .din     (_zz_1184[35:0]        ), //i
    .dout    (fixTo_223_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_224 (
    .din     (_zz_1185[35:0]        ), //i
    .dout    (fixTo_224_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_225 (
    .din     (_zz_1186[35:0]        ), //i
    .dout    (fixTo_225_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_226 (
    .din     (_zz_1187[35:0]        ), //i
    .dout    (fixTo_226_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_227 (
    .din     (_zz_1188[35:0]        ), //i
    .dout    (fixTo_227_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_228 (
    .din     (_zz_1189[35:0]        ), //i
    .dout    (fixTo_228_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_229 (
    .din     (_zz_1190[35:0]        ), //i
    .dout    (fixTo_229_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_230 (
    .din     (_zz_1191[35:0]        ), //i
    .dout    (fixTo_230_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_231 (
    .din     (_zz_1192[35:0]        ), //i
    .dout    (fixTo_231_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_232 (
    .din     (_zz_1193[35:0]        ), //i
    .dout    (fixTo_232_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_233 (
    .din     (_zz_1194[35:0]        ), //i
    .dout    (fixTo_233_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_234 (
    .din     (_zz_1195[35:0]        ), //i
    .dout    (fixTo_234_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_235 (
    .din     (_zz_1196[35:0]        ), //i
    .dout    (fixTo_235_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_236 (
    .din     (_zz_1197[35:0]        ), //i
    .dout    (fixTo_236_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_237 (
    .din     (_zz_1198[35:0]        ), //i
    .dout    (fixTo_237_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_238 (
    .din     (_zz_1199[35:0]        ), //i
    .dout    (fixTo_238_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_239 (
    .din     (_zz_1200[35:0]        ), //i
    .dout    (fixTo_239_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_240 (
    .din     (_zz_1201[35:0]        ), //i
    .dout    (fixTo_240_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_241 (
    .din     (_zz_1202[35:0]        ), //i
    .dout    (fixTo_241_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_242 (
    .din     (_zz_1203[35:0]        ), //i
    .dout    (fixTo_242_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_243 (
    .din     (_zz_1204[35:0]        ), //i
    .dout    (fixTo_243_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_244 (
    .din     (_zz_1205[35:0]        ), //i
    .dout    (fixTo_244_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_245 (
    .din     (_zz_1206[35:0]        ), //i
    .dout    (fixTo_245_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_246 (
    .din     (_zz_1207[35:0]        ), //i
    .dout    (fixTo_246_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_247 (
    .din     (_zz_1208[35:0]        ), //i
    .dout    (fixTo_247_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_248 (
    .din     (_zz_1209[35:0]        ), //i
    .dout    (fixTo_248_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_249 (
    .din     (_zz_1210[35:0]        ), //i
    .dout    (fixTo_249_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_250 (
    .din     (_zz_1211[35:0]        ), //i
    .dout    (fixTo_250_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_251 (
    .din     (_zz_1212[35:0]        ), //i
    .dout    (fixTo_251_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_252 (
    .din     (_zz_1213[35:0]        ), //i
    .dout    (fixTo_252_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_253 (
    .din     (_zz_1214[35:0]        ), //i
    .dout    (fixTo_253_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_254 (
    .din     (_zz_1215[35:0]        ), //i
    .dout    (fixTo_254_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_255 (
    .din     (_zz_1216[35:0]        ), //i
    .dout    (fixTo_255_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_256 (
    .din     (_zz_1217[35:0]        ), //i
    .dout    (fixTo_256_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_257 (
    .din     (_zz_1218[35:0]        ), //i
    .dout    (fixTo_257_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_258 (
    .din     (_zz_1219[35:0]        ), //i
    .dout    (fixTo_258_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_259 (
    .din     (_zz_1220[35:0]        ), //i
    .dout    (fixTo_259_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_260 (
    .din     (_zz_1221[35:0]        ), //i
    .dout    (fixTo_260_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_261 (
    .din     (_zz_1222[35:0]        ), //i
    .dout    (fixTo_261_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_262 (
    .din     (_zz_1223[35:0]        ), //i
    .dout    (fixTo_262_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_263 (
    .din     (_zz_1224[35:0]        ), //i
    .dout    (fixTo_263_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_264 (
    .din     (_zz_1225[35:0]        ), //i
    .dout    (fixTo_264_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_265 (
    .din     (_zz_1226[35:0]        ), //i
    .dout    (fixTo_265_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_266 (
    .din     (_zz_1227[35:0]        ), //i
    .dout    (fixTo_266_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_267 (
    .din     (_zz_1228[35:0]        ), //i
    .dout    (fixTo_267_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_268 (
    .din     (_zz_1229[35:0]        ), //i
    .dout    (fixTo_268_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_269 (
    .din     (_zz_1230[35:0]        ), //i
    .dout    (fixTo_269_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_270 (
    .din     (_zz_1231[35:0]        ), //i
    .dout    (fixTo_270_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_271 (
    .din     (_zz_1232[35:0]        ), //i
    .dout    (fixTo_271_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_272 (
    .din     (_zz_1233[35:0]        ), //i
    .dout    (fixTo_272_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_273 (
    .din     (_zz_1234[35:0]        ), //i
    .dout    (fixTo_273_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_274 (
    .din     (_zz_1235[35:0]        ), //i
    .dout    (fixTo_274_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_275 (
    .din     (_zz_1236[35:0]        ), //i
    .dout    (fixTo_275_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_276 (
    .din     (_zz_1237[35:0]        ), //i
    .dout    (fixTo_276_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_277 (
    .din     (_zz_1238[35:0]        ), //i
    .dout    (fixTo_277_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_278 (
    .din     (_zz_1239[35:0]        ), //i
    .dout    (fixTo_278_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_279 (
    .din     (_zz_1240[35:0]        ), //i
    .dout    (fixTo_279_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_280 (
    .din     (_zz_1241[35:0]        ), //i
    .dout    (fixTo_280_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_281 (
    .din     (_zz_1242[35:0]        ), //i
    .dout    (fixTo_281_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_282 (
    .din     (_zz_1243[35:0]        ), //i
    .dout    (fixTo_282_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_283 (
    .din     (_zz_1244[35:0]        ), //i
    .dout    (fixTo_283_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_284 (
    .din     (_zz_1245[35:0]        ), //i
    .dout    (fixTo_284_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_285 (
    .din     (_zz_1246[35:0]        ), //i
    .dout    (fixTo_285_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_286 (
    .din     (_zz_1247[35:0]        ), //i
    .dout    (fixTo_286_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_287 (
    .din     (_zz_1248[35:0]        ), //i
    .dout    (fixTo_287_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_288 (
    .din     (_zz_1249[35:0]        ), //i
    .dout    (fixTo_288_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_289 (
    .din     (_zz_1250[35:0]        ), //i
    .dout    (fixTo_289_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_290 (
    .din     (_zz_1251[35:0]        ), //i
    .dout    (fixTo_290_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_291 (
    .din     (_zz_1252[35:0]        ), //i
    .dout    (fixTo_291_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_292 (
    .din     (_zz_1253[35:0]        ), //i
    .dout    (fixTo_292_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_293 (
    .din     (_zz_1254[35:0]        ), //i
    .dout    (fixTo_293_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_294 (
    .din     (_zz_1255[35:0]        ), //i
    .dout    (fixTo_294_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_295 (
    .din     (_zz_1256[35:0]        ), //i
    .dout    (fixTo_295_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_296 (
    .din     (_zz_1257[35:0]        ), //i
    .dout    (fixTo_296_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_297 (
    .din     (_zz_1258[35:0]        ), //i
    .dout    (fixTo_297_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_298 (
    .din     (_zz_1259[35:0]        ), //i
    .dout    (fixTo_298_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_299 (
    .din     (_zz_1260[35:0]        ), //i
    .dout    (fixTo_299_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_300 (
    .din     (_zz_1261[35:0]        ), //i
    .dout    (fixTo_300_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_301 (
    .din     (_zz_1262[35:0]        ), //i
    .dout    (fixTo_301_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_302 (
    .din     (_zz_1263[35:0]        ), //i
    .dout    (fixTo_302_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_303 (
    .din     (_zz_1264[35:0]        ), //i
    .dout    (fixTo_303_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_304 (
    .din     (_zz_1265[35:0]        ), //i
    .dout    (fixTo_304_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_305 (
    .din     (_zz_1266[35:0]        ), //i
    .dout    (fixTo_305_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_306 (
    .din     (_zz_1267[35:0]        ), //i
    .dout    (fixTo_306_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_307 (
    .din     (_zz_1268[35:0]        ), //i
    .dout    (fixTo_307_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_308 (
    .din     (_zz_1269[35:0]        ), //i
    .dout    (fixTo_308_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_309 (
    .din     (_zz_1270[35:0]        ), //i
    .dout    (fixTo_309_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_310 (
    .din     (_zz_1271[35:0]        ), //i
    .dout    (fixTo_310_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_311 (
    .din     (_zz_1272[35:0]        ), //i
    .dout    (fixTo_311_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_312 (
    .din     (_zz_1273[35:0]        ), //i
    .dout    (fixTo_312_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_313 (
    .din     (_zz_1274[35:0]        ), //i
    .dout    (fixTo_313_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_314 (
    .din     (_zz_1275[35:0]        ), //i
    .dout    (fixTo_314_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_315 (
    .din     (_zz_1276[35:0]        ), //i
    .dout    (fixTo_315_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_316 (
    .din     (_zz_1277[35:0]        ), //i
    .dout    (fixTo_316_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_317 (
    .din     (_zz_1278[35:0]        ), //i
    .dout    (fixTo_317_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_318 (
    .din     (_zz_1279[35:0]        ), //i
    .dout    (fixTo_318_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_319 (
    .din     (_zz_1280[35:0]        ), //i
    .dout    (fixTo_319_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_320 (
    .din     (_zz_1281[35:0]        ), //i
    .dout    (fixTo_320_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_321 (
    .din     (_zz_1282[35:0]        ), //i
    .dout    (fixTo_321_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_322 (
    .din     (_zz_1283[35:0]        ), //i
    .dout    (fixTo_322_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_323 (
    .din     (_zz_1284[35:0]        ), //i
    .dout    (fixTo_323_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_324 (
    .din     (_zz_1285[35:0]        ), //i
    .dout    (fixTo_324_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_325 (
    .din     (_zz_1286[35:0]        ), //i
    .dout    (fixTo_325_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_326 (
    .din     (_zz_1287[35:0]        ), //i
    .dout    (fixTo_326_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_327 (
    .din     (_zz_1288[35:0]        ), //i
    .dout    (fixTo_327_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_328 (
    .din     (_zz_1289[35:0]        ), //i
    .dout    (fixTo_328_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_329 (
    .din     (_zz_1290[35:0]        ), //i
    .dout    (fixTo_329_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_330 (
    .din     (_zz_1291[35:0]        ), //i
    .dout    (fixTo_330_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_331 (
    .din     (_zz_1292[35:0]        ), //i
    .dout    (fixTo_331_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_332 (
    .din     (_zz_1293[35:0]        ), //i
    .dout    (fixTo_332_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_333 (
    .din     (_zz_1294[35:0]        ), //i
    .dout    (fixTo_333_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_334 (
    .din     (_zz_1295[35:0]        ), //i
    .dout    (fixTo_334_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_335 (
    .din     (_zz_1296[35:0]        ), //i
    .dout    (fixTo_335_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_336 (
    .din     (_zz_1297[35:0]        ), //i
    .dout    (fixTo_336_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_337 (
    .din     (_zz_1298[35:0]        ), //i
    .dout    (fixTo_337_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_338 (
    .din     (_zz_1299[35:0]        ), //i
    .dout    (fixTo_338_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_339 (
    .din     (_zz_1300[35:0]        ), //i
    .dout    (fixTo_339_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_340 (
    .din     (_zz_1301[35:0]        ), //i
    .dout    (fixTo_340_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_341 (
    .din     (_zz_1302[35:0]        ), //i
    .dout    (fixTo_341_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_342 (
    .din     (_zz_1303[35:0]        ), //i
    .dout    (fixTo_342_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_343 (
    .din     (_zz_1304[35:0]        ), //i
    .dout    (fixTo_343_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_344 (
    .din     (_zz_1305[35:0]        ), //i
    .dout    (fixTo_344_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_345 (
    .din     (_zz_1306[35:0]        ), //i
    .dout    (fixTo_345_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_346 (
    .din     (_zz_1307[35:0]        ), //i
    .dout    (fixTo_346_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_347 (
    .din     (_zz_1308[35:0]        ), //i
    .dout    (fixTo_347_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_348 (
    .din     (_zz_1309[35:0]        ), //i
    .dout    (fixTo_348_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_349 (
    .din     (_zz_1310[35:0]        ), //i
    .dout    (fixTo_349_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_350 (
    .din     (_zz_1311[35:0]        ), //i
    .dout    (fixTo_350_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_351 (
    .din     (_zz_1312[35:0]        ), //i
    .dout    (fixTo_351_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_352 (
    .din     (_zz_1313[35:0]        ), //i
    .dout    (fixTo_352_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_353 (
    .din     (_zz_1314[35:0]        ), //i
    .dout    (fixTo_353_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_354 (
    .din     (_zz_1315[35:0]        ), //i
    .dout    (fixTo_354_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_355 (
    .din     (_zz_1316[35:0]        ), //i
    .dout    (fixTo_355_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_356 (
    .din     (_zz_1317[35:0]        ), //i
    .dout    (fixTo_356_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_357 (
    .din     (_zz_1318[35:0]        ), //i
    .dout    (fixTo_357_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_358 (
    .din     (_zz_1319[35:0]        ), //i
    .dout    (fixTo_358_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_359 (
    .din     (_zz_1320[35:0]        ), //i
    .dout    (fixTo_359_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_360 (
    .din     (_zz_1321[35:0]        ), //i
    .dout    (fixTo_360_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_361 (
    .din     (_zz_1322[35:0]        ), //i
    .dout    (fixTo_361_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_362 (
    .din     (_zz_1323[35:0]        ), //i
    .dout    (fixTo_362_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_363 (
    .din     (_zz_1324[35:0]        ), //i
    .dout    (fixTo_363_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_364 (
    .din     (_zz_1325[35:0]        ), //i
    .dout    (fixTo_364_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_365 (
    .din     (_zz_1326[35:0]        ), //i
    .dout    (fixTo_365_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_366 (
    .din     (_zz_1327[35:0]        ), //i
    .dout    (fixTo_366_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_367 (
    .din     (_zz_1328[35:0]        ), //i
    .dout    (fixTo_367_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_368 (
    .din     (_zz_1329[35:0]        ), //i
    .dout    (fixTo_368_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_369 (
    .din     (_zz_1330[35:0]        ), //i
    .dout    (fixTo_369_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_370 (
    .din     (_zz_1331[35:0]        ), //i
    .dout    (fixTo_370_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_371 (
    .din     (_zz_1332[35:0]        ), //i
    .dout    (fixTo_371_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_372 (
    .din     (_zz_1333[35:0]        ), //i
    .dout    (fixTo_372_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_373 (
    .din     (_zz_1334[35:0]        ), //i
    .dout    (fixTo_373_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_374 (
    .din     (_zz_1335[35:0]        ), //i
    .dout    (fixTo_374_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_375 (
    .din     (_zz_1336[35:0]        ), //i
    .dout    (fixTo_375_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_376 (
    .din     (_zz_1337[35:0]        ), //i
    .dout    (fixTo_376_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_377 (
    .din     (_zz_1338[35:0]        ), //i
    .dout    (fixTo_377_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_378 (
    .din     (_zz_1339[35:0]        ), //i
    .dout    (fixTo_378_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_379 (
    .din     (_zz_1340[35:0]        ), //i
    .dout    (fixTo_379_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_380 (
    .din     (_zz_1341[35:0]        ), //i
    .dout    (fixTo_380_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_381 (
    .din     (_zz_1342[35:0]        ), //i
    .dout    (fixTo_381_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_382 (
    .din     (_zz_1343[35:0]        ), //i
    .dout    (fixTo_382_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_383 (
    .din     (_zz_1344[35:0]        ), //i
    .dout    (fixTo_383_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_384 (
    .din     (_zz_1345[35:0]        ), //i
    .dout    (fixTo_384_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_385 (
    .din     (_zz_1346[35:0]        ), //i
    .dout    (fixTo_385_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_386 (
    .din     (_zz_1347[35:0]        ), //i
    .dout    (fixTo_386_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_387 (
    .din     (_zz_1348[35:0]        ), //i
    .dout    (fixTo_387_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_388 (
    .din     (_zz_1349[35:0]        ), //i
    .dout    (fixTo_388_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_389 (
    .din     (_zz_1350[35:0]        ), //i
    .dout    (fixTo_389_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_390 (
    .din     (_zz_1351[35:0]        ), //i
    .dout    (fixTo_390_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_391 (
    .din     (_zz_1352[35:0]        ), //i
    .dout    (fixTo_391_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_392 (
    .din     (_zz_1353[35:0]        ), //i
    .dout    (fixTo_392_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_393 (
    .din     (_zz_1354[35:0]        ), //i
    .dout    (fixTo_393_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_394 (
    .din     (_zz_1355[35:0]        ), //i
    .dout    (fixTo_394_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_395 (
    .din     (_zz_1356[35:0]        ), //i
    .dout    (fixTo_395_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_396 (
    .din     (_zz_1357[35:0]        ), //i
    .dout    (fixTo_396_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_397 (
    .din     (_zz_1358[35:0]        ), //i
    .dout    (fixTo_397_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_398 (
    .din     (_zz_1359[35:0]        ), //i
    .dout    (fixTo_398_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_399 (
    .din     (_zz_1360[35:0]        ), //i
    .dout    (fixTo_399_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_400 (
    .din     (_zz_1361[35:0]        ), //i
    .dout    (fixTo_400_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_401 (
    .din     (_zz_1362[35:0]        ), //i
    .dout    (fixTo_401_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_402 (
    .din     (_zz_1363[35:0]        ), //i
    .dout    (fixTo_402_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_403 (
    .din     (_zz_1364[35:0]        ), //i
    .dout    (fixTo_403_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_404 (
    .din     (_zz_1365[35:0]        ), //i
    .dout    (fixTo_404_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_405 (
    .din     (_zz_1366[35:0]        ), //i
    .dout    (fixTo_405_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_406 (
    .din     (_zz_1367[35:0]        ), //i
    .dout    (fixTo_406_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_407 (
    .din     (_zz_1368[35:0]        ), //i
    .dout    (fixTo_407_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_408 (
    .din     (_zz_1369[35:0]        ), //i
    .dout    (fixTo_408_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_409 (
    .din     (_zz_1370[35:0]        ), //i
    .dout    (fixTo_409_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_410 (
    .din     (_zz_1371[35:0]        ), //i
    .dout    (fixTo_410_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_411 (
    .din     (_zz_1372[35:0]        ), //i
    .dout    (fixTo_411_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_412 (
    .din     (_zz_1373[35:0]        ), //i
    .dout    (fixTo_412_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_413 (
    .din     (_zz_1374[35:0]        ), //i
    .dout    (fixTo_413_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_414 (
    .din     (_zz_1375[35:0]        ), //i
    .dout    (fixTo_414_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_415 (
    .din     (_zz_1376[35:0]        ), //i
    .dout    (fixTo_415_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_416 (
    .din     (_zz_1377[35:0]        ), //i
    .dout    (fixTo_416_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_417 (
    .din     (_zz_1378[35:0]        ), //i
    .dout    (fixTo_417_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_418 (
    .din     (_zz_1379[35:0]        ), //i
    .dout    (fixTo_418_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_419 (
    .din     (_zz_1380[35:0]        ), //i
    .dout    (fixTo_419_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_420 (
    .din     (_zz_1381[35:0]        ), //i
    .dout    (fixTo_420_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_421 (
    .din     (_zz_1382[35:0]        ), //i
    .dout    (fixTo_421_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_422 (
    .din     (_zz_1383[35:0]        ), //i
    .dout    (fixTo_422_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_423 (
    .din     (_zz_1384[35:0]        ), //i
    .dout    (fixTo_423_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_424 (
    .din     (_zz_1385[35:0]        ), //i
    .dout    (fixTo_424_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_425 (
    .din     (_zz_1386[35:0]        ), //i
    .dout    (fixTo_425_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_426 (
    .din     (_zz_1387[35:0]        ), //i
    .dout    (fixTo_426_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_427 (
    .din     (_zz_1388[35:0]        ), //i
    .dout    (fixTo_427_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_428 (
    .din     (_zz_1389[35:0]        ), //i
    .dout    (fixTo_428_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_429 (
    .din     (_zz_1390[35:0]        ), //i
    .dout    (fixTo_429_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_430 (
    .din     (_zz_1391[35:0]        ), //i
    .dout    (fixTo_430_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_431 (
    .din     (_zz_1392[35:0]        ), //i
    .dout    (fixTo_431_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_432 (
    .din     (_zz_1393[35:0]        ), //i
    .dout    (fixTo_432_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_433 (
    .din     (_zz_1394[35:0]        ), //i
    .dout    (fixTo_433_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_434 (
    .din     (_zz_1395[35:0]        ), //i
    .dout    (fixTo_434_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_435 (
    .din     (_zz_1396[35:0]        ), //i
    .dout    (fixTo_435_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_436 (
    .din     (_zz_1397[35:0]        ), //i
    .dout    (fixTo_436_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_437 (
    .din     (_zz_1398[35:0]        ), //i
    .dout    (fixTo_437_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_438 (
    .din     (_zz_1399[35:0]        ), //i
    .dout    (fixTo_438_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_439 (
    .din     (_zz_1400[35:0]        ), //i
    .dout    (fixTo_439_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_440 (
    .din     (_zz_1401[35:0]        ), //i
    .dout    (fixTo_440_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_441 (
    .din     (_zz_1402[35:0]        ), //i
    .dout    (fixTo_441_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_442 (
    .din     (_zz_1403[35:0]        ), //i
    .dout    (fixTo_442_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_443 (
    .din     (_zz_1404[35:0]        ), //i
    .dout    (fixTo_443_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_444 (
    .din     (_zz_1405[35:0]        ), //i
    .dout    (fixTo_444_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_445 (
    .din     (_zz_1406[35:0]        ), //i
    .dout    (fixTo_445_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_446 (
    .din     (_zz_1407[35:0]        ), //i
    .dout    (fixTo_446_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_447 (
    .din     (_zz_1408[35:0]        ), //i
    .dout    (fixTo_447_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_448 (
    .din     (_zz_1409[35:0]        ), //i
    .dout    (fixTo_448_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_449 (
    .din     (_zz_1410[35:0]        ), //i
    .dout    (fixTo_449_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_450 (
    .din     (_zz_1411[35:0]        ), //i
    .dout    (fixTo_450_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_451 (
    .din     (_zz_1412[35:0]        ), //i
    .dout    (fixTo_451_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_452 (
    .din     (_zz_1413[35:0]        ), //i
    .dout    (fixTo_452_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_453 (
    .din     (_zz_1414[35:0]        ), //i
    .dout    (fixTo_453_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_454 (
    .din     (_zz_1415[35:0]        ), //i
    .dout    (fixTo_454_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_455 (
    .din     (_zz_1416[35:0]        ), //i
    .dout    (fixTo_455_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_456 (
    .din     (_zz_1417[35:0]        ), //i
    .dout    (fixTo_456_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_457 (
    .din     (_zz_1418[35:0]        ), //i
    .dout    (fixTo_457_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_458 (
    .din     (_zz_1419[35:0]        ), //i
    .dout    (fixTo_458_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_459 (
    .din     (_zz_1420[35:0]        ), //i
    .dout    (fixTo_459_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_460 (
    .din     (_zz_1421[35:0]        ), //i
    .dout    (fixTo_460_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_461 (
    .din     (_zz_1422[35:0]        ), //i
    .dout    (fixTo_461_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_462 (
    .din     (_zz_1423[35:0]        ), //i
    .dout    (fixTo_462_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_463 (
    .din     (_zz_1424[35:0]        ), //i
    .dout    (fixTo_463_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_464 (
    .din     (_zz_1425[35:0]        ), //i
    .dout    (fixTo_464_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_465 (
    .din     (_zz_1426[35:0]        ), //i
    .dout    (fixTo_465_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_466 (
    .din     (_zz_1427[35:0]        ), //i
    .dout    (fixTo_466_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_467 (
    .din     (_zz_1428[35:0]        ), //i
    .dout    (fixTo_467_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_468 (
    .din     (_zz_1429[35:0]        ), //i
    .dout    (fixTo_468_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_469 (
    .din     (_zz_1430[35:0]        ), //i
    .dout    (fixTo_469_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_470 (
    .din     (_zz_1431[35:0]        ), //i
    .dout    (fixTo_470_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_471 (
    .din     (_zz_1432[35:0]        ), //i
    .dout    (fixTo_471_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_472 (
    .din     (_zz_1433[35:0]        ), //i
    .dout    (fixTo_472_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_473 (
    .din     (_zz_1434[35:0]        ), //i
    .dout    (fixTo_473_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_474 (
    .din     (_zz_1435[35:0]        ), //i
    .dout    (fixTo_474_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_475 (
    .din     (_zz_1436[35:0]        ), //i
    .dout    (fixTo_475_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_476 (
    .din     (_zz_1437[35:0]        ), //i
    .dout    (fixTo_476_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_477 (
    .din     (_zz_1438[35:0]        ), //i
    .dout    (fixTo_477_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_478 (
    .din     (_zz_1439[35:0]        ), //i
    .dout    (fixTo_478_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_479 (
    .din     (_zz_1440[35:0]        ), //i
    .dout    (fixTo_479_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_480 (
    .din     (_zz_1441[35:0]        ), //i
    .dout    (fixTo_480_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_481 (
    .din     (_zz_1442[35:0]        ), //i
    .dout    (fixTo_481_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_482 (
    .din     (_zz_1443[35:0]        ), //i
    .dout    (fixTo_482_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_483 (
    .din     (_zz_1444[35:0]        ), //i
    .dout    (fixTo_483_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_484 (
    .din     (_zz_1445[35:0]        ), //i
    .dout    (fixTo_484_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_485 (
    .din     (_zz_1446[35:0]        ), //i
    .dout    (fixTo_485_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_486 (
    .din     (_zz_1447[35:0]        ), //i
    .dout    (fixTo_486_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_487 (
    .din     (_zz_1448[35:0]        ), //i
    .dout    (fixTo_487_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_488 (
    .din     (_zz_1449[35:0]        ), //i
    .dout    (fixTo_488_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_489 (
    .din     (_zz_1450[35:0]        ), //i
    .dout    (fixTo_489_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_490 (
    .din     (_zz_1451[35:0]        ), //i
    .dout    (fixTo_490_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_491 (
    .din     (_zz_1452[35:0]        ), //i
    .dout    (fixTo_491_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_492 (
    .din     (_zz_1453[35:0]        ), //i
    .dout    (fixTo_492_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_493 (
    .din     (_zz_1454[35:0]        ), //i
    .dout    (fixTo_493_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_494 (
    .din     (_zz_1455[35:0]        ), //i
    .dout    (fixTo_494_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_495 (
    .din     (_zz_1456[35:0]        ), //i
    .dout    (fixTo_495_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_496 (
    .din     (_zz_1457[35:0]        ), //i
    .dout    (fixTo_496_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_497 (
    .din     (_zz_1458[35:0]        ), //i
    .dout    (fixTo_497_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_498 (
    .din     (_zz_1459[35:0]        ), //i
    .dout    (fixTo_498_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_499 (
    .din     (_zz_1460[35:0]        ), //i
    .dout    (fixTo_499_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_500 (
    .din     (_zz_1461[35:0]        ), //i
    .dout    (fixTo_500_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_501 (
    .din     (_zz_1462[35:0]        ), //i
    .dout    (fixTo_501_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_502 (
    .din     (_zz_1463[35:0]        ), //i
    .dout    (fixTo_502_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_503 (
    .din     (_zz_1464[35:0]        ), //i
    .dout    (fixTo_503_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_504 (
    .din     (_zz_1465[35:0]        ), //i
    .dout    (fixTo_504_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_505 (
    .din     (_zz_1466[35:0]        ), //i
    .dout    (fixTo_505_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_506 (
    .din     (_zz_1467[35:0]        ), //i
    .dout    (fixTo_506_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_507 (
    .din     (_zz_1468[35:0]        ), //i
    .dout    (fixTo_507_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_508 (
    .din     (_zz_1469[35:0]        ), //i
    .dout    (fixTo_508_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_509 (
    .din     (_zz_1470[35:0]        ), //i
    .dout    (fixTo_509_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_510 (
    .din     (_zz_1471[35:0]        ), //i
    .dout    (fixTo_510_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_511 (
    .din     (_zz_1472[35:0]        ), //i
    .dout    (fixTo_511_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_512 (
    .din     (_zz_1473[35:0]        ), //i
    .dout    (fixTo_512_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_513 (
    .din     (_zz_1474[35:0]        ), //i
    .dout    (fixTo_513_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_514 (
    .din     (_zz_1475[35:0]        ), //i
    .dout    (fixTo_514_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_515 (
    .din     (_zz_1476[35:0]        ), //i
    .dout    (fixTo_515_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_516 (
    .din     (_zz_1477[35:0]        ), //i
    .dout    (fixTo_516_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_517 (
    .din     (_zz_1478[35:0]        ), //i
    .dout    (fixTo_517_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_518 (
    .din     (_zz_1479[35:0]        ), //i
    .dout    (fixTo_518_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_519 (
    .din     (_zz_1480[35:0]        ), //i
    .dout    (fixTo_519_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_520 (
    .din     (_zz_1481[35:0]        ), //i
    .dout    (fixTo_520_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_521 (
    .din     (_zz_1482[35:0]        ), //i
    .dout    (fixTo_521_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_522 (
    .din     (_zz_1483[35:0]        ), //i
    .dout    (fixTo_522_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_523 (
    .din     (_zz_1484[35:0]        ), //i
    .dout    (fixTo_523_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_524 (
    .din     (_zz_1485[35:0]        ), //i
    .dout    (fixTo_524_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_525 (
    .din     (_zz_1486[35:0]        ), //i
    .dout    (fixTo_525_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_526 (
    .din     (_zz_1487[35:0]        ), //i
    .dout    (fixTo_526_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_527 (
    .din     (_zz_1488[35:0]        ), //i
    .dout    (fixTo_527_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_528 (
    .din     (_zz_1489[35:0]        ), //i
    .dout    (fixTo_528_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_529 (
    .din     (_zz_1490[35:0]        ), //i
    .dout    (fixTo_529_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_530 (
    .din     (_zz_1491[35:0]        ), //i
    .dout    (fixTo_530_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_531 (
    .din     (_zz_1492[35:0]        ), //i
    .dout    (fixTo_531_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_532 (
    .din     (_zz_1493[35:0]        ), //i
    .dout    (fixTo_532_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_533 (
    .din     (_zz_1494[35:0]        ), //i
    .dout    (fixTo_533_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_534 (
    .din     (_zz_1495[35:0]        ), //i
    .dout    (fixTo_534_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_535 (
    .din     (_zz_1496[35:0]        ), //i
    .dout    (fixTo_535_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_536 (
    .din     (_zz_1497[35:0]        ), //i
    .dout    (fixTo_536_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_537 (
    .din     (_zz_1498[35:0]        ), //i
    .dout    (fixTo_537_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_538 (
    .din     (_zz_1499[35:0]        ), //i
    .dout    (fixTo_538_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_539 (
    .din     (_zz_1500[35:0]        ), //i
    .dout    (fixTo_539_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_540 (
    .din     (_zz_1501[35:0]        ), //i
    .dout    (fixTo_540_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_541 (
    .din     (_zz_1502[35:0]        ), //i
    .dout    (fixTo_541_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_542 (
    .din     (_zz_1503[35:0]        ), //i
    .dout    (fixTo_542_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_543 (
    .din     (_zz_1504[35:0]        ), //i
    .dout    (fixTo_543_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_544 (
    .din     (_zz_1505[35:0]        ), //i
    .dout    (fixTo_544_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_545 (
    .din     (_zz_1506[35:0]        ), //i
    .dout    (fixTo_545_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_546 (
    .din     (_zz_1507[35:0]        ), //i
    .dout    (fixTo_546_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_547 (
    .din     (_zz_1508[35:0]        ), //i
    .dout    (fixTo_547_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_548 (
    .din     (_zz_1509[35:0]        ), //i
    .dout    (fixTo_548_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_549 (
    .din     (_zz_1510[35:0]        ), //i
    .dout    (fixTo_549_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_550 (
    .din     (_zz_1511[35:0]        ), //i
    .dout    (fixTo_550_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_551 (
    .din     (_zz_1512[35:0]        ), //i
    .dout    (fixTo_551_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_552 (
    .din     (_zz_1513[35:0]        ), //i
    .dout    (fixTo_552_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_553 (
    .din     (_zz_1514[35:0]        ), //i
    .dout    (fixTo_553_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_554 (
    .din     (_zz_1515[35:0]        ), //i
    .dout    (fixTo_554_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_555 (
    .din     (_zz_1516[35:0]        ), //i
    .dout    (fixTo_555_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_556 (
    .din     (_zz_1517[35:0]        ), //i
    .dout    (fixTo_556_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_557 (
    .din     (_zz_1518[35:0]        ), //i
    .dout    (fixTo_557_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_558 (
    .din     (_zz_1519[35:0]        ), //i
    .dout    (fixTo_558_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_559 (
    .din     (_zz_1520[35:0]        ), //i
    .dout    (fixTo_559_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_560 (
    .din     (_zz_1521[35:0]        ), //i
    .dout    (fixTo_560_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_561 (
    .din     (_zz_1522[35:0]        ), //i
    .dout    (fixTo_561_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_562 (
    .din     (_zz_1523[35:0]        ), //i
    .dout    (fixTo_562_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_563 (
    .din     (_zz_1524[35:0]        ), //i
    .dout    (fixTo_563_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_564 (
    .din     (_zz_1525[35:0]        ), //i
    .dout    (fixTo_564_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_565 (
    .din     (_zz_1526[35:0]        ), //i
    .dout    (fixTo_565_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_566 (
    .din     (_zz_1527[35:0]        ), //i
    .dout    (fixTo_566_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_567 (
    .din     (_zz_1528[35:0]        ), //i
    .dout    (fixTo_567_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_568 (
    .din     (_zz_1529[35:0]        ), //i
    .dout    (fixTo_568_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_569 (
    .din     (_zz_1530[35:0]        ), //i
    .dout    (fixTo_569_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_570 (
    .din     (_zz_1531[35:0]        ), //i
    .dout    (fixTo_570_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_571 (
    .din     (_zz_1532[35:0]        ), //i
    .dout    (fixTo_571_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_572 (
    .din     (_zz_1533[35:0]        ), //i
    .dout    (fixTo_572_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_573 (
    .din     (_zz_1534[35:0]        ), //i
    .dout    (fixTo_573_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_574 (
    .din     (_zz_1535[35:0]        ), //i
    .dout    (fixTo_574_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_575 (
    .din     (_zz_1536[35:0]        ), //i
    .dout    (fixTo_575_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_576 (
    .din     (_zz_1537[35:0]        ), //i
    .dout    (fixTo_576_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_577 (
    .din     (_zz_1538[35:0]        ), //i
    .dout    (fixTo_577_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_578 (
    .din     (_zz_1539[35:0]        ), //i
    .dout    (fixTo_578_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_579 (
    .din     (_zz_1540[35:0]        ), //i
    .dout    (fixTo_579_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_580 (
    .din     (_zz_1541[35:0]        ), //i
    .dout    (fixTo_580_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_581 (
    .din     (_zz_1542[35:0]        ), //i
    .dout    (fixTo_581_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_582 (
    .din     (_zz_1543[35:0]        ), //i
    .dout    (fixTo_582_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_583 (
    .din     (_zz_1544[35:0]        ), //i
    .dout    (fixTo_583_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_584 (
    .din     (_zz_1545[35:0]        ), //i
    .dout    (fixTo_584_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_585 (
    .din     (_zz_1546[35:0]        ), //i
    .dout    (fixTo_585_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_586 (
    .din     (_zz_1547[35:0]        ), //i
    .dout    (fixTo_586_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_587 (
    .din     (_zz_1548[35:0]        ), //i
    .dout    (fixTo_587_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_588 (
    .din     (_zz_1549[35:0]        ), //i
    .dout    (fixTo_588_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_589 (
    .din     (_zz_1550[35:0]        ), //i
    .dout    (fixTo_589_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_590 (
    .din     (_zz_1551[35:0]        ), //i
    .dout    (fixTo_590_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_591 (
    .din     (_zz_1552[35:0]        ), //i
    .dout    (fixTo_591_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_592 (
    .din     (_zz_1553[35:0]        ), //i
    .dout    (fixTo_592_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_593 (
    .din     (_zz_1554[35:0]        ), //i
    .dout    (fixTo_593_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_594 (
    .din     (_zz_1555[35:0]        ), //i
    .dout    (fixTo_594_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_595 (
    .din     (_zz_1556[35:0]        ), //i
    .dout    (fixTo_595_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_596 (
    .din     (_zz_1557[35:0]        ), //i
    .dout    (fixTo_596_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_597 (
    .din     (_zz_1558[35:0]        ), //i
    .dout    (fixTo_597_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_598 (
    .din     (_zz_1559[35:0]        ), //i
    .dout    (fixTo_598_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_599 (
    .din     (_zz_1560[35:0]        ), //i
    .dout    (fixTo_599_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_600 (
    .din     (_zz_1561[35:0]        ), //i
    .dout    (fixTo_600_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_601 (
    .din     (_zz_1562[35:0]        ), //i
    .dout    (fixTo_601_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_602 (
    .din     (_zz_1563[35:0]        ), //i
    .dout    (fixTo_602_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_603 (
    .din     (_zz_1564[35:0]        ), //i
    .dout    (fixTo_603_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_604 (
    .din     (_zz_1565[35:0]        ), //i
    .dout    (fixTo_604_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_605 (
    .din     (_zz_1566[35:0]        ), //i
    .dout    (fixTo_605_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_606 (
    .din     (_zz_1567[35:0]        ), //i
    .dout    (fixTo_606_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_607 (
    .din     (_zz_1568[35:0]        ), //i
    .dout    (fixTo_607_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_608 (
    .din     (_zz_1569[35:0]        ), //i
    .dout    (fixTo_608_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_609 (
    .din     (_zz_1570[35:0]        ), //i
    .dout    (fixTo_609_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_610 (
    .din     (_zz_1571[35:0]        ), //i
    .dout    (fixTo_610_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_611 (
    .din     (_zz_1572[35:0]        ), //i
    .dout    (fixTo_611_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_612 (
    .din     (_zz_1573[35:0]        ), //i
    .dout    (fixTo_612_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_613 (
    .din     (_zz_1574[35:0]        ), //i
    .dout    (fixTo_613_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_614 (
    .din     (_zz_1575[35:0]        ), //i
    .dout    (fixTo_614_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_615 (
    .din     (_zz_1576[35:0]        ), //i
    .dout    (fixTo_615_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_616 (
    .din     (_zz_1577[35:0]        ), //i
    .dout    (fixTo_616_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_617 (
    .din     (_zz_1578[35:0]        ), //i
    .dout    (fixTo_617_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_618 (
    .din     (_zz_1579[35:0]        ), //i
    .dout    (fixTo_618_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_619 (
    .din     (_zz_1580[35:0]        ), //i
    .dout    (fixTo_619_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_620 (
    .din     (_zz_1581[35:0]        ), //i
    .dout    (fixTo_620_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_621 (
    .din     (_zz_1582[35:0]        ), //i
    .dout    (fixTo_621_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_622 (
    .din     (_zz_1583[35:0]        ), //i
    .dout    (fixTo_622_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_623 (
    .din     (_zz_1584[35:0]        ), //i
    .dout    (fixTo_623_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_624 (
    .din     (_zz_1585[35:0]        ), //i
    .dout    (fixTo_624_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_625 (
    .din     (_zz_1586[35:0]        ), //i
    .dout    (fixTo_625_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_626 (
    .din     (_zz_1587[35:0]        ), //i
    .dout    (fixTo_626_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_627 (
    .din     (_zz_1588[35:0]        ), //i
    .dout    (fixTo_627_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_628 (
    .din     (_zz_1589[35:0]        ), //i
    .dout    (fixTo_628_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_629 (
    .din     (_zz_1590[35:0]        ), //i
    .dout    (fixTo_629_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_630 (
    .din     (_zz_1591[35:0]        ), //i
    .dout    (fixTo_630_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_631 (
    .din     (_zz_1592[35:0]        ), //i
    .dout    (fixTo_631_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_632 (
    .din     (_zz_1593[35:0]        ), //i
    .dout    (fixTo_632_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_633 (
    .din     (_zz_1594[35:0]        ), //i
    .dout    (fixTo_633_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_634 (
    .din     (_zz_1595[35:0]        ), //i
    .dout    (fixTo_634_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_635 (
    .din     (_zz_1596[35:0]        ), //i
    .dout    (fixTo_635_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_636 (
    .din     (_zz_1597[35:0]        ), //i
    .dout    (fixTo_636_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_637 (
    .din     (_zz_1598[35:0]        ), //i
    .dout    (fixTo_637_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_638 (
    .din     (_zz_1599[35:0]        ), //i
    .dout    (fixTo_638_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_639 (
    .din     (_zz_1600[35:0]        ), //i
    .dout    (fixTo_639_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_640 (
    .din     (_zz_1601[35:0]        ), //i
    .dout    (fixTo_640_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_641 (
    .din     (_zz_1602[35:0]        ), //i
    .dout    (fixTo_641_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_642 (
    .din     (_zz_1603[35:0]        ), //i
    .dout    (fixTo_642_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_643 (
    .din     (_zz_1604[35:0]        ), //i
    .dout    (fixTo_643_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_644 (
    .din     (_zz_1605[35:0]        ), //i
    .dout    (fixTo_644_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_645 (
    .din     (_zz_1606[35:0]        ), //i
    .dout    (fixTo_645_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_646 (
    .din     (_zz_1607[35:0]        ), //i
    .dout    (fixTo_646_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_647 (
    .din     (_zz_1608[35:0]        ), //i
    .dout    (fixTo_647_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_648 (
    .din     (_zz_1609[35:0]        ), //i
    .dout    (fixTo_648_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_649 (
    .din     (_zz_1610[35:0]        ), //i
    .dout    (fixTo_649_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_650 (
    .din     (_zz_1611[35:0]        ), //i
    .dout    (fixTo_650_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_651 (
    .din     (_zz_1612[35:0]        ), //i
    .dout    (fixTo_651_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_652 (
    .din     (_zz_1613[35:0]        ), //i
    .dout    (fixTo_652_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_653 (
    .din     (_zz_1614[35:0]        ), //i
    .dout    (fixTo_653_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_654 (
    .din     (_zz_1615[35:0]        ), //i
    .dout    (fixTo_654_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_655 (
    .din     (_zz_1616[35:0]        ), //i
    .dout    (fixTo_655_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_656 (
    .din     (_zz_1617[35:0]        ), //i
    .dout    (fixTo_656_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_657 (
    .din     (_zz_1618[35:0]        ), //i
    .dout    (fixTo_657_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_658 (
    .din     (_zz_1619[35:0]        ), //i
    .dout    (fixTo_658_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_659 (
    .din     (_zz_1620[35:0]        ), //i
    .dout    (fixTo_659_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_660 (
    .din     (_zz_1621[35:0]        ), //i
    .dout    (fixTo_660_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_661 (
    .din     (_zz_1622[35:0]        ), //i
    .dout    (fixTo_661_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_662 (
    .din     (_zz_1623[35:0]        ), //i
    .dout    (fixTo_662_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_663 (
    .din     (_zz_1624[35:0]        ), //i
    .dout    (fixTo_663_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_664 (
    .din     (_zz_1625[35:0]        ), //i
    .dout    (fixTo_664_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_665 (
    .din     (_zz_1626[35:0]        ), //i
    .dout    (fixTo_665_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_666 (
    .din     (_zz_1627[35:0]        ), //i
    .dout    (fixTo_666_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_667 (
    .din     (_zz_1628[35:0]        ), //i
    .dout    (fixTo_667_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_668 (
    .din     (_zz_1629[35:0]        ), //i
    .dout    (fixTo_668_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_669 (
    .din     (_zz_1630[35:0]        ), //i
    .dout    (fixTo_669_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_670 (
    .din     (_zz_1631[35:0]        ), //i
    .dout    (fixTo_670_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_671 (
    .din     (_zz_1632[35:0]        ), //i
    .dout    (fixTo_671_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_672 (
    .din     (_zz_1633[35:0]        ), //i
    .dout    (fixTo_672_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_673 (
    .din     (_zz_1634[35:0]        ), //i
    .dout    (fixTo_673_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_674 (
    .din     (_zz_1635[35:0]        ), //i
    .dout    (fixTo_674_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_675 (
    .din     (_zz_1636[35:0]        ), //i
    .dout    (fixTo_675_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_676 (
    .din     (_zz_1637[35:0]        ), //i
    .dout    (fixTo_676_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_677 (
    .din     (_zz_1638[35:0]        ), //i
    .dout    (fixTo_677_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_678 (
    .din     (_zz_1639[35:0]        ), //i
    .dout    (fixTo_678_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_679 (
    .din     (_zz_1640[35:0]        ), //i
    .dout    (fixTo_679_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_680 (
    .din     (_zz_1641[35:0]        ), //i
    .dout    (fixTo_680_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_681 (
    .din     (_zz_1642[35:0]        ), //i
    .dout    (fixTo_681_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_682 (
    .din     (_zz_1643[35:0]        ), //i
    .dout    (fixTo_682_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_683 (
    .din     (_zz_1644[35:0]        ), //i
    .dout    (fixTo_683_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_684 (
    .din     (_zz_1645[35:0]        ), //i
    .dout    (fixTo_684_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_685 (
    .din     (_zz_1646[35:0]        ), //i
    .dout    (fixTo_685_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_686 (
    .din     (_zz_1647[35:0]        ), //i
    .dout    (fixTo_686_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_687 (
    .din     (_zz_1648[35:0]        ), //i
    .dout    (fixTo_687_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_688 (
    .din     (_zz_1649[35:0]        ), //i
    .dout    (fixTo_688_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_689 (
    .din     (_zz_1650[35:0]        ), //i
    .dout    (fixTo_689_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_690 (
    .din     (_zz_1651[35:0]        ), //i
    .dout    (fixTo_690_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_691 (
    .din     (_zz_1652[35:0]        ), //i
    .dout    (fixTo_691_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_692 (
    .din     (_zz_1653[35:0]        ), //i
    .dout    (fixTo_692_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_693 (
    .din     (_zz_1654[35:0]        ), //i
    .dout    (fixTo_693_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_694 (
    .din     (_zz_1655[35:0]        ), //i
    .dout    (fixTo_694_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_695 (
    .din     (_zz_1656[35:0]        ), //i
    .dout    (fixTo_695_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_696 (
    .din     (_zz_1657[35:0]        ), //i
    .dout    (fixTo_696_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_697 (
    .din     (_zz_1658[35:0]        ), //i
    .dout    (fixTo_697_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_698 (
    .din     (_zz_1659[35:0]        ), //i
    .dout    (fixTo_698_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_699 (
    .din     (_zz_1660[35:0]        ), //i
    .dout    (fixTo_699_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_700 (
    .din     (_zz_1661[35:0]        ), //i
    .dout    (fixTo_700_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_701 (
    .din     (_zz_1662[35:0]        ), //i
    .dout    (fixTo_701_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_702 (
    .din     (_zz_1663[35:0]        ), //i
    .dout    (fixTo_702_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_703 (
    .din     (_zz_1664[35:0]        ), //i
    .dout    (fixTo_703_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_704 (
    .din     (_zz_1665[35:0]        ), //i
    .dout    (fixTo_704_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_705 (
    .din     (_zz_1666[35:0]        ), //i
    .dout    (fixTo_705_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_706 (
    .din     (_zz_1667[35:0]        ), //i
    .dout    (fixTo_706_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_707 (
    .din     (_zz_1668[35:0]        ), //i
    .dout    (fixTo_707_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_708 (
    .din     (_zz_1669[35:0]        ), //i
    .dout    (fixTo_708_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_709 (
    .din     (_zz_1670[35:0]        ), //i
    .dout    (fixTo_709_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_710 (
    .din     (_zz_1671[35:0]        ), //i
    .dout    (fixTo_710_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_711 (
    .din     (_zz_1672[35:0]        ), //i
    .dout    (fixTo_711_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_712 (
    .din     (_zz_1673[35:0]        ), //i
    .dout    (fixTo_712_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_713 (
    .din     (_zz_1674[35:0]        ), //i
    .dout    (fixTo_713_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_714 (
    .din     (_zz_1675[35:0]        ), //i
    .dout    (fixTo_714_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_715 (
    .din     (_zz_1676[35:0]        ), //i
    .dout    (fixTo_715_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_716 (
    .din     (_zz_1677[35:0]        ), //i
    .dout    (fixTo_716_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_717 (
    .din     (_zz_1678[35:0]        ), //i
    .dout    (fixTo_717_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_718 (
    .din     (_zz_1679[35:0]        ), //i
    .dout    (fixTo_718_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_719 (
    .din     (_zz_1680[35:0]        ), //i
    .dout    (fixTo_719_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_720 (
    .din     (_zz_1681[35:0]        ), //i
    .dout    (fixTo_720_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_721 (
    .din     (_zz_1682[35:0]        ), //i
    .dout    (fixTo_721_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_722 (
    .din     (_zz_1683[35:0]        ), //i
    .dout    (fixTo_722_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_723 (
    .din     (_zz_1684[35:0]        ), //i
    .dout    (fixTo_723_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_724 (
    .din     (_zz_1685[35:0]        ), //i
    .dout    (fixTo_724_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_725 (
    .din     (_zz_1686[35:0]        ), //i
    .dout    (fixTo_725_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_726 (
    .din     (_zz_1687[35:0]        ), //i
    .dout    (fixTo_726_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_727 (
    .din     (_zz_1688[35:0]        ), //i
    .dout    (fixTo_727_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_728 (
    .din     (_zz_1689[35:0]        ), //i
    .dout    (fixTo_728_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_729 (
    .din     (_zz_1690[35:0]        ), //i
    .dout    (fixTo_729_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_730 (
    .din     (_zz_1691[35:0]        ), //i
    .dout    (fixTo_730_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_731 (
    .din     (_zz_1692[35:0]        ), //i
    .dout    (fixTo_731_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_732 (
    .din     (_zz_1693[35:0]        ), //i
    .dout    (fixTo_732_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_733 (
    .din     (_zz_1694[35:0]        ), //i
    .dout    (fixTo_733_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_734 (
    .din     (_zz_1695[35:0]        ), //i
    .dout    (fixTo_734_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_735 (
    .din     (_zz_1696[35:0]        ), //i
    .dout    (fixTo_735_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_736 (
    .din     (_zz_1697[35:0]        ), //i
    .dout    (fixTo_736_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_737 (
    .din     (_zz_1698[35:0]        ), //i
    .dout    (fixTo_737_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_738 (
    .din     (_zz_1699[35:0]        ), //i
    .dout    (fixTo_738_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_739 (
    .din     (_zz_1700[35:0]        ), //i
    .dout    (fixTo_739_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_740 (
    .din     (_zz_1701[35:0]        ), //i
    .dout    (fixTo_740_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_741 (
    .din     (_zz_1702[35:0]        ), //i
    .dout    (fixTo_741_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_742 (
    .din     (_zz_1703[35:0]        ), //i
    .dout    (fixTo_742_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_743 (
    .din     (_zz_1704[35:0]        ), //i
    .dout    (fixTo_743_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_744 (
    .din     (_zz_1705[35:0]        ), //i
    .dout    (fixTo_744_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_745 (
    .din     (_zz_1706[35:0]        ), //i
    .dout    (fixTo_745_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_746 (
    .din     (_zz_1707[35:0]        ), //i
    .dout    (fixTo_746_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_747 (
    .din     (_zz_1708[35:0]        ), //i
    .dout    (fixTo_747_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_748 (
    .din     (_zz_1709[35:0]        ), //i
    .dout    (fixTo_748_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_749 (
    .din     (_zz_1710[35:0]        ), //i
    .dout    (fixTo_749_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_750 (
    .din     (_zz_1711[35:0]        ), //i
    .dout    (fixTo_750_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_751 (
    .din     (_zz_1712[35:0]        ), //i
    .dout    (fixTo_751_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_752 (
    .din     (_zz_1713[35:0]        ), //i
    .dout    (fixTo_752_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_753 (
    .din     (_zz_1714[35:0]        ), //i
    .dout    (fixTo_753_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_754 (
    .din     (_zz_1715[35:0]        ), //i
    .dout    (fixTo_754_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_755 (
    .din     (_zz_1716[35:0]        ), //i
    .dout    (fixTo_755_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_756 (
    .din     (_zz_1717[35:0]        ), //i
    .dout    (fixTo_756_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_757 (
    .din     (_zz_1718[35:0]        ), //i
    .dout    (fixTo_757_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_758 (
    .din     (_zz_1719[35:0]        ), //i
    .dout    (fixTo_758_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_759 (
    .din     (_zz_1720[35:0]        ), //i
    .dout    (fixTo_759_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_760 (
    .din     (_zz_1721[35:0]        ), //i
    .dout    (fixTo_760_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_761 (
    .din     (_zz_1722[35:0]        ), //i
    .dout    (fixTo_761_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_762 (
    .din     (_zz_1723[35:0]        ), //i
    .dout    (fixTo_762_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_763 (
    .din     (_zz_1724[35:0]        ), //i
    .dout    (fixTo_763_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_764 (
    .din     (_zz_1725[35:0]        ), //i
    .dout    (fixTo_764_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_765 (
    .din     (_zz_1726[35:0]        ), //i
    .dout    (fixTo_765_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_766 (
    .din     (_zz_1727[35:0]        ), //i
    .dout    (fixTo_766_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_767 (
    .din     (_zz_1728[35:0]        ), //i
    .dout    (fixTo_767_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_768 (
    .din     (_zz_1729[35:0]        ), //i
    .dout    (fixTo_768_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_769 (
    .din     (_zz_1730[35:0]        ), //i
    .dout    (fixTo_769_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_770 (
    .din     (_zz_1731[35:0]        ), //i
    .dout    (fixTo_770_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_771 (
    .din     (_zz_1732[35:0]        ), //i
    .dout    (fixTo_771_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_772 (
    .din     (_zz_1733[35:0]        ), //i
    .dout    (fixTo_772_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_773 (
    .din     (_zz_1734[35:0]        ), //i
    .dout    (fixTo_773_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_774 (
    .din     (_zz_1735[35:0]        ), //i
    .dout    (fixTo_774_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_775 (
    .din     (_zz_1736[35:0]        ), //i
    .dout    (fixTo_775_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_776 (
    .din     (_zz_1737[35:0]        ), //i
    .dout    (fixTo_776_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_777 (
    .din     (_zz_1738[35:0]        ), //i
    .dout    (fixTo_777_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_778 (
    .din     (_zz_1739[35:0]        ), //i
    .dout    (fixTo_778_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_779 (
    .din     (_zz_1740[35:0]        ), //i
    .dout    (fixTo_779_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_780 (
    .din     (_zz_1741[35:0]        ), //i
    .dout    (fixTo_780_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_781 (
    .din     (_zz_1742[35:0]        ), //i
    .dout    (fixTo_781_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_782 (
    .din     (_zz_1743[35:0]        ), //i
    .dout    (fixTo_782_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_783 (
    .din     (_zz_1744[35:0]        ), //i
    .dout    (fixTo_783_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_784 (
    .din     (_zz_1745[35:0]        ), //i
    .dout    (fixTo_784_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_785 (
    .din     (_zz_1746[35:0]        ), //i
    .dout    (fixTo_785_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_786 (
    .din     (_zz_1747[35:0]        ), //i
    .dout    (fixTo_786_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_787 (
    .din     (_zz_1748[35:0]        ), //i
    .dout    (fixTo_787_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_788 (
    .din     (_zz_1749[35:0]        ), //i
    .dout    (fixTo_788_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_789 (
    .din     (_zz_1750[35:0]        ), //i
    .dout    (fixTo_789_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_790 (
    .din     (_zz_1751[35:0]        ), //i
    .dout    (fixTo_790_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_791 (
    .din     (_zz_1752[35:0]        ), //i
    .dout    (fixTo_791_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_792 (
    .din     (_zz_1753[35:0]        ), //i
    .dout    (fixTo_792_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_793 (
    .din     (_zz_1754[35:0]        ), //i
    .dout    (fixTo_793_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_794 (
    .din     (_zz_1755[35:0]        ), //i
    .dout    (fixTo_794_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_795 (
    .din     (_zz_1756[35:0]        ), //i
    .dout    (fixTo_795_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_796 (
    .din     (_zz_1757[35:0]        ), //i
    .dout    (fixTo_796_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_797 (
    .din     (_zz_1758[35:0]        ), //i
    .dout    (fixTo_797_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_798 (
    .din     (_zz_1759[35:0]        ), //i
    .dout    (fixTo_798_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_799 (
    .din     (_zz_1760[35:0]        ), //i
    .dout    (fixTo_799_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_800 (
    .din     (_zz_1761[35:0]        ), //i
    .dout    (fixTo_800_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_801 (
    .din     (_zz_1762[35:0]        ), //i
    .dout    (fixTo_801_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_802 (
    .din     (_zz_1763[35:0]        ), //i
    .dout    (fixTo_802_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_803 (
    .din     (_zz_1764[35:0]        ), //i
    .dout    (fixTo_803_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_804 (
    .din     (_zz_1765[35:0]        ), //i
    .dout    (fixTo_804_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_805 (
    .din     (_zz_1766[35:0]        ), //i
    .dout    (fixTo_805_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_806 (
    .din     (_zz_1767[35:0]        ), //i
    .dout    (fixTo_806_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_807 (
    .din     (_zz_1768[35:0]        ), //i
    .dout    (fixTo_807_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_808 (
    .din     (_zz_1769[35:0]        ), //i
    .dout    (fixTo_808_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_809 (
    .din     (_zz_1770[35:0]        ), //i
    .dout    (fixTo_809_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_810 (
    .din     (_zz_1771[35:0]        ), //i
    .dout    (fixTo_810_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_811 (
    .din     (_zz_1772[35:0]        ), //i
    .dout    (fixTo_811_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_812 (
    .din     (_zz_1773[35:0]        ), //i
    .dout    (fixTo_812_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_813 (
    .din     (_zz_1774[35:0]        ), //i
    .dout    (fixTo_813_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_814 (
    .din     (_zz_1775[35:0]        ), //i
    .dout    (fixTo_814_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_815 (
    .din     (_zz_1776[35:0]        ), //i
    .dout    (fixTo_815_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_816 (
    .din     (_zz_1777[35:0]        ), //i
    .dout    (fixTo_816_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_817 (
    .din     (_zz_1778[35:0]        ), //i
    .dout    (fixTo_817_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_818 (
    .din     (_zz_1779[35:0]        ), //i
    .dout    (fixTo_818_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_819 (
    .din     (_zz_1780[35:0]        ), //i
    .dout    (fixTo_819_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_820 (
    .din     (_zz_1781[35:0]        ), //i
    .dout    (fixTo_820_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_821 (
    .din     (_zz_1782[35:0]        ), //i
    .dout    (fixTo_821_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_822 (
    .din     (_zz_1783[35:0]        ), //i
    .dout    (fixTo_822_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_823 (
    .din     (_zz_1784[35:0]        ), //i
    .dout    (fixTo_823_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_824 (
    .din     (_zz_1785[35:0]        ), //i
    .dout    (fixTo_824_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_825 (
    .din     (_zz_1786[35:0]        ), //i
    .dout    (fixTo_825_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_826 (
    .din     (_zz_1787[35:0]        ), //i
    .dout    (fixTo_826_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_827 (
    .din     (_zz_1788[35:0]        ), //i
    .dout    (fixTo_827_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_828 (
    .din     (_zz_1789[35:0]        ), //i
    .dout    (fixTo_828_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_829 (
    .din     (_zz_1790[35:0]        ), //i
    .dout    (fixTo_829_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_830 (
    .din     (_zz_1791[35:0]        ), //i
    .dout    (fixTo_830_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_831 (
    .din     (_zz_1792[35:0]        ), //i
    .dout    (fixTo_831_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_832 (
    .din     (_zz_1793[35:0]        ), //i
    .dout    (fixTo_832_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_833 (
    .din     (_zz_1794[35:0]        ), //i
    .dout    (fixTo_833_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_834 (
    .din     (_zz_1795[35:0]        ), //i
    .dout    (fixTo_834_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_835 (
    .din     (_zz_1796[35:0]        ), //i
    .dout    (fixTo_835_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_836 (
    .din     (_zz_1797[35:0]        ), //i
    .dout    (fixTo_836_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_837 (
    .din     (_zz_1798[35:0]        ), //i
    .dout    (fixTo_837_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_838 (
    .din     (_zz_1799[35:0]        ), //i
    .dout    (fixTo_838_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_839 (
    .din     (_zz_1800[35:0]        ), //i
    .dout    (fixTo_839_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_840 (
    .din     (_zz_1801[35:0]        ), //i
    .dout    (fixTo_840_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_841 (
    .din     (_zz_1802[35:0]        ), //i
    .dout    (fixTo_841_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_842 (
    .din     (_zz_1803[35:0]        ), //i
    .dout    (fixTo_842_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_843 (
    .din     (_zz_1804[35:0]        ), //i
    .dout    (fixTo_843_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_844 (
    .din     (_zz_1805[35:0]        ), //i
    .dout    (fixTo_844_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_845 (
    .din     (_zz_1806[35:0]        ), //i
    .dout    (fixTo_845_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_846 (
    .din     (_zz_1807[35:0]        ), //i
    .dout    (fixTo_846_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_847 (
    .din     (_zz_1808[35:0]        ), //i
    .dout    (fixTo_847_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_848 (
    .din     (_zz_1809[35:0]        ), //i
    .dout    (fixTo_848_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_849 (
    .din     (_zz_1810[35:0]        ), //i
    .dout    (fixTo_849_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_850 (
    .din     (_zz_1811[35:0]        ), //i
    .dout    (fixTo_850_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_851 (
    .din     (_zz_1812[35:0]        ), //i
    .dout    (fixTo_851_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_852 (
    .din     (_zz_1813[35:0]        ), //i
    .dout    (fixTo_852_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_853 (
    .din     (_zz_1814[35:0]        ), //i
    .dout    (fixTo_853_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_854 (
    .din     (_zz_1815[35:0]        ), //i
    .dout    (fixTo_854_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_855 (
    .din     (_zz_1816[35:0]        ), //i
    .dout    (fixTo_855_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_856 (
    .din     (_zz_1817[35:0]        ), //i
    .dout    (fixTo_856_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_857 (
    .din     (_zz_1818[35:0]        ), //i
    .dout    (fixTo_857_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_858 (
    .din     (_zz_1819[35:0]        ), //i
    .dout    (fixTo_858_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_859 (
    .din     (_zz_1820[35:0]        ), //i
    .dout    (fixTo_859_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_860 (
    .din     (_zz_1821[35:0]        ), //i
    .dout    (fixTo_860_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_861 (
    .din     (_zz_1822[35:0]        ), //i
    .dout    (fixTo_861_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_862 (
    .din     (_zz_1823[35:0]        ), //i
    .dout    (fixTo_862_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_863 (
    .din     (_zz_1824[35:0]        ), //i
    .dout    (fixTo_863_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_864 (
    .din     (_zz_1825[35:0]        ), //i
    .dout    (fixTo_864_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_865 (
    .din     (_zz_1826[35:0]        ), //i
    .dout    (fixTo_865_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_866 (
    .din     (_zz_1827[35:0]        ), //i
    .dout    (fixTo_866_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_867 (
    .din     (_zz_1828[35:0]        ), //i
    .dout    (fixTo_867_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_868 (
    .din     (_zz_1829[35:0]        ), //i
    .dout    (fixTo_868_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_869 (
    .din     (_zz_1830[35:0]        ), //i
    .dout    (fixTo_869_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_870 (
    .din     (_zz_1831[35:0]        ), //i
    .dout    (fixTo_870_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_871 (
    .din     (_zz_1832[35:0]        ), //i
    .dout    (fixTo_871_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_872 (
    .din     (_zz_1833[35:0]        ), //i
    .dout    (fixTo_872_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_873 (
    .din     (_zz_1834[35:0]        ), //i
    .dout    (fixTo_873_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_874 (
    .din     (_zz_1835[35:0]        ), //i
    .dout    (fixTo_874_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_875 (
    .din     (_zz_1836[35:0]        ), //i
    .dout    (fixTo_875_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_876 (
    .din     (_zz_1837[35:0]        ), //i
    .dout    (fixTo_876_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_877 (
    .din     (_zz_1838[35:0]        ), //i
    .dout    (fixTo_877_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_878 (
    .din     (_zz_1839[35:0]        ), //i
    .dout    (fixTo_878_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_879 (
    .din     (_zz_1840[35:0]        ), //i
    .dout    (fixTo_879_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_880 (
    .din     (_zz_1841[35:0]        ), //i
    .dout    (fixTo_880_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_881 (
    .din     (_zz_1842[35:0]        ), //i
    .dout    (fixTo_881_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_882 (
    .din     (_zz_1843[35:0]        ), //i
    .dout    (fixTo_882_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_883 (
    .din     (_zz_1844[35:0]        ), //i
    .dout    (fixTo_883_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_884 (
    .din     (_zz_1845[35:0]        ), //i
    .dout    (fixTo_884_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_885 (
    .din     (_zz_1846[35:0]        ), //i
    .dout    (fixTo_885_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_886 (
    .din     (_zz_1847[35:0]        ), //i
    .dout    (fixTo_886_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_887 (
    .din     (_zz_1848[35:0]        ), //i
    .dout    (fixTo_887_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_888 (
    .din     (_zz_1849[35:0]        ), //i
    .dout    (fixTo_888_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_889 (
    .din     (_zz_1850[35:0]        ), //i
    .dout    (fixTo_889_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_890 (
    .din     (_zz_1851[35:0]        ), //i
    .dout    (fixTo_890_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_891 (
    .din     (_zz_1852[35:0]        ), //i
    .dout    (fixTo_891_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_892 (
    .din     (_zz_1853[35:0]        ), //i
    .dout    (fixTo_892_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_893 (
    .din     (_zz_1854[35:0]        ), //i
    .dout    (fixTo_893_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_894 (
    .din     (_zz_1855[35:0]        ), //i
    .dout    (fixTo_894_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_895 (
    .din     (_zz_1856[35:0]        ), //i
    .dout    (fixTo_895_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_896 (
    .din     (_zz_1857[35:0]        ), //i
    .dout    (fixTo_896_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_897 (
    .din     (_zz_1858[35:0]        ), //i
    .dout    (fixTo_897_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_898 (
    .din     (_zz_1859[35:0]        ), //i
    .dout    (fixTo_898_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_899 (
    .din     (_zz_1860[35:0]        ), //i
    .dout    (fixTo_899_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_900 (
    .din     (_zz_1861[35:0]        ), //i
    .dout    (fixTo_900_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_901 (
    .din     (_zz_1862[35:0]        ), //i
    .dout    (fixTo_901_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_902 (
    .din     (_zz_1863[35:0]        ), //i
    .dout    (fixTo_902_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_903 (
    .din     (_zz_1864[35:0]        ), //i
    .dout    (fixTo_903_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_904 (
    .din     (_zz_1865[35:0]        ), //i
    .dout    (fixTo_904_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_905 (
    .din     (_zz_1866[35:0]        ), //i
    .dout    (fixTo_905_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_906 (
    .din     (_zz_1867[35:0]        ), //i
    .dout    (fixTo_906_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_907 (
    .din     (_zz_1868[35:0]        ), //i
    .dout    (fixTo_907_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_908 (
    .din     (_zz_1869[35:0]        ), //i
    .dout    (fixTo_908_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_909 (
    .din     (_zz_1870[35:0]        ), //i
    .dout    (fixTo_909_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_910 (
    .din     (_zz_1871[35:0]        ), //i
    .dout    (fixTo_910_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_911 (
    .din     (_zz_1872[35:0]        ), //i
    .dout    (fixTo_911_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_912 (
    .din     (_zz_1873[35:0]        ), //i
    .dout    (fixTo_912_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_913 (
    .din     (_zz_1874[35:0]        ), //i
    .dout    (fixTo_913_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_914 (
    .din     (_zz_1875[35:0]        ), //i
    .dout    (fixTo_914_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_915 (
    .din     (_zz_1876[35:0]        ), //i
    .dout    (fixTo_915_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_916 (
    .din     (_zz_1877[35:0]        ), //i
    .dout    (fixTo_916_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_917 (
    .din     (_zz_1878[35:0]        ), //i
    .dout    (fixTo_917_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_918 (
    .din     (_zz_1879[35:0]        ), //i
    .dout    (fixTo_918_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_919 (
    .din     (_zz_1880[35:0]        ), //i
    .dout    (fixTo_919_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_920 (
    .din     (_zz_1881[35:0]        ), //i
    .dout    (fixTo_920_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_921 (
    .din     (_zz_1882[35:0]        ), //i
    .dout    (fixTo_921_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_922 (
    .din     (_zz_1883[35:0]        ), //i
    .dout    (fixTo_922_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_923 (
    .din     (_zz_1884[35:0]        ), //i
    .dout    (fixTo_923_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_924 (
    .din     (_zz_1885[35:0]        ), //i
    .dout    (fixTo_924_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_925 (
    .din     (_zz_1886[35:0]        ), //i
    .dout    (fixTo_925_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_926 (
    .din     (_zz_1887[35:0]        ), //i
    .dout    (fixTo_926_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_927 (
    .din     (_zz_1888[35:0]        ), //i
    .dout    (fixTo_927_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_928 (
    .din     (_zz_1889[35:0]        ), //i
    .dout    (fixTo_928_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_929 (
    .din     (_zz_1890[35:0]        ), //i
    .dout    (fixTo_929_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_930 (
    .din     (_zz_1891[35:0]        ), //i
    .dout    (fixTo_930_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_931 (
    .din     (_zz_1892[35:0]        ), //i
    .dout    (fixTo_931_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_932 (
    .din     (_zz_1893[35:0]        ), //i
    .dout    (fixTo_932_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_933 (
    .din     (_zz_1894[35:0]        ), //i
    .dout    (fixTo_933_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_934 (
    .din     (_zz_1895[35:0]        ), //i
    .dout    (fixTo_934_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_935 (
    .din     (_zz_1896[35:0]        ), //i
    .dout    (fixTo_935_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_936 (
    .din     (_zz_1897[35:0]        ), //i
    .dout    (fixTo_936_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_937 (
    .din     (_zz_1898[35:0]        ), //i
    .dout    (fixTo_937_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_938 (
    .din     (_zz_1899[35:0]        ), //i
    .dout    (fixTo_938_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_939 (
    .din     (_zz_1900[35:0]        ), //i
    .dout    (fixTo_939_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_940 (
    .din     (_zz_1901[35:0]        ), //i
    .dout    (fixTo_940_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_941 (
    .din     (_zz_1902[35:0]        ), //i
    .dout    (fixTo_941_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_942 (
    .din     (_zz_1903[35:0]        ), //i
    .dout    (fixTo_942_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_943 (
    .din     (_zz_1904[35:0]        ), //i
    .dout    (fixTo_943_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_944 (
    .din     (_zz_1905[35:0]        ), //i
    .dout    (fixTo_944_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_945 (
    .din     (_zz_1906[35:0]        ), //i
    .dout    (fixTo_945_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_946 (
    .din     (_zz_1907[35:0]        ), //i
    .dout    (fixTo_946_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_947 (
    .din     (_zz_1908[35:0]        ), //i
    .dout    (fixTo_947_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_948 (
    .din     (_zz_1909[35:0]        ), //i
    .dout    (fixTo_948_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_949 (
    .din     (_zz_1910[35:0]        ), //i
    .dout    (fixTo_949_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_950 (
    .din     (_zz_1911[35:0]        ), //i
    .dout    (fixTo_950_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_951 (
    .din     (_zz_1912[35:0]        ), //i
    .dout    (fixTo_951_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_952 (
    .din     (_zz_1913[35:0]        ), //i
    .dout    (fixTo_952_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_953 (
    .din     (_zz_1914[35:0]        ), //i
    .dout    (fixTo_953_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_954 (
    .din     (_zz_1915[35:0]        ), //i
    .dout    (fixTo_954_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_955 (
    .din     (_zz_1916[35:0]        ), //i
    .dout    (fixTo_955_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_956 (
    .din     (_zz_1917[35:0]        ), //i
    .dout    (fixTo_956_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_957 (
    .din     (_zz_1918[35:0]        ), //i
    .dout    (fixTo_957_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_958 (
    .din     (_zz_1919[35:0]        ), //i
    .dout    (fixTo_958_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_959 (
    .din     (_zz_1920[35:0]        ), //i
    .dout    (fixTo_959_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_960 (
    .din     (_zz_1921[35:0]        ), //i
    .dout    (fixTo_960_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_961 (
    .din     (_zz_1922[35:0]        ), //i
    .dout    (fixTo_961_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_962 (
    .din     (_zz_1923[35:0]        ), //i
    .dout    (fixTo_962_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_963 (
    .din     (_zz_1924[35:0]        ), //i
    .dout    (fixTo_963_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_964 (
    .din     (_zz_1925[35:0]        ), //i
    .dout    (fixTo_964_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_965 (
    .din     (_zz_1926[35:0]        ), //i
    .dout    (fixTo_965_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_966 (
    .din     (_zz_1927[35:0]        ), //i
    .dout    (fixTo_966_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_967 (
    .din     (_zz_1928[35:0]        ), //i
    .dout    (fixTo_967_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_968 (
    .din     (_zz_1929[35:0]        ), //i
    .dout    (fixTo_968_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_969 (
    .din     (_zz_1930[35:0]        ), //i
    .dout    (fixTo_969_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_970 (
    .din     (_zz_1931[35:0]        ), //i
    .dout    (fixTo_970_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_971 (
    .din     (_zz_1932[35:0]        ), //i
    .dout    (fixTo_971_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_972 (
    .din     (_zz_1933[35:0]        ), //i
    .dout    (fixTo_972_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_973 (
    .din     (_zz_1934[35:0]        ), //i
    .dout    (fixTo_973_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_974 (
    .din     (_zz_1935[35:0]        ), //i
    .dout    (fixTo_974_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_975 (
    .din     (_zz_1936[35:0]        ), //i
    .dout    (fixTo_975_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_976 (
    .din     (_zz_1937[35:0]        ), //i
    .dout    (fixTo_976_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_977 (
    .din     (_zz_1938[35:0]        ), //i
    .dout    (fixTo_977_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_978 (
    .din     (_zz_1939[35:0]        ), //i
    .dout    (fixTo_978_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_979 (
    .din     (_zz_1940[35:0]        ), //i
    .dout    (fixTo_979_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_980 (
    .din     (_zz_1941[35:0]        ), //i
    .dout    (fixTo_980_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_981 (
    .din     (_zz_1942[35:0]        ), //i
    .dout    (fixTo_981_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_982 (
    .din     (_zz_1943[35:0]        ), //i
    .dout    (fixTo_982_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_983 (
    .din     (_zz_1944[35:0]        ), //i
    .dout    (fixTo_983_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_984 (
    .din     (_zz_1945[35:0]        ), //i
    .dout    (fixTo_984_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_985 (
    .din     (_zz_1946[35:0]        ), //i
    .dout    (fixTo_985_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_986 (
    .din     (_zz_1947[35:0]        ), //i
    .dout    (fixTo_986_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_987 (
    .din     (_zz_1948[35:0]        ), //i
    .dout    (fixTo_987_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_988 (
    .din     (_zz_1949[35:0]        ), //i
    .dout    (fixTo_988_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_989 (
    .din     (_zz_1950[35:0]        ), //i
    .dout    (fixTo_989_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_990 (
    .din     (_zz_1951[35:0]        ), //i
    .dout    (fixTo_990_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_991 (
    .din     (_zz_1952[35:0]        ), //i
    .dout    (fixTo_991_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_992 (
    .din     (_zz_1953[35:0]        ), //i
    .dout    (fixTo_992_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_993 (
    .din     (_zz_1954[35:0]        ), //i
    .dout    (fixTo_993_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_994 (
    .din     (_zz_1955[35:0]        ), //i
    .dout    (fixTo_994_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_995 (
    .din     (_zz_1956[35:0]        ), //i
    .dout    (fixTo_995_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_996 (
    .din     (_zz_1957[35:0]        ), //i
    .dout    (fixTo_996_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_997 (
    .din     (_zz_1958[35:0]        ), //i
    .dout    (fixTo_997_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_998 (
    .din     (_zz_1959[35:0]        ), //i
    .dout    (fixTo_998_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_999 (
    .din     (_zz_1960[35:0]        ), //i
    .dout    (fixTo_999_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1000 (
    .din     (_zz_1961[35:0]         ), //i
    .dout    (fixTo_1000_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1001 (
    .din     (_zz_1962[35:0]         ), //i
    .dout    (fixTo_1001_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1002 (
    .din     (_zz_1963[35:0]         ), //i
    .dout    (fixTo_1002_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1003 (
    .din     (_zz_1964[35:0]         ), //i
    .dout    (fixTo_1003_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1004 (
    .din     (_zz_1965[35:0]         ), //i
    .dout    (fixTo_1004_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1005 (
    .din     (_zz_1966[35:0]         ), //i
    .dout    (fixTo_1005_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1006 (
    .din     (_zz_1967[35:0]         ), //i
    .dout    (fixTo_1006_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1007 (
    .din     (_zz_1968[35:0]         ), //i
    .dout    (fixTo_1007_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1008 (
    .din     (_zz_1969[35:0]         ), //i
    .dout    (fixTo_1008_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1009 (
    .din     (_zz_1970[35:0]         ), //i
    .dout    (fixTo_1009_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1010 (
    .din     (_zz_1971[35:0]         ), //i
    .dout    (fixTo_1010_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1011 (
    .din     (_zz_1972[35:0]         ), //i
    .dout    (fixTo_1011_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1012 (
    .din     (_zz_1973[35:0]         ), //i
    .dout    (fixTo_1012_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1013 (
    .din     (_zz_1974[35:0]         ), //i
    .dout    (fixTo_1013_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1014 (
    .din     (_zz_1975[35:0]         ), //i
    .dout    (fixTo_1014_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1015 (
    .din     (_zz_1976[35:0]         ), //i
    .dout    (fixTo_1015_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1016 (
    .din     (_zz_1977[35:0]         ), //i
    .dout    (fixTo_1016_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1017 (
    .din     (_zz_1978[35:0]         ), //i
    .dout    (fixTo_1017_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1018 (
    .din     (_zz_1979[35:0]         ), //i
    .dout    (fixTo_1018_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1019 (
    .din     (_zz_1980[35:0]         ), //i
    .dout    (fixTo_1019_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1020 (
    .din     (_zz_1981[35:0]         ), //i
    .dout    (fixTo_1020_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1021 (
    .din     (_zz_1982[35:0]         ), //i
    .dout    (fixTo_1021_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1022 (
    .din     (_zz_1983[35:0]         ), //i
    .dout    (fixTo_1022_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1023 (
    .din     (_zz_1984[35:0]         ), //i
    .dout    (fixTo_1023_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1024 (
    .din     (_zz_1985[35:0]         ), //i
    .dout    (fixTo_1024_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1025 (
    .din     (_zz_1986[35:0]         ), //i
    .dout    (fixTo_1025_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1026 (
    .din     (_zz_1987[35:0]         ), //i
    .dout    (fixTo_1026_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1027 (
    .din     (_zz_1988[35:0]         ), //i
    .dout    (fixTo_1027_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1028 (
    .din     (_zz_1989[35:0]         ), //i
    .dout    (fixTo_1028_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1029 (
    .din     (_zz_1990[35:0]         ), //i
    .dout    (fixTo_1029_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1030 (
    .din     (_zz_1991[35:0]         ), //i
    .dout    (fixTo_1030_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1031 (
    .din     (_zz_1992[35:0]         ), //i
    .dout    (fixTo_1031_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1032 (
    .din     (_zz_1993[35:0]         ), //i
    .dout    (fixTo_1032_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1033 (
    .din     (_zz_1994[35:0]         ), //i
    .dout    (fixTo_1033_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1034 (
    .din     (_zz_1995[35:0]         ), //i
    .dout    (fixTo_1034_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1035 (
    .din     (_zz_1996[35:0]         ), //i
    .dout    (fixTo_1035_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1036 (
    .din     (_zz_1997[35:0]         ), //i
    .dout    (fixTo_1036_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1037 (
    .din     (_zz_1998[35:0]         ), //i
    .dout    (fixTo_1037_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1038 (
    .din     (_zz_1999[35:0]         ), //i
    .dout    (fixTo_1038_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1039 (
    .din     (_zz_2000[35:0]         ), //i
    .dout    (fixTo_1039_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1040 (
    .din     (_zz_2001[35:0]         ), //i
    .dout    (fixTo_1040_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1041 (
    .din     (_zz_2002[35:0]         ), //i
    .dout    (fixTo_1041_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1042 (
    .din     (_zz_2003[35:0]         ), //i
    .dout    (fixTo_1042_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1043 (
    .din     (_zz_2004[35:0]         ), //i
    .dout    (fixTo_1043_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1044 (
    .din     (_zz_2005[35:0]         ), //i
    .dout    (fixTo_1044_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1045 (
    .din     (_zz_2006[35:0]         ), //i
    .dout    (fixTo_1045_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1046 (
    .din     (_zz_2007[35:0]         ), //i
    .dout    (fixTo_1046_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1047 (
    .din     (_zz_2008[35:0]         ), //i
    .dout    (fixTo_1047_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1048 (
    .din     (_zz_2009[35:0]         ), //i
    .dout    (fixTo_1048_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1049 (
    .din     (_zz_2010[35:0]         ), //i
    .dout    (fixTo_1049_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1050 (
    .din     (_zz_2011[35:0]         ), //i
    .dout    (fixTo_1050_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1051 (
    .din     (_zz_2012[35:0]         ), //i
    .dout    (fixTo_1051_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1052 (
    .din     (_zz_2013[35:0]         ), //i
    .dout    (fixTo_1052_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1053 (
    .din     (_zz_2014[35:0]         ), //i
    .dout    (fixTo_1053_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1054 (
    .din     (_zz_2015[35:0]         ), //i
    .dout    (fixTo_1054_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1055 (
    .din     (_zz_2016[35:0]         ), //i
    .dout    (fixTo_1055_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1056 (
    .din     (_zz_2017[35:0]         ), //i
    .dout    (fixTo_1056_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1057 (
    .din     (_zz_2018[35:0]         ), //i
    .dout    (fixTo_1057_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1058 (
    .din     (_zz_2019[35:0]         ), //i
    .dout    (fixTo_1058_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1059 (
    .din     (_zz_2020[35:0]         ), //i
    .dout    (fixTo_1059_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1060 (
    .din     (_zz_2021[35:0]         ), //i
    .dout    (fixTo_1060_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1061 (
    .din     (_zz_2022[35:0]         ), //i
    .dout    (fixTo_1061_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1062 (
    .din     (_zz_2023[35:0]         ), //i
    .dout    (fixTo_1062_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1063 (
    .din     (_zz_2024[35:0]         ), //i
    .dout    (fixTo_1063_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1064 (
    .din     (_zz_2025[35:0]         ), //i
    .dout    (fixTo_1064_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1065 (
    .din     (_zz_2026[35:0]         ), //i
    .dout    (fixTo_1065_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1066 (
    .din     (_zz_2027[35:0]         ), //i
    .dout    (fixTo_1066_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1067 (
    .din     (_zz_2028[35:0]         ), //i
    .dout    (fixTo_1067_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1068 (
    .din     (_zz_2029[35:0]         ), //i
    .dout    (fixTo_1068_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1069 (
    .din     (_zz_2030[35:0]         ), //i
    .dout    (fixTo_1069_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1070 (
    .din     (_zz_2031[35:0]         ), //i
    .dout    (fixTo_1070_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1071 (
    .din     (_zz_2032[35:0]         ), //i
    .dout    (fixTo_1071_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1072 (
    .din     (_zz_2033[35:0]         ), //i
    .dout    (fixTo_1072_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1073 (
    .din     (_zz_2034[35:0]         ), //i
    .dout    (fixTo_1073_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1074 (
    .din     (_zz_2035[35:0]         ), //i
    .dout    (fixTo_1074_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1075 (
    .din     (_zz_2036[35:0]         ), //i
    .dout    (fixTo_1075_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1076 (
    .din     (_zz_2037[35:0]         ), //i
    .dout    (fixTo_1076_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1077 (
    .din     (_zz_2038[35:0]         ), //i
    .dout    (fixTo_1077_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1078 (
    .din     (_zz_2039[35:0]         ), //i
    .dout    (fixTo_1078_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1079 (
    .din     (_zz_2040[35:0]         ), //i
    .dout    (fixTo_1079_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1080 (
    .din     (_zz_2041[35:0]         ), //i
    .dout    (fixTo_1080_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1081 (
    .din     (_zz_2042[35:0]         ), //i
    .dout    (fixTo_1081_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1082 (
    .din     (_zz_2043[35:0]         ), //i
    .dout    (fixTo_1082_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1083 (
    .din     (_zz_2044[35:0]         ), //i
    .dout    (fixTo_1083_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1084 (
    .din     (_zz_2045[35:0]         ), //i
    .dout    (fixTo_1084_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1085 (
    .din     (_zz_2046[35:0]         ), //i
    .dout    (fixTo_1085_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1086 (
    .din     (_zz_2047[35:0]         ), //i
    .dout    (fixTo_1086_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1087 (
    .din     (_zz_2048[35:0]         ), //i
    .dout    (fixTo_1087_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1088 (
    .din     (_zz_2049[35:0]         ), //i
    .dout    (fixTo_1088_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1089 (
    .din     (_zz_2050[35:0]         ), //i
    .dout    (fixTo_1089_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1090 (
    .din     (_zz_2051[35:0]         ), //i
    .dout    (fixTo_1090_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1091 (
    .din     (_zz_2052[35:0]         ), //i
    .dout    (fixTo_1091_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1092 (
    .din     (_zz_2053[35:0]         ), //i
    .dout    (fixTo_1092_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1093 (
    .din     (_zz_2054[35:0]         ), //i
    .dout    (fixTo_1093_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1094 (
    .din     (_zz_2055[35:0]         ), //i
    .dout    (fixTo_1094_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1095 (
    .din     (_zz_2056[35:0]         ), //i
    .dout    (fixTo_1095_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1096 (
    .din     (_zz_2057[35:0]         ), //i
    .dout    (fixTo_1096_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1097 (
    .din     (_zz_2058[35:0]         ), //i
    .dout    (fixTo_1097_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1098 (
    .din     (_zz_2059[35:0]         ), //i
    .dout    (fixTo_1098_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1099 (
    .din     (_zz_2060[35:0]         ), //i
    .dout    (fixTo_1099_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1100 (
    .din     (_zz_2061[35:0]         ), //i
    .dout    (fixTo_1100_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1101 (
    .din     (_zz_2062[35:0]         ), //i
    .dout    (fixTo_1101_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1102 (
    .din     (_zz_2063[35:0]         ), //i
    .dout    (fixTo_1102_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1103 (
    .din     (_zz_2064[35:0]         ), //i
    .dout    (fixTo_1103_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1104 (
    .din     (_zz_2065[35:0]         ), //i
    .dout    (fixTo_1104_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1105 (
    .din     (_zz_2066[35:0]         ), //i
    .dout    (fixTo_1105_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1106 (
    .din     (_zz_2067[35:0]         ), //i
    .dout    (fixTo_1106_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1107 (
    .din     (_zz_2068[35:0]         ), //i
    .dout    (fixTo_1107_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1108 (
    .din     (_zz_2069[35:0]         ), //i
    .dout    (fixTo_1108_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1109 (
    .din     (_zz_2070[35:0]         ), //i
    .dout    (fixTo_1109_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1110 (
    .din     (_zz_2071[35:0]         ), //i
    .dout    (fixTo_1110_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1111 (
    .din     (_zz_2072[35:0]         ), //i
    .dout    (fixTo_1111_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1112 (
    .din     (_zz_2073[35:0]         ), //i
    .dout    (fixTo_1112_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1113 (
    .din     (_zz_2074[35:0]         ), //i
    .dout    (fixTo_1113_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1114 (
    .din     (_zz_2075[35:0]         ), //i
    .dout    (fixTo_1114_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1115 (
    .din     (_zz_2076[35:0]         ), //i
    .dout    (fixTo_1115_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1116 (
    .din     (_zz_2077[35:0]         ), //i
    .dout    (fixTo_1116_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1117 (
    .din     (_zz_2078[35:0]         ), //i
    .dout    (fixTo_1117_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1118 (
    .din     (_zz_2079[35:0]         ), //i
    .dout    (fixTo_1118_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1119 (
    .din     (_zz_2080[35:0]         ), //i
    .dout    (fixTo_1119_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1120 (
    .din     (_zz_2081[35:0]         ), //i
    .dout    (fixTo_1120_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1121 (
    .din     (_zz_2082[35:0]         ), //i
    .dout    (fixTo_1121_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1122 (
    .din     (_zz_2083[35:0]         ), //i
    .dout    (fixTo_1122_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1123 (
    .din     (_zz_2084[35:0]         ), //i
    .dout    (fixTo_1123_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1124 (
    .din     (_zz_2085[35:0]         ), //i
    .dout    (fixTo_1124_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1125 (
    .din     (_zz_2086[35:0]         ), //i
    .dout    (fixTo_1125_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1126 (
    .din     (_zz_2087[35:0]         ), //i
    .dout    (fixTo_1126_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1127 (
    .din     (_zz_2088[35:0]         ), //i
    .dout    (fixTo_1127_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1128 (
    .din     (_zz_2089[35:0]         ), //i
    .dout    (fixTo_1128_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1129 (
    .din     (_zz_2090[35:0]         ), //i
    .dout    (fixTo_1129_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1130 (
    .din     (_zz_2091[35:0]         ), //i
    .dout    (fixTo_1130_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1131 (
    .din     (_zz_2092[35:0]         ), //i
    .dout    (fixTo_1131_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1132 (
    .din     (_zz_2093[35:0]         ), //i
    .dout    (fixTo_1132_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1133 (
    .din     (_zz_2094[35:0]         ), //i
    .dout    (fixTo_1133_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1134 (
    .din     (_zz_2095[35:0]         ), //i
    .dout    (fixTo_1134_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1135 (
    .din     (_zz_2096[35:0]         ), //i
    .dout    (fixTo_1135_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1136 (
    .din     (_zz_2097[35:0]         ), //i
    .dout    (fixTo_1136_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1137 (
    .din     (_zz_2098[35:0]         ), //i
    .dout    (fixTo_1137_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1138 (
    .din     (_zz_2099[35:0]         ), //i
    .dout    (fixTo_1138_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1139 (
    .din     (_zz_2100[35:0]         ), //i
    .dout    (fixTo_1139_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1140 (
    .din     (_zz_2101[35:0]         ), //i
    .dout    (fixTo_1140_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1141 (
    .din     (_zz_2102[35:0]         ), //i
    .dout    (fixTo_1141_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1142 (
    .din     (_zz_2103[35:0]         ), //i
    .dout    (fixTo_1142_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1143 (
    .din     (_zz_2104[35:0]         ), //i
    .dout    (fixTo_1143_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1144 (
    .din     (_zz_2105[35:0]         ), //i
    .dout    (fixTo_1144_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1145 (
    .din     (_zz_2106[35:0]         ), //i
    .dout    (fixTo_1145_dout[17:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1146 (
    .din     (_zz_2107[35:0]         ), //i
    .dout    (fixTo_1146_dout[35:0]  )  //o
  );
  SInt36fixTo35_0_ROUNDTOINF fixTo_1147 (
    .din     (_zz_2108[35:0]         ), //i
    .dout    (fixTo_1147_dout[35:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1148 (
    .din     (_zz_2109[35:0]         ), //i
    .dout    (fixTo_1148_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1149 (
    .din     (_zz_2110[35:0]         ), //i
    .dout    (fixTo_1149_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1150 (
    .din     (_zz_2111[35:0]         ), //i
    .dout    (fixTo_1150_dout[17:0]  )  //o
  );
  SInt36fixTo26_9_ROUNDTOINF fixTo_1151 (
    .din     (_zz_2112[35:0]         ), //i
    .dout    (fixTo_1151_dout[17:0]  )  //o
  );
  assign twiddle_factor_table_0_real = 18'h00200;
  assign twiddle_factor_table_0_imag = 18'h0;
  assign twiddle_factor_table_1_real = 18'h00200;
  assign twiddle_factor_table_1_imag = 18'h0;
  assign twiddle_factor_table_2_real = 18'h0;
  assign twiddle_factor_table_2_imag = 18'h3fe00;
  assign twiddle_factor_table_3_real = 18'h00200;
  assign twiddle_factor_table_3_imag = 18'h0;
  assign twiddle_factor_table_4_real = 18'h0016a;
  assign twiddle_factor_table_4_imag = 18'h3fe96;
  assign twiddle_factor_table_5_real = 18'h0;
  assign twiddle_factor_table_5_imag = 18'h3fe00;
  assign twiddle_factor_table_6_real = 18'h3fe96;
  assign twiddle_factor_table_6_imag = 18'h3fe96;
  assign twiddle_factor_table_7_real = 18'h00200;
  assign twiddle_factor_table_7_imag = 18'h0;
  assign twiddle_factor_table_8_real = 18'h001d9;
  assign twiddle_factor_table_8_imag = 18'h3ff3d;
  assign twiddle_factor_table_9_real = 18'h0016a;
  assign twiddle_factor_table_9_imag = 18'h3fe96;
  assign twiddle_factor_table_10_real = 18'h000c3;
  assign twiddle_factor_table_10_imag = 18'h3fe27;
  assign twiddle_factor_table_11_real = 18'h0;
  assign twiddle_factor_table_11_imag = 18'h3fe00;
  assign twiddle_factor_table_12_real = 18'h3ff3d;
  assign twiddle_factor_table_12_imag = 18'h3fe27;
  assign twiddle_factor_table_13_real = 18'h3fe96;
  assign twiddle_factor_table_13_imag = 18'h3fe96;
  assign twiddle_factor_table_14_real = 18'h3fe27;
  assign twiddle_factor_table_14_imag = 18'h3ff3d;
  assign twiddle_factor_table_15_real = 18'h00200;
  assign twiddle_factor_table_15_imag = 18'h0;
  assign twiddle_factor_table_16_real = 18'h001f6;
  assign twiddle_factor_table_16_imag = 18'h3ff9d;
  assign twiddle_factor_table_17_real = 18'h001d9;
  assign twiddle_factor_table_17_imag = 18'h3ff3d;
  assign twiddle_factor_table_18_real = 18'h001a9;
  assign twiddle_factor_table_18_imag = 18'h3fee4;
  assign twiddle_factor_table_19_real = 18'h0016a;
  assign twiddle_factor_table_19_imag = 18'h3fe96;
  assign twiddle_factor_table_20_real = 18'h0011c;
  assign twiddle_factor_table_20_imag = 18'h3fe57;
  assign twiddle_factor_table_21_real = 18'h000c3;
  assign twiddle_factor_table_21_imag = 18'h3fe27;
  assign twiddle_factor_table_22_real = 18'h00063;
  assign twiddle_factor_table_22_imag = 18'h3fe0a;
  assign twiddle_factor_table_23_real = 18'h0;
  assign twiddle_factor_table_23_imag = 18'h3fe00;
  assign twiddle_factor_table_24_real = 18'h3ff9d;
  assign twiddle_factor_table_24_imag = 18'h3fe0a;
  assign twiddle_factor_table_25_real = 18'h3ff3d;
  assign twiddle_factor_table_25_imag = 18'h3fe27;
  assign twiddle_factor_table_26_real = 18'h3fee4;
  assign twiddle_factor_table_26_imag = 18'h3fe57;
  assign twiddle_factor_table_27_real = 18'h3fe96;
  assign twiddle_factor_table_27_imag = 18'h3fe96;
  assign twiddle_factor_table_28_real = 18'h3fe57;
  assign twiddle_factor_table_28_imag = 18'h3fee4;
  assign twiddle_factor_table_29_real = 18'h3fe27;
  assign twiddle_factor_table_29_imag = 18'h3ff3d;
  assign twiddle_factor_table_30_real = 18'h3fe0a;
  assign twiddle_factor_table_30_imag = 18'h3ff9d;
  assign twiddle_factor_table_31_real = 18'h00200;
  assign twiddle_factor_table_31_imag = 18'h0;
  assign twiddle_factor_table_32_real = 18'h001fd;
  assign twiddle_factor_table_32_imag = 18'h3ffce;
  assign twiddle_factor_table_33_real = 18'h001f6;
  assign twiddle_factor_table_33_imag = 18'h3ff9d;
  assign twiddle_factor_table_34_real = 18'h001e9;
  assign twiddle_factor_table_34_imag = 18'h3ff6c;
  assign twiddle_factor_table_35_real = 18'h001d9;
  assign twiddle_factor_table_35_imag = 18'h3ff3d;
  assign twiddle_factor_table_36_real = 18'h001c3;
  assign twiddle_factor_table_36_imag = 18'h3ff0f;
  assign twiddle_factor_table_37_real = 18'h001a9;
  assign twiddle_factor_table_37_imag = 18'h3fee4;
  assign twiddle_factor_table_38_real = 18'h0018b;
  assign twiddle_factor_table_38_imag = 18'h3febc;
  assign twiddle_factor_table_39_real = 18'h0016a;
  assign twiddle_factor_table_39_imag = 18'h3fe96;
  assign twiddle_factor_table_40_real = 18'h00144;
  assign twiddle_factor_table_40_imag = 18'h3fe75;
  assign twiddle_factor_table_41_real = 18'h0011c;
  assign twiddle_factor_table_41_imag = 18'h3fe57;
  assign twiddle_factor_table_42_real = 18'h000f1;
  assign twiddle_factor_table_42_imag = 18'h3fe3d;
  assign twiddle_factor_table_43_real = 18'h000c3;
  assign twiddle_factor_table_43_imag = 18'h3fe27;
  assign twiddle_factor_table_44_real = 18'h00094;
  assign twiddle_factor_table_44_imag = 18'h3fe17;
  assign twiddle_factor_table_45_real = 18'h00063;
  assign twiddle_factor_table_45_imag = 18'h3fe0a;
  assign twiddle_factor_table_46_real = 18'h00032;
  assign twiddle_factor_table_46_imag = 18'h3fe03;
  assign twiddle_factor_table_47_real = 18'h0;
  assign twiddle_factor_table_47_imag = 18'h3fe00;
  assign twiddle_factor_table_48_real = 18'h3ffce;
  assign twiddle_factor_table_48_imag = 18'h3fe03;
  assign twiddle_factor_table_49_real = 18'h3ff9d;
  assign twiddle_factor_table_49_imag = 18'h3fe0a;
  assign twiddle_factor_table_50_real = 18'h3ff6c;
  assign twiddle_factor_table_50_imag = 18'h3fe17;
  assign twiddle_factor_table_51_real = 18'h3ff3d;
  assign twiddle_factor_table_51_imag = 18'h3fe27;
  assign twiddle_factor_table_52_real = 18'h3ff0f;
  assign twiddle_factor_table_52_imag = 18'h3fe3d;
  assign twiddle_factor_table_53_real = 18'h3fee4;
  assign twiddle_factor_table_53_imag = 18'h3fe57;
  assign twiddle_factor_table_54_real = 18'h3febc;
  assign twiddle_factor_table_54_imag = 18'h3fe75;
  assign twiddle_factor_table_55_real = 18'h3fe96;
  assign twiddle_factor_table_55_imag = 18'h3fe96;
  assign twiddle_factor_table_56_real = 18'h3fe75;
  assign twiddle_factor_table_56_imag = 18'h3febc;
  assign twiddle_factor_table_57_real = 18'h3fe57;
  assign twiddle_factor_table_57_imag = 18'h3fee4;
  assign twiddle_factor_table_58_real = 18'h3fe3d;
  assign twiddle_factor_table_58_imag = 18'h3ff0f;
  assign twiddle_factor_table_59_real = 18'h3fe27;
  assign twiddle_factor_table_59_imag = 18'h3ff3d;
  assign twiddle_factor_table_60_real = 18'h3fe17;
  assign twiddle_factor_table_60_imag = 18'h3ff6c;
  assign twiddle_factor_table_61_real = 18'h3fe0a;
  assign twiddle_factor_table_61_imag = 18'h3ff9d;
  assign twiddle_factor_table_62_real = 18'h3fe03;
  assign twiddle_factor_table_62_imag = 18'h3ffce;
  assign data_reorder_0_real = data_in_0_real;
  assign data_reorder_0_imag = data_in_0_imag;
  assign data_reorder_32_real = data_in_1_real;
  assign data_reorder_32_imag = data_in_1_imag;
  assign data_reorder_16_real = data_in_2_real;
  assign data_reorder_16_imag = data_in_2_imag;
  assign data_reorder_48_real = data_in_3_real;
  assign data_reorder_48_imag = data_in_3_imag;
  assign data_reorder_8_real = data_in_4_real;
  assign data_reorder_8_imag = data_in_4_imag;
  assign data_reorder_40_real = data_in_5_real;
  assign data_reorder_40_imag = data_in_5_imag;
  assign data_reorder_24_real = data_in_6_real;
  assign data_reorder_24_imag = data_in_6_imag;
  assign data_reorder_56_real = data_in_7_real;
  assign data_reorder_56_imag = data_in_7_imag;
  assign data_reorder_4_real = data_in_8_real;
  assign data_reorder_4_imag = data_in_8_imag;
  assign data_reorder_36_real = data_in_9_real;
  assign data_reorder_36_imag = data_in_9_imag;
  assign data_reorder_20_real = data_in_10_real;
  assign data_reorder_20_imag = data_in_10_imag;
  assign data_reorder_52_real = data_in_11_real;
  assign data_reorder_52_imag = data_in_11_imag;
  assign data_reorder_12_real = data_in_12_real;
  assign data_reorder_12_imag = data_in_12_imag;
  assign data_reorder_44_real = data_in_13_real;
  assign data_reorder_44_imag = data_in_13_imag;
  assign data_reorder_28_real = data_in_14_real;
  assign data_reorder_28_imag = data_in_14_imag;
  assign data_reorder_60_real = data_in_15_real;
  assign data_reorder_60_imag = data_in_15_imag;
  assign data_reorder_2_real = data_in_16_real;
  assign data_reorder_2_imag = data_in_16_imag;
  assign data_reorder_34_real = data_in_17_real;
  assign data_reorder_34_imag = data_in_17_imag;
  assign data_reorder_18_real = data_in_18_real;
  assign data_reorder_18_imag = data_in_18_imag;
  assign data_reorder_50_real = data_in_19_real;
  assign data_reorder_50_imag = data_in_19_imag;
  assign data_reorder_10_real = data_in_20_real;
  assign data_reorder_10_imag = data_in_20_imag;
  assign data_reorder_42_real = data_in_21_real;
  assign data_reorder_42_imag = data_in_21_imag;
  assign data_reorder_26_real = data_in_22_real;
  assign data_reorder_26_imag = data_in_22_imag;
  assign data_reorder_58_real = data_in_23_real;
  assign data_reorder_58_imag = data_in_23_imag;
  assign data_reorder_6_real = data_in_24_real;
  assign data_reorder_6_imag = data_in_24_imag;
  assign data_reorder_38_real = data_in_25_real;
  assign data_reorder_38_imag = data_in_25_imag;
  assign data_reorder_22_real = data_in_26_real;
  assign data_reorder_22_imag = data_in_26_imag;
  assign data_reorder_54_real = data_in_27_real;
  assign data_reorder_54_imag = data_in_27_imag;
  assign data_reorder_14_real = data_in_28_real;
  assign data_reorder_14_imag = data_in_28_imag;
  assign data_reorder_46_real = data_in_29_real;
  assign data_reorder_46_imag = data_in_29_imag;
  assign data_reorder_30_real = data_in_30_real;
  assign data_reorder_30_imag = data_in_30_imag;
  assign data_reorder_62_real = data_in_31_real;
  assign data_reorder_62_imag = data_in_31_imag;
  assign data_reorder_1_real = data_in_32_real;
  assign data_reorder_1_imag = data_in_32_imag;
  assign data_reorder_33_real = data_in_33_real;
  assign data_reorder_33_imag = data_in_33_imag;
  assign data_reorder_17_real = data_in_34_real;
  assign data_reorder_17_imag = data_in_34_imag;
  assign data_reorder_49_real = data_in_35_real;
  assign data_reorder_49_imag = data_in_35_imag;
  assign data_reorder_9_real = data_in_36_real;
  assign data_reorder_9_imag = data_in_36_imag;
  assign data_reorder_41_real = data_in_37_real;
  assign data_reorder_41_imag = data_in_37_imag;
  assign data_reorder_25_real = data_in_38_real;
  assign data_reorder_25_imag = data_in_38_imag;
  assign data_reorder_57_real = data_in_39_real;
  assign data_reorder_57_imag = data_in_39_imag;
  assign data_reorder_5_real = data_in_40_real;
  assign data_reorder_5_imag = data_in_40_imag;
  assign data_reorder_37_real = data_in_41_real;
  assign data_reorder_37_imag = data_in_41_imag;
  assign data_reorder_21_real = data_in_42_real;
  assign data_reorder_21_imag = data_in_42_imag;
  assign data_reorder_53_real = data_in_43_real;
  assign data_reorder_53_imag = data_in_43_imag;
  assign data_reorder_13_real = data_in_44_real;
  assign data_reorder_13_imag = data_in_44_imag;
  assign data_reorder_45_real = data_in_45_real;
  assign data_reorder_45_imag = data_in_45_imag;
  assign data_reorder_29_real = data_in_46_real;
  assign data_reorder_29_imag = data_in_46_imag;
  assign data_reorder_61_real = data_in_47_real;
  assign data_reorder_61_imag = data_in_47_imag;
  assign data_reorder_3_real = data_in_48_real;
  assign data_reorder_3_imag = data_in_48_imag;
  assign data_reorder_35_real = data_in_49_real;
  assign data_reorder_35_imag = data_in_49_imag;
  assign data_reorder_19_real = data_in_50_real;
  assign data_reorder_19_imag = data_in_50_imag;
  assign data_reorder_51_real = data_in_51_real;
  assign data_reorder_51_imag = data_in_51_imag;
  assign data_reorder_11_real = data_in_52_real;
  assign data_reorder_11_imag = data_in_52_imag;
  assign data_reorder_43_real = data_in_53_real;
  assign data_reorder_43_imag = data_in_53_imag;
  assign data_reorder_27_real = data_in_54_real;
  assign data_reorder_27_imag = data_in_54_imag;
  assign data_reorder_59_real = data_in_55_real;
  assign data_reorder_59_imag = data_in_55_imag;
  assign data_reorder_7_real = data_in_56_real;
  assign data_reorder_7_imag = data_in_56_imag;
  assign data_reorder_39_real = data_in_57_real;
  assign data_reorder_39_imag = data_in_57_imag;
  assign data_reorder_23_real = data_in_58_real;
  assign data_reorder_23_imag = data_in_58_imag;
  assign data_reorder_55_real = data_in_59_real;
  assign data_reorder_55_imag = data_in_59_imag;
  assign data_reorder_15_real = data_in_60_real;
  assign data_reorder_15_imag = data_in_60_imag;
  assign data_reorder_47_real = data_in_61_real;
  assign data_reorder_47_imag = data_in_61_imag;
  assign data_reorder_31_real = data_in_62_real;
  assign data_reorder_31_imag = data_in_62_imag;
  assign data_reorder_63_real = data_in_63_real;
  assign data_reorder_63_imag = data_in_63_imag;
  assign _zz_3 = ($signed(_zz_2113) * $signed(data_mid_0_1_real));
  assign _zz_961 = _zz_2114;
  assign _zz_1 = _zz_2117[35 : 0];
  assign _zz_962 = _zz_2118;
  assign _zz_2 = _zz_2121[35 : 0];
  assign _zz_4 = 1'b1;
  assign _zz_963 = _zz_2122;
  assign _zz_964 = _zz_2130;
  assign _zz_5 = 1'b1;
  assign _zz_965 = _zz_2138;
  assign _zz_966 = _zz_2146;
  assign _zz_8 = ($signed(_zz_2154) * $signed(data_mid_0_3_real));
  assign _zz_967 = _zz_2155;
  assign _zz_6 = _zz_2158[35 : 0];
  assign _zz_968 = _zz_2159;
  assign _zz_7 = _zz_2162[35 : 0];
  assign _zz_9 = 1'b1;
  assign _zz_969 = _zz_2163;
  assign _zz_970 = _zz_2171;
  assign _zz_10 = 1'b1;
  assign _zz_971 = _zz_2179;
  assign _zz_972 = _zz_2187;
  assign _zz_13 = ($signed(_zz_2195) * $signed(data_mid_0_5_real));
  assign _zz_973 = _zz_2196;
  assign _zz_11 = _zz_2199[35 : 0];
  assign _zz_974 = _zz_2200;
  assign _zz_12 = _zz_2203[35 : 0];
  assign _zz_14 = 1'b1;
  assign _zz_975 = _zz_2204;
  assign _zz_976 = _zz_2212;
  assign _zz_15 = 1'b1;
  assign _zz_977 = _zz_2220;
  assign _zz_978 = _zz_2228;
  assign _zz_18 = ($signed(_zz_2236) * $signed(data_mid_0_7_real));
  assign _zz_979 = _zz_2237;
  assign _zz_16 = _zz_2240[35 : 0];
  assign _zz_980 = _zz_2241;
  assign _zz_17 = _zz_2244[35 : 0];
  assign _zz_19 = 1'b1;
  assign _zz_981 = _zz_2245;
  assign _zz_982 = _zz_2253;
  assign _zz_20 = 1'b1;
  assign _zz_983 = _zz_2261;
  assign _zz_984 = _zz_2269;
  assign _zz_23 = ($signed(_zz_2277) * $signed(data_mid_0_9_real));
  assign _zz_985 = _zz_2278;
  assign _zz_21 = _zz_2281[35 : 0];
  assign _zz_986 = _zz_2282;
  assign _zz_22 = _zz_2285[35 : 0];
  assign _zz_24 = 1'b1;
  assign _zz_987 = _zz_2286;
  assign _zz_988 = _zz_2294;
  assign _zz_25 = 1'b1;
  assign _zz_989 = _zz_2302;
  assign _zz_990 = _zz_2310;
  assign _zz_28 = ($signed(_zz_2318) * $signed(data_mid_0_11_real));
  assign _zz_991 = _zz_2319;
  assign _zz_26 = _zz_2322[35 : 0];
  assign _zz_992 = _zz_2323;
  assign _zz_27 = _zz_2326[35 : 0];
  assign _zz_29 = 1'b1;
  assign _zz_993 = _zz_2327;
  assign _zz_994 = _zz_2335;
  assign _zz_30 = 1'b1;
  assign _zz_995 = _zz_2343;
  assign _zz_996 = _zz_2351;
  assign _zz_33 = ($signed(_zz_2359) * $signed(data_mid_0_13_real));
  assign _zz_997 = _zz_2360;
  assign _zz_31 = _zz_2363[35 : 0];
  assign _zz_998 = _zz_2364;
  assign _zz_32 = _zz_2367[35 : 0];
  assign _zz_34 = 1'b1;
  assign _zz_999 = _zz_2368;
  assign _zz_1000 = _zz_2376;
  assign _zz_35 = 1'b1;
  assign _zz_1001 = _zz_2384;
  assign _zz_1002 = _zz_2392;
  assign _zz_38 = ($signed(_zz_2400) * $signed(data_mid_0_15_real));
  assign _zz_1003 = _zz_2401;
  assign _zz_36 = _zz_2404[35 : 0];
  assign _zz_1004 = _zz_2405;
  assign _zz_37 = _zz_2408[35 : 0];
  assign _zz_39 = 1'b1;
  assign _zz_1005 = _zz_2409;
  assign _zz_1006 = _zz_2417;
  assign _zz_40 = 1'b1;
  assign _zz_1007 = _zz_2425;
  assign _zz_1008 = _zz_2433;
  assign _zz_43 = ($signed(_zz_2441) * $signed(data_mid_0_17_real));
  assign _zz_1009 = _zz_2442;
  assign _zz_41 = _zz_2445[35 : 0];
  assign _zz_1010 = _zz_2446;
  assign _zz_42 = _zz_2449[35 : 0];
  assign _zz_44 = 1'b1;
  assign _zz_1011 = _zz_2450;
  assign _zz_1012 = _zz_2458;
  assign _zz_45 = 1'b1;
  assign _zz_1013 = _zz_2466;
  assign _zz_1014 = _zz_2474;
  assign _zz_48 = ($signed(_zz_2482) * $signed(data_mid_0_19_real));
  assign _zz_1015 = _zz_2483;
  assign _zz_46 = _zz_2486[35 : 0];
  assign _zz_1016 = _zz_2487;
  assign _zz_47 = _zz_2490[35 : 0];
  assign _zz_49 = 1'b1;
  assign _zz_1017 = _zz_2491;
  assign _zz_1018 = _zz_2499;
  assign _zz_50 = 1'b1;
  assign _zz_1019 = _zz_2507;
  assign _zz_1020 = _zz_2515;
  assign _zz_53 = ($signed(_zz_2523) * $signed(data_mid_0_21_real));
  assign _zz_1021 = _zz_2524;
  assign _zz_51 = _zz_2527[35 : 0];
  assign _zz_1022 = _zz_2528;
  assign _zz_52 = _zz_2531[35 : 0];
  assign _zz_54 = 1'b1;
  assign _zz_1023 = _zz_2532;
  assign _zz_1024 = _zz_2540;
  assign _zz_55 = 1'b1;
  assign _zz_1025 = _zz_2548;
  assign _zz_1026 = _zz_2556;
  assign _zz_58 = ($signed(_zz_2564) * $signed(data_mid_0_23_real));
  assign _zz_1027 = _zz_2565;
  assign _zz_56 = _zz_2568[35 : 0];
  assign _zz_1028 = _zz_2569;
  assign _zz_57 = _zz_2572[35 : 0];
  assign _zz_59 = 1'b1;
  assign _zz_1029 = _zz_2573;
  assign _zz_1030 = _zz_2581;
  assign _zz_60 = 1'b1;
  assign _zz_1031 = _zz_2589;
  assign _zz_1032 = _zz_2597;
  assign _zz_63 = ($signed(_zz_2605) * $signed(data_mid_0_25_real));
  assign _zz_1033 = _zz_2606;
  assign _zz_61 = _zz_2609[35 : 0];
  assign _zz_1034 = _zz_2610;
  assign _zz_62 = _zz_2613[35 : 0];
  assign _zz_64 = 1'b1;
  assign _zz_1035 = _zz_2614;
  assign _zz_1036 = _zz_2622;
  assign _zz_65 = 1'b1;
  assign _zz_1037 = _zz_2630;
  assign _zz_1038 = _zz_2638;
  assign _zz_68 = ($signed(_zz_2646) * $signed(data_mid_0_27_real));
  assign _zz_1039 = _zz_2647;
  assign _zz_66 = _zz_2650[35 : 0];
  assign _zz_1040 = _zz_2651;
  assign _zz_67 = _zz_2654[35 : 0];
  assign _zz_69 = 1'b1;
  assign _zz_1041 = _zz_2655;
  assign _zz_1042 = _zz_2663;
  assign _zz_70 = 1'b1;
  assign _zz_1043 = _zz_2671;
  assign _zz_1044 = _zz_2679;
  assign _zz_73 = ($signed(_zz_2687) * $signed(data_mid_0_29_real));
  assign _zz_1045 = _zz_2688;
  assign _zz_71 = _zz_2691[35 : 0];
  assign _zz_1046 = _zz_2692;
  assign _zz_72 = _zz_2695[35 : 0];
  assign _zz_74 = 1'b1;
  assign _zz_1047 = _zz_2696;
  assign _zz_1048 = _zz_2704;
  assign _zz_75 = 1'b1;
  assign _zz_1049 = _zz_2712;
  assign _zz_1050 = _zz_2720;
  assign _zz_78 = ($signed(_zz_2728) * $signed(data_mid_0_31_real));
  assign _zz_1051 = _zz_2729;
  assign _zz_76 = _zz_2732[35 : 0];
  assign _zz_1052 = _zz_2733;
  assign _zz_77 = _zz_2736[35 : 0];
  assign _zz_79 = 1'b1;
  assign _zz_1053 = _zz_2737;
  assign _zz_1054 = _zz_2745;
  assign _zz_80 = 1'b1;
  assign _zz_1055 = _zz_2753;
  assign _zz_1056 = _zz_2761;
  assign _zz_83 = ($signed(_zz_2769) * $signed(data_mid_0_33_real));
  assign _zz_1057 = _zz_2770;
  assign _zz_81 = _zz_2773[35 : 0];
  assign _zz_1058 = _zz_2774;
  assign _zz_82 = _zz_2777[35 : 0];
  assign _zz_84 = 1'b1;
  assign _zz_1059 = _zz_2778;
  assign _zz_1060 = _zz_2786;
  assign _zz_85 = 1'b1;
  assign _zz_1061 = _zz_2794;
  assign _zz_1062 = _zz_2802;
  assign _zz_88 = ($signed(_zz_2810) * $signed(data_mid_0_35_real));
  assign _zz_1063 = _zz_2811;
  assign _zz_86 = _zz_2814[35 : 0];
  assign _zz_1064 = _zz_2815;
  assign _zz_87 = _zz_2818[35 : 0];
  assign _zz_89 = 1'b1;
  assign _zz_1065 = _zz_2819;
  assign _zz_1066 = _zz_2827;
  assign _zz_90 = 1'b1;
  assign _zz_1067 = _zz_2835;
  assign _zz_1068 = _zz_2843;
  assign _zz_93 = ($signed(_zz_2851) * $signed(data_mid_0_37_real));
  assign _zz_1069 = _zz_2852;
  assign _zz_91 = _zz_2855[35 : 0];
  assign _zz_1070 = _zz_2856;
  assign _zz_92 = _zz_2859[35 : 0];
  assign _zz_94 = 1'b1;
  assign _zz_1071 = _zz_2860;
  assign _zz_1072 = _zz_2868;
  assign _zz_95 = 1'b1;
  assign _zz_1073 = _zz_2876;
  assign _zz_1074 = _zz_2884;
  assign _zz_98 = ($signed(_zz_2892) * $signed(data_mid_0_39_real));
  assign _zz_1075 = _zz_2893;
  assign _zz_96 = _zz_2896[35 : 0];
  assign _zz_1076 = _zz_2897;
  assign _zz_97 = _zz_2900[35 : 0];
  assign _zz_99 = 1'b1;
  assign _zz_1077 = _zz_2901;
  assign _zz_1078 = _zz_2909;
  assign _zz_100 = 1'b1;
  assign _zz_1079 = _zz_2917;
  assign _zz_1080 = _zz_2925;
  assign _zz_103 = ($signed(_zz_2933) * $signed(data_mid_0_41_real));
  assign _zz_1081 = _zz_2934;
  assign _zz_101 = _zz_2937[35 : 0];
  assign _zz_1082 = _zz_2938;
  assign _zz_102 = _zz_2941[35 : 0];
  assign _zz_104 = 1'b1;
  assign _zz_1083 = _zz_2942;
  assign _zz_1084 = _zz_2950;
  assign _zz_105 = 1'b1;
  assign _zz_1085 = _zz_2958;
  assign _zz_1086 = _zz_2966;
  assign _zz_108 = ($signed(_zz_2974) * $signed(data_mid_0_43_real));
  assign _zz_1087 = _zz_2975;
  assign _zz_106 = _zz_2978[35 : 0];
  assign _zz_1088 = _zz_2979;
  assign _zz_107 = _zz_2982[35 : 0];
  assign _zz_109 = 1'b1;
  assign _zz_1089 = _zz_2983;
  assign _zz_1090 = _zz_2991;
  assign _zz_110 = 1'b1;
  assign _zz_1091 = _zz_2999;
  assign _zz_1092 = _zz_3007;
  assign _zz_113 = ($signed(_zz_3015) * $signed(data_mid_0_45_real));
  assign _zz_1093 = _zz_3016;
  assign _zz_111 = _zz_3019[35 : 0];
  assign _zz_1094 = _zz_3020;
  assign _zz_112 = _zz_3023[35 : 0];
  assign _zz_114 = 1'b1;
  assign _zz_1095 = _zz_3024;
  assign _zz_1096 = _zz_3032;
  assign _zz_115 = 1'b1;
  assign _zz_1097 = _zz_3040;
  assign _zz_1098 = _zz_3048;
  assign _zz_118 = ($signed(_zz_3056) * $signed(data_mid_0_47_real));
  assign _zz_1099 = _zz_3057;
  assign _zz_116 = _zz_3060[35 : 0];
  assign _zz_1100 = _zz_3061;
  assign _zz_117 = _zz_3064[35 : 0];
  assign _zz_119 = 1'b1;
  assign _zz_1101 = _zz_3065;
  assign _zz_1102 = _zz_3073;
  assign _zz_120 = 1'b1;
  assign _zz_1103 = _zz_3081;
  assign _zz_1104 = _zz_3089;
  assign _zz_123 = ($signed(_zz_3097) * $signed(data_mid_0_49_real));
  assign _zz_1105 = _zz_3098;
  assign _zz_121 = _zz_3101[35 : 0];
  assign _zz_1106 = _zz_3102;
  assign _zz_122 = _zz_3105[35 : 0];
  assign _zz_124 = 1'b1;
  assign _zz_1107 = _zz_3106;
  assign _zz_1108 = _zz_3114;
  assign _zz_125 = 1'b1;
  assign _zz_1109 = _zz_3122;
  assign _zz_1110 = _zz_3130;
  assign _zz_128 = ($signed(_zz_3138) * $signed(data_mid_0_51_real));
  assign _zz_1111 = _zz_3139;
  assign _zz_126 = _zz_3142[35 : 0];
  assign _zz_1112 = _zz_3143;
  assign _zz_127 = _zz_3146[35 : 0];
  assign _zz_129 = 1'b1;
  assign _zz_1113 = _zz_3147;
  assign _zz_1114 = _zz_3155;
  assign _zz_130 = 1'b1;
  assign _zz_1115 = _zz_3163;
  assign _zz_1116 = _zz_3171;
  assign _zz_133 = ($signed(_zz_3179) * $signed(data_mid_0_53_real));
  assign _zz_1117 = _zz_3180;
  assign _zz_131 = _zz_3183[35 : 0];
  assign _zz_1118 = _zz_3184;
  assign _zz_132 = _zz_3187[35 : 0];
  assign _zz_134 = 1'b1;
  assign _zz_1119 = _zz_3188;
  assign _zz_1120 = _zz_3196;
  assign _zz_135 = 1'b1;
  assign _zz_1121 = _zz_3204;
  assign _zz_1122 = _zz_3212;
  assign _zz_138 = ($signed(_zz_3220) * $signed(data_mid_0_55_real));
  assign _zz_1123 = _zz_3221;
  assign _zz_136 = _zz_3224[35 : 0];
  assign _zz_1124 = _zz_3225;
  assign _zz_137 = _zz_3228[35 : 0];
  assign _zz_139 = 1'b1;
  assign _zz_1125 = _zz_3229;
  assign _zz_1126 = _zz_3237;
  assign _zz_140 = 1'b1;
  assign _zz_1127 = _zz_3245;
  assign _zz_1128 = _zz_3253;
  assign _zz_143 = ($signed(_zz_3261) * $signed(data_mid_0_57_real));
  assign _zz_1129 = _zz_3262;
  assign _zz_141 = _zz_3265[35 : 0];
  assign _zz_1130 = _zz_3266;
  assign _zz_142 = _zz_3269[35 : 0];
  assign _zz_144 = 1'b1;
  assign _zz_1131 = _zz_3270;
  assign _zz_1132 = _zz_3278;
  assign _zz_145 = 1'b1;
  assign _zz_1133 = _zz_3286;
  assign _zz_1134 = _zz_3294;
  assign _zz_148 = ($signed(_zz_3302) * $signed(data_mid_0_59_real));
  assign _zz_1135 = _zz_3303;
  assign _zz_146 = _zz_3306[35 : 0];
  assign _zz_1136 = _zz_3307;
  assign _zz_147 = _zz_3310[35 : 0];
  assign _zz_149 = 1'b1;
  assign _zz_1137 = _zz_3311;
  assign _zz_1138 = _zz_3319;
  assign _zz_150 = 1'b1;
  assign _zz_1139 = _zz_3327;
  assign _zz_1140 = _zz_3335;
  assign _zz_153 = ($signed(_zz_3343) * $signed(data_mid_0_61_real));
  assign _zz_1141 = _zz_3344;
  assign _zz_151 = _zz_3347[35 : 0];
  assign _zz_1142 = _zz_3348;
  assign _zz_152 = _zz_3351[35 : 0];
  assign _zz_154 = 1'b1;
  assign _zz_1143 = _zz_3352;
  assign _zz_1144 = _zz_3360;
  assign _zz_155 = 1'b1;
  assign _zz_1145 = _zz_3368;
  assign _zz_1146 = _zz_3376;
  assign _zz_158 = ($signed(_zz_3384) * $signed(data_mid_0_63_real));
  assign _zz_1147 = _zz_3385;
  assign _zz_156 = _zz_3388[35 : 0];
  assign _zz_1148 = _zz_3389;
  assign _zz_157 = _zz_3392[35 : 0];
  assign _zz_159 = 1'b1;
  assign _zz_1149 = _zz_3393;
  assign _zz_1150 = _zz_3401;
  assign _zz_160 = 1'b1;
  assign _zz_1151 = _zz_3409;
  assign _zz_1152 = _zz_3417;
  assign _zz_163 = ($signed(_zz_3425) * $signed(data_mid_1_2_real));
  assign _zz_1153 = _zz_3426;
  assign _zz_161 = _zz_3429[35 : 0];
  assign _zz_1154 = _zz_3430;
  assign _zz_162 = _zz_3433[35 : 0];
  assign _zz_164 = 1'b1;
  assign _zz_1155 = _zz_3434;
  assign _zz_1156 = _zz_3442;
  assign _zz_165 = 1'b1;
  assign _zz_1157 = _zz_3450;
  assign _zz_1158 = _zz_3458;
  assign _zz_168 = ($signed(_zz_3466) * $signed(data_mid_1_3_real));
  assign _zz_1159 = _zz_3467;
  assign _zz_166 = _zz_3470[35 : 0];
  assign _zz_1160 = _zz_3471;
  assign _zz_167 = _zz_3474[35 : 0];
  assign _zz_169 = 1'b1;
  assign _zz_1161 = _zz_3475;
  assign _zz_1162 = _zz_3483;
  assign _zz_170 = 1'b1;
  assign _zz_1163 = _zz_3491;
  assign _zz_1164 = _zz_3499;
  assign _zz_173 = ($signed(_zz_3507) * $signed(data_mid_1_6_real));
  assign _zz_1165 = _zz_3508;
  assign _zz_171 = _zz_3511[35 : 0];
  assign _zz_1166 = _zz_3512;
  assign _zz_172 = _zz_3515[35 : 0];
  assign _zz_174 = 1'b1;
  assign _zz_1167 = _zz_3516;
  assign _zz_1168 = _zz_3524;
  assign _zz_175 = 1'b1;
  assign _zz_1169 = _zz_3532;
  assign _zz_1170 = _zz_3540;
  assign _zz_178 = ($signed(_zz_3548) * $signed(data_mid_1_7_real));
  assign _zz_1171 = _zz_3549;
  assign _zz_176 = _zz_3552[35 : 0];
  assign _zz_1172 = _zz_3553;
  assign _zz_177 = _zz_3556[35 : 0];
  assign _zz_179 = 1'b1;
  assign _zz_1173 = _zz_3557;
  assign _zz_1174 = _zz_3565;
  assign _zz_180 = 1'b1;
  assign _zz_1175 = _zz_3573;
  assign _zz_1176 = _zz_3581;
  assign _zz_183 = ($signed(_zz_3589) * $signed(data_mid_1_10_real));
  assign _zz_1177 = _zz_3590;
  assign _zz_181 = _zz_3593[35 : 0];
  assign _zz_1178 = _zz_3594;
  assign _zz_182 = _zz_3597[35 : 0];
  assign _zz_184 = 1'b1;
  assign _zz_1179 = _zz_3598;
  assign _zz_1180 = _zz_3606;
  assign _zz_185 = 1'b1;
  assign _zz_1181 = _zz_3614;
  assign _zz_1182 = _zz_3622;
  assign _zz_188 = ($signed(_zz_3630) * $signed(data_mid_1_11_real));
  assign _zz_1183 = _zz_3631;
  assign _zz_186 = _zz_3634[35 : 0];
  assign _zz_1184 = _zz_3635;
  assign _zz_187 = _zz_3638[35 : 0];
  assign _zz_189 = 1'b1;
  assign _zz_1185 = _zz_3639;
  assign _zz_1186 = _zz_3647;
  assign _zz_190 = 1'b1;
  assign _zz_1187 = _zz_3655;
  assign _zz_1188 = _zz_3663;
  assign _zz_193 = ($signed(_zz_3671) * $signed(data_mid_1_14_real));
  assign _zz_1189 = _zz_3672;
  assign _zz_191 = _zz_3675[35 : 0];
  assign _zz_1190 = _zz_3676;
  assign _zz_192 = _zz_3679[35 : 0];
  assign _zz_194 = 1'b1;
  assign _zz_1191 = _zz_3680;
  assign _zz_1192 = _zz_3688;
  assign _zz_195 = 1'b1;
  assign _zz_1193 = _zz_3696;
  assign _zz_1194 = _zz_3704;
  assign _zz_198 = ($signed(_zz_3712) * $signed(data_mid_1_15_real));
  assign _zz_1195 = _zz_3713;
  assign _zz_196 = _zz_3716[35 : 0];
  assign _zz_1196 = _zz_3717;
  assign _zz_197 = _zz_3720[35 : 0];
  assign _zz_199 = 1'b1;
  assign _zz_1197 = _zz_3721;
  assign _zz_1198 = _zz_3729;
  assign _zz_200 = 1'b1;
  assign _zz_1199 = _zz_3737;
  assign _zz_1200 = _zz_3745;
  assign _zz_203 = ($signed(_zz_3753) * $signed(data_mid_1_18_real));
  assign _zz_1201 = _zz_3754;
  assign _zz_201 = _zz_3757[35 : 0];
  assign _zz_1202 = _zz_3758;
  assign _zz_202 = _zz_3761[35 : 0];
  assign _zz_204 = 1'b1;
  assign _zz_1203 = _zz_3762;
  assign _zz_1204 = _zz_3770;
  assign _zz_205 = 1'b1;
  assign _zz_1205 = _zz_3778;
  assign _zz_1206 = _zz_3786;
  assign _zz_208 = ($signed(_zz_3794) * $signed(data_mid_1_19_real));
  assign _zz_1207 = _zz_3795;
  assign _zz_206 = _zz_3798[35 : 0];
  assign _zz_1208 = _zz_3799;
  assign _zz_207 = _zz_3802[35 : 0];
  assign _zz_209 = 1'b1;
  assign _zz_1209 = _zz_3803;
  assign _zz_1210 = _zz_3811;
  assign _zz_210 = 1'b1;
  assign _zz_1211 = _zz_3819;
  assign _zz_1212 = _zz_3827;
  assign _zz_213 = ($signed(_zz_3835) * $signed(data_mid_1_22_real));
  assign _zz_1213 = _zz_3836;
  assign _zz_211 = _zz_3839[35 : 0];
  assign _zz_1214 = _zz_3840;
  assign _zz_212 = _zz_3843[35 : 0];
  assign _zz_214 = 1'b1;
  assign _zz_1215 = _zz_3844;
  assign _zz_1216 = _zz_3852;
  assign _zz_215 = 1'b1;
  assign _zz_1217 = _zz_3860;
  assign _zz_1218 = _zz_3868;
  assign _zz_218 = ($signed(_zz_3876) * $signed(data_mid_1_23_real));
  assign _zz_1219 = _zz_3877;
  assign _zz_216 = _zz_3880[35 : 0];
  assign _zz_1220 = _zz_3881;
  assign _zz_217 = _zz_3884[35 : 0];
  assign _zz_219 = 1'b1;
  assign _zz_1221 = _zz_3885;
  assign _zz_1222 = _zz_3893;
  assign _zz_220 = 1'b1;
  assign _zz_1223 = _zz_3901;
  assign _zz_1224 = _zz_3909;
  assign _zz_223 = ($signed(_zz_3917) * $signed(data_mid_1_26_real));
  assign _zz_1225 = _zz_3918;
  assign _zz_221 = _zz_3921[35 : 0];
  assign _zz_1226 = _zz_3922;
  assign _zz_222 = _zz_3925[35 : 0];
  assign _zz_224 = 1'b1;
  assign _zz_1227 = _zz_3926;
  assign _zz_1228 = _zz_3934;
  assign _zz_225 = 1'b1;
  assign _zz_1229 = _zz_3942;
  assign _zz_1230 = _zz_3950;
  assign _zz_228 = ($signed(_zz_3958) * $signed(data_mid_1_27_real));
  assign _zz_1231 = _zz_3959;
  assign _zz_226 = _zz_3962[35 : 0];
  assign _zz_1232 = _zz_3963;
  assign _zz_227 = _zz_3966[35 : 0];
  assign _zz_229 = 1'b1;
  assign _zz_1233 = _zz_3967;
  assign _zz_1234 = _zz_3975;
  assign _zz_230 = 1'b1;
  assign _zz_1235 = _zz_3983;
  assign _zz_1236 = _zz_3991;
  assign _zz_233 = ($signed(_zz_3999) * $signed(data_mid_1_30_real));
  assign _zz_1237 = _zz_4000;
  assign _zz_231 = _zz_4003[35 : 0];
  assign _zz_1238 = _zz_4004;
  assign _zz_232 = _zz_4007[35 : 0];
  assign _zz_234 = 1'b1;
  assign _zz_1239 = _zz_4008;
  assign _zz_1240 = _zz_4016;
  assign _zz_235 = 1'b1;
  assign _zz_1241 = _zz_4024;
  assign _zz_1242 = _zz_4032;
  assign _zz_238 = ($signed(_zz_4040) * $signed(data_mid_1_31_real));
  assign _zz_1243 = _zz_4041;
  assign _zz_236 = _zz_4044[35 : 0];
  assign _zz_1244 = _zz_4045;
  assign _zz_237 = _zz_4048[35 : 0];
  assign _zz_239 = 1'b1;
  assign _zz_1245 = _zz_4049;
  assign _zz_1246 = _zz_4057;
  assign _zz_240 = 1'b1;
  assign _zz_1247 = _zz_4065;
  assign _zz_1248 = _zz_4073;
  assign _zz_243 = ($signed(_zz_4081) * $signed(data_mid_1_34_real));
  assign _zz_1249 = _zz_4082;
  assign _zz_241 = _zz_4085[35 : 0];
  assign _zz_1250 = _zz_4086;
  assign _zz_242 = _zz_4089[35 : 0];
  assign _zz_244 = 1'b1;
  assign _zz_1251 = _zz_4090;
  assign _zz_1252 = _zz_4098;
  assign _zz_245 = 1'b1;
  assign _zz_1253 = _zz_4106;
  assign _zz_1254 = _zz_4114;
  assign _zz_248 = ($signed(_zz_4122) * $signed(data_mid_1_35_real));
  assign _zz_1255 = _zz_4123;
  assign _zz_246 = _zz_4126[35 : 0];
  assign _zz_1256 = _zz_4127;
  assign _zz_247 = _zz_4130[35 : 0];
  assign _zz_249 = 1'b1;
  assign _zz_1257 = _zz_4131;
  assign _zz_1258 = _zz_4139;
  assign _zz_250 = 1'b1;
  assign _zz_1259 = _zz_4147;
  assign _zz_1260 = _zz_4155;
  assign _zz_253 = ($signed(_zz_4163) * $signed(data_mid_1_38_real));
  assign _zz_1261 = _zz_4164;
  assign _zz_251 = _zz_4167[35 : 0];
  assign _zz_1262 = _zz_4168;
  assign _zz_252 = _zz_4171[35 : 0];
  assign _zz_254 = 1'b1;
  assign _zz_1263 = _zz_4172;
  assign _zz_1264 = _zz_4180;
  assign _zz_255 = 1'b1;
  assign _zz_1265 = _zz_4188;
  assign _zz_1266 = _zz_4196;
  assign _zz_258 = ($signed(_zz_4204) * $signed(data_mid_1_39_real));
  assign _zz_1267 = _zz_4205;
  assign _zz_256 = _zz_4208[35 : 0];
  assign _zz_1268 = _zz_4209;
  assign _zz_257 = _zz_4212[35 : 0];
  assign _zz_259 = 1'b1;
  assign _zz_1269 = _zz_4213;
  assign _zz_1270 = _zz_4221;
  assign _zz_260 = 1'b1;
  assign _zz_1271 = _zz_4229;
  assign _zz_1272 = _zz_4237;
  assign _zz_263 = ($signed(_zz_4245) * $signed(data_mid_1_42_real));
  assign _zz_1273 = _zz_4246;
  assign _zz_261 = _zz_4249[35 : 0];
  assign _zz_1274 = _zz_4250;
  assign _zz_262 = _zz_4253[35 : 0];
  assign _zz_264 = 1'b1;
  assign _zz_1275 = _zz_4254;
  assign _zz_1276 = _zz_4262;
  assign _zz_265 = 1'b1;
  assign _zz_1277 = _zz_4270;
  assign _zz_1278 = _zz_4278;
  assign _zz_268 = ($signed(_zz_4286) * $signed(data_mid_1_43_real));
  assign _zz_1279 = _zz_4287;
  assign _zz_266 = _zz_4290[35 : 0];
  assign _zz_1280 = _zz_4291;
  assign _zz_267 = _zz_4294[35 : 0];
  assign _zz_269 = 1'b1;
  assign _zz_1281 = _zz_4295;
  assign _zz_1282 = _zz_4303;
  assign _zz_270 = 1'b1;
  assign _zz_1283 = _zz_4311;
  assign _zz_1284 = _zz_4319;
  assign _zz_273 = ($signed(_zz_4327) * $signed(data_mid_1_46_real));
  assign _zz_1285 = _zz_4328;
  assign _zz_271 = _zz_4331[35 : 0];
  assign _zz_1286 = _zz_4332;
  assign _zz_272 = _zz_4335[35 : 0];
  assign _zz_274 = 1'b1;
  assign _zz_1287 = _zz_4336;
  assign _zz_1288 = _zz_4344;
  assign _zz_275 = 1'b1;
  assign _zz_1289 = _zz_4352;
  assign _zz_1290 = _zz_4360;
  assign _zz_278 = ($signed(_zz_4368) * $signed(data_mid_1_47_real));
  assign _zz_1291 = _zz_4369;
  assign _zz_276 = _zz_4372[35 : 0];
  assign _zz_1292 = _zz_4373;
  assign _zz_277 = _zz_4376[35 : 0];
  assign _zz_279 = 1'b1;
  assign _zz_1293 = _zz_4377;
  assign _zz_1294 = _zz_4385;
  assign _zz_280 = 1'b1;
  assign _zz_1295 = _zz_4393;
  assign _zz_1296 = _zz_4401;
  assign _zz_283 = ($signed(_zz_4409) * $signed(data_mid_1_50_real));
  assign _zz_1297 = _zz_4410;
  assign _zz_281 = _zz_4413[35 : 0];
  assign _zz_1298 = _zz_4414;
  assign _zz_282 = _zz_4417[35 : 0];
  assign _zz_284 = 1'b1;
  assign _zz_1299 = _zz_4418;
  assign _zz_1300 = _zz_4426;
  assign _zz_285 = 1'b1;
  assign _zz_1301 = _zz_4434;
  assign _zz_1302 = _zz_4442;
  assign _zz_288 = ($signed(_zz_4450) * $signed(data_mid_1_51_real));
  assign _zz_1303 = _zz_4451;
  assign _zz_286 = _zz_4454[35 : 0];
  assign _zz_1304 = _zz_4455;
  assign _zz_287 = _zz_4458[35 : 0];
  assign _zz_289 = 1'b1;
  assign _zz_1305 = _zz_4459;
  assign _zz_1306 = _zz_4467;
  assign _zz_290 = 1'b1;
  assign _zz_1307 = _zz_4475;
  assign _zz_1308 = _zz_4483;
  assign _zz_293 = ($signed(_zz_4491) * $signed(data_mid_1_54_real));
  assign _zz_1309 = _zz_4492;
  assign _zz_291 = _zz_4495[35 : 0];
  assign _zz_1310 = _zz_4496;
  assign _zz_292 = _zz_4499[35 : 0];
  assign _zz_294 = 1'b1;
  assign _zz_1311 = _zz_4500;
  assign _zz_1312 = _zz_4508;
  assign _zz_295 = 1'b1;
  assign _zz_1313 = _zz_4516;
  assign _zz_1314 = _zz_4524;
  assign _zz_298 = ($signed(_zz_4532) * $signed(data_mid_1_55_real));
  assign _zz_1315 = _zz_4533;
  assign _zz_296 = _zz_4536[35 : 0];
  assign _zz_1316 = _zz_4537;
  assign _zz_297 = _zz_4540[35 : 0];
  assign _zz_299 = 1'b1;
  assign _zz_1317 = _zz_4541;
  assign _zz_1318 = _zz_4549;
  assign _zz_300 = 1'b1;
  assign _zz_1319 = _zz_4557;
  assign _zz_1320 = _zz_4565;
  assign _zz_303 = ($signed(_zz_4573) * $signed(data_mid_1_58_real));
  assign _zz_1321 = _zz_4574;
  assign _zz_301 = _zz_4577[35 : 0];
  assign _zz_1322 = _zz_4578;
  assign _zz_302 = _zz_4581[35 : 0];
  assign _zz_304 = 1'b1;
  assign _zz_1323 = _zz_4582;
  assign _zz_1324 = _zz_4590;
  assign _zz_305 = 1'b1;
  assign _zz_1325 = _zz_4598;
  assign _zz_1326 = _zz_4606;
  assign _zz_308 = ($signed(_zz_4614) * $signed(data_mid_1_59_real));
  assign _zz_1327 = _zz_4615;
  assign _zz_306 = _zz_4618[35 : 0];
  assign _zz_1328 = _zz_4619;
  assign _zz_307 = _zz_4622[35 : 0];
  assign _zz_309 = 1'b1;
  assign _zz_1329 = _zz_4623;
  assign _zz_1330 = _zz_4631;
  assign _zz_310 = 1'b1;
  assign _zz_1331 = _zz_4639;
  assign _zz_1332 = _zz_4647;
  assign _zz_313 = ($signed(_zz_4655) * $signed(data_mid_1_62_real));
  assign _zz_1333 = _zz_4656;
  assign _zz_311 = _zz_4659[35 : 0];
  assign _zz_1334 = _zz_4660;
  assign _zz_312 = _zz_4663[35 : 0];
  assign _zz_314 = 1'b1;
  assign _zz_1335 = _zz_4664;
  assign _zz_1336 = _zz_4672;
  assign _zz_315 = 1'b1;
  assign _zz_1337 = _zz_4680;
  assign _zz_1338 = _zz_4688;
  assign _zz_318 = ($signed(_zz_4696) * $signed(data_mid_1_63_real));
  assign _zz_1339 = _zz_4697;
  assign _zz_316 = _zz_4700[35 : 0];
  assign _zz_1340 = _zz_4701;
  assign _zz_317 = _zz_4704[35 : 0];
  assign _zz_319 = 1'b1;
  assign _zz_1341 = _zz_4705;
  assign _zz_1342 = _zz_4713;
  assign _zz_320 = 1'b1;
  assign _zz_1343 = _zz_4721;
  assign _zz_1344 = _zz_4729;
  assign _zz_323 = ($signed(_zz_4737) * $signed(data_mid_2_4_real));
  assign _zz_1345 = _zz_4738;
  assign _zz_321 = _zz_4741[35 : 0];
  assign _zz_1346 = _zz_4742;
  assign _zz_322 = _zz_4745[35 : 0];
  assign _zz_324 = 1'b1;
  assign _zz_1347 = _zz_4746;
  assign _zz_1348 = _zz_4754;
  assign _zz_325 = 1'b1;
  assign _zz_1349 = _zz_4762;
  assign _zz_1350 = _zz_4770;
  assign _zz_328 = ($signed(_zz_4778) * $signed(data_mid_2_5_real));
  assign _zz_1351 = _zz_4779;
  assign _zz_326 = _zz_4782[35 : 0];
  assign _zz_1352 = _zz_4783;
  assign _zz_327 = _zz_4786[35 : 0];
  assign _zz_329 = 1'b1;
  assign _zz_1353 = _zz_4787;
  assign _zz_1354 = _zz_4795;
  assign _zz_330 = 1'b1;
  assign _zz_1355 = _zz_4803;
  assign _zz_1356 = _zz_4811;
  assign _zz_333 = ($signed(_zz_4819) * $signed(data_mid_2_6_real));
  assign _zz_1357 = _zz_4820;
  assign _zz_331 = _zz_4823[35 : 0];
  assign _zz_1358 = _zz_4824;
  assign _zz_332 = _zz_4827[35 : 0];
  assign _zz_334 = 1'b1;
  assign _zz_1359 = _zz_4828;
  assign _zz_1360 = _zz_4836;
  assign _zz_335 = 1'b1;
  assign _zz_1361 = _zz_4844;
  assign _zz_1362 = _zz_4852;
  assign _zz_338 = ($signed(_zz_4860) * $signed(data_mid_2_7_real));
  assign _zz_1363 = _zz_4861;
  assign _zz_336 = _zz_4864[35 : 0];
  assign _zz_1364 = _zz_4865;
  assign _zz_337 = _zz_4868[35 : 0];
  assign _zz_339 = 1'b1;
  assign _zz_1365 = _zz_4869;
  assign _zz_1366 = _zz_4877;
  assign _zz_340 = 1'b1;
  assign _zz_1367 = _zz_4885;
  assign _zz_1368 = _zz_4893;
  assign _zz_343 = ($signed(_zz_4901) * $signed(data_mid_2_12_real));
  assign _zz_1369 = _zz_4902;
  assign _zz_341 = _zz_4905[35 : 0];
  assign _zz_1370 = _zz_4906;
  assign _zz_342 = _zz_4909[35 : 0];
  assign _zz_344 = 1'b1;
  assign _zz_1371 = _zz_4910;
  assign _zz_1372 = _zz_4918;
  assign _zz_345 = 1'b1;
  assign _zz_1373 = _zz_4926;
  assign _zz_1374 = _zz_4934;
  assign _zz_348 = ($signed(_zz_4942) * $signed(data_mid_2_13_real));
  assign _zz_1375 = _zz_4943;
  assign _zz_346 = _zz_4946[35 : 0];
  assign _zz_1376 = _zz_4947;
  assign _zz_347 = _zz_4950[35 : 0];
  assign _zz_349 = 1'b1;
  assign _zz_1377 = _zz_4951;
  assign _zz_1378 = _zz_4959;
  assign _zz_350 = 1'b1;
  assign _zz_1379 = _zz_4967;
  assign _zz_1380 = _zz_4975;
  assign _zz_353 = ($signed(_zz_4983) * $signed(data_mid_2_14_real));
  assign _zz_1381 = _zz_4984;
  assign _zz_351 = _zz_4987[35 : 0];
  assign _zz_1382 = _zz_4988;
  assign _zz_352 = _zz_4991[35 : 0];
  assign _zz_354 = 1'b1;
  assign _zz_1383 = _zz_4992;
  assign _zz_1384 = _zz_5000;
  assign _zz_355 = 1'b1;
  assign _zz_1385 = _zz_5008;
  assign _zz_1386 = _zz_5016;
  assign _zz_358 = ($signed(_zz_5024) * $signed(data_mid_2_15_real));
  assign _zz_1387 = _zz_5025;
  assign _zz_356 = _zz_5028[35 : 0];
  assign _zz_1388 = _zz_5029;
  assign _zz_357 = _zz_5032[35 : 0];
  assign _zz_359 = 1'b1;
  assign _zz_1389 = _zz_5033;
  assign _zz_1390 = _zz_5041;
  assign _zz_360 = 1'b1;
  assign _zz_1391 = _zz_5049;
  assign _zz_1392 = _zz_5057;
  assign _zz_363 = ($signed(_zz_5065) * $signed(data_mid_2_20_real));
  assign _zz_1393 = _zz_5066;
  assign _zz_361 = _zz_5069[35 : 0];
  assign _zz_1394 = _zz_5070;
  assign _zz_362 = _zz_5073[35 : 0];
  assign _zz_364 = 1'b1;
  assign _zz_1395 = _zz_5074;
  assign _zz_1396 = _zz_5082;
  assign _zz_365 = 1'b1;
  assign _zz_1397 = _zz_5090;
  assign _zz_1398 = _zz_5098;
  assign _zz_368 = ($signed(_zz_5106) * $signed(data_mid_2_21_real));
  assign _zz_1399 = _zz_5107;
  assign _zz_366 = _zz_5110[35 : 0];
  assign _zz_1400 = _zz_5111;
  assign _zz_367 = _zz_5114[35 : 0];
  assign _zz_369 = 1'b1;
  assign _zz_1401 = _zz_5115;
  assign _zz_1402 = _zz_5123;
  assign _zz_370 = 1'b1;
  assign _zz_1403 = _zz_5131;
  assign _zz_1404 = _zz_5139;
  assign _zz_373 = ($signed(_zz_5147) * $signed(data_mid_2_22_real));
  assign _zz_1405 = _zz_5148;
  assign _zz_371 = _zz_5151[35 : 0];
  assign _zz_1406 = _zz_5152;
  assign _zz_372 = _zz_5155[35 : 0];
  assign _zz_374 = 1'b1;
  assign _zz_1407 = _zz_5156;
  assign _zz_1408 = _zz_5164;
  assign _zz_375 = 1'b1;
  assign _zz_1409 = _zz_5172;
  assign _zz_1410 = _zz_5180;
  assign _zz_378 = ($signed(_zz_5188) * $signed(data_mid_2_23_real));
  assign _zz_1411 = _zz_5189;
  assign _zz_376 = _zz_5192[35 : 0];
  assign _zz_1412 = _zz_5193;
  assign _zz_377 = _zz_5196[35 : 0];
  assign _zz_379 = 1'b1;
  assign _zz_1413 = _zz_5197;
  assign _zz_1414 = _zz_5205;
  assign _zz_380 = 1'b1;
  assign _zz_1415 = _zz_5213;
  assign _zz_1416 = _zz_5221;
  assign _zz_383 = ($signed(_zz_5229) * $signed(data_mid_2_28_real));
  assign _zz_1417 = _zz_5230;
  assign _zz_381 = _zz_5233[35 : 0];
  assign _zz_1418 = _zz_5234;
  assign _zz_382 = _zz_5237[35 : 0];
  assign _zz_384 = 1'b1;
  assign _zz_1419 = _zz_5238;
  assign _zz_1420 = _zz_5246;
  assign _zz_385 = 1'b1;
  assign _zz_1421 = _zz_5254;
  assign _zz_1422 = _zz_5262;
  assign _zz_388 = ($signed(_zz_5270) * $signed(data_mid_2_29_real));
  assign _zz_1423 = _zz_5271;
  assign _zz_386 = _zz_5274[35 : 0];
  assign _zz_1424 = _zz_5275;
  assign _zz_387 = _zz_5278[35 : 0];
  assign _zz_389 = 1'b1;
  assign _zz_1425 = _zz_5279;
  assign _zz_1426 = _zz_5287;
  assign _zz_390 = 1'b1;
  assign _zz_1427 = _zz_5295;
  assign _zz_1428 = _zz_5303;
  assign _zz_393 = ($signed(_zz_5311) * $signed(data_mid_2_30_real));
  assign _zz_1429 = _zz_5312;
  assign _zz_391 = _zz_5315[35 : 0];
  assign _zz_1430 = _zz_5316;
  assign _zz_392 = _zz_5319[35 : 0];
  assign _zz_394 = 1'b1;
  assign _zz_1431 = _zz_5320;
  assign _zz_1432 = _zz_5328;
  assign _zz_395 = 1'b1;
  assign _zz_1433 = _zz_5336;
  assign _zz_1434 = _zz_5344;
  assign _zz_398 = ($signed(_zz_5352) * $signed(data_mid_2_31_real));
  assign _zz_1435 = _zz_5353;
  assign _zz_396 = _zz_5356[35 : 0];
  assign _zz_1436 = _zz_5357;
  assign _zz_397 = _zz_5360[35 : 0];
  assign _zz_399 = 1'b1;
  assign _zz_1437 = _zz_5361;
  assign _zz_1438 = _zz_5369;
  assign _zz_400 = 1'b1;
  assign _zz_1439 = _zz_5377;
  assign _zz_1440 = _zz_5385;
  assign _zz_403 = ($signed(_zz_5393) * $signed(data_mid_2_36_real));
  assign _zz_1441 = _zz_5394;
  assign _zz_401 = _zz_5397[35 : 0];
  assign _zz_1442 = _zz_5398;
  assign _zz_402 = _zz_5401[35 : 0];
  assign _zz_404 = 1'b1;
  assign _zz_1443 = _zz_5402;
  assign _zz_1444 = _zz_5410;
  assign _zz_405 = 1'b1;
  assign _zz_1445 = _zz_5418;
  assign _zz_1446 = _zz_5426;
  assign _zz_408 = ($signed(_zz_5434) * $signed(data_mid_2_37_real));
  assign _zz_1447 = _zz_5435;
  assign _zz_406 = _zz_5438[35 : 0];
  assign _zz_1448 = _zz_5439;
  assign _zz_407 = _zz_5442[35 : 0];
  assign _zz_409 = 1'b1;
  assign _zz_1449 = _zz_5443;
  assign _zz_1450 = _zz_5451;
  assign _zz_410 = 1'b1;
  assign _zz_1451 = _zz_5459;
  assign _zz_1452 = _zz_5467;
  assign _zz_413 = ($signed(_zz_5475) * $signed(data_mid_2_38_real));
  assign _zz_1453 = _zz_5476;
  assign _zz_411 = _zz_5479[35 : 0];
  assign _zz_1454 = _zz_5480;
  assign _zz_412 = _zz_5483[35 : 0];
  assign _zz_414 = 1'b1;
  assign _zz_1455 = _zz_5484;
  assign _zz_1456 = _zz_5492;
  assign _zz_415 = 1'b1;
  assign _zz_1457 = _zz_5500;
  assign _zz_1458 = _zz_5508;
  assign _zz_418 = ($signed(_zz_5516) * $signed(data_mid_2_39_real));
  assign _zz_1459 = _zz_5517;
  assign _zz_416 = _zz_5520[35 : 0];
  assign _zz_1460 = _zz_5521;
  assign _zz_417 = _zz_5524[35 : 0];
  assign _zz_419 = 1'b1;
  assign _zz_1461 = _zz_5525;
  assign _zz_1462 = _zz_5533;
  assign _zz_420 = 1'b1;
  assign _zz_1463 = _zz_5541;
  assign _zz_1464 = _zz_5549;
  assign _zz_423 = ($signed(_zz_5557) * $signed(data_mid_2_44_real));
  assign _zz_1465 = _zz_5558;
  assign _zz_421 = _zz_5561[35 : 0];
  assign _zz_1466 = _zz_5562;
  assign _zz_422 = _zz_5565[35 : 0];
  assign _zz_424 = 1'b1;
  assign _zz_1467 = _zz_5566;
  assign _zz_1468 = _zz_5574;
  assign _zz_425 = 1'b1;
  assign _zz_1469 = _zz_5582;
  assign _zz_1470 = _zz_5590;
  assign _zz_428 = ($signed(_zz_5598) * $signed(data_mid_2_45_real));
  assign _zz_1471 = _zz_5599;
  assign _zz_426 = _zz_5602[35 : 0];
  assign _zz_1472 = _zz_5603;
  assign _zz_427 = _zz_5606[35 : 0];
  assign _zz_429 = 1'b1;
  assign _zz_1473 = _zz_5607;
  assign _zz_1474 = _zz_5615;
  assign _zz_430 = 1'b1;
  assign _zz_1475 = _zz_5623;
  assign _zz_1476 = _zz_5631;
  assign _zz_433 = ($signed(_zz_5639) * $signed(data_mid_2_46_real));
  assign _zz_1477 = _zz_5640;
  assign _zz_431 = _zz_5643[35 : 0];
  assign _zz_1478 = _zz_5644;
  assign _zz_432 = _zz_5647[35 : 0];
  assign _zz_434 = 1'b1;
  assign _zz_1479 = _zz_5648;
  assign _zz_1480 = _zz_5656;
  assign _zz_435 = 1'b1;
  assign _zz_1481 = _zz_5664;
  assign _zz_1482 = _zz_5672;
  assign _zz_438 = ($signed(_zz_5680) * $signed(data_mid_2_47_real));
  assign _zz_1483 = _zz_5681;
  assign _zz_436 = _zz_5684[35 : 0];
  assign _zz_1484 = _zz_5685;
  assign _zz_437 = _zz_5688[35 : 0];
  assign _zz_439 = 1'b1;
  assign _zz_1485 = _zz_5689;
  assign _zz_1486 = _zz_5697;
  assign _zz_440 = 1'b1;
  assign _zz_1487 = _zz_5705;
  assign _zz_1488 = _zz_5713;
  assign _zz_443 = ($signed(_zz_5721) * $signed(data_mid_2_52_real));
  assign _zz_1489 = _zz_5722;
  assign _zz_441 = _zz_5725[35 : 0];
  assign _zz_1490 = _zz_5726;
  assign _zz_442 = _zz_5729[35 : 0];
  assign _zz_444 = 1'b1;
  assign _zz_1491 = _zz_5730;
  assign _zz_1492 = _zz_5738;
  assign _zz_445 = 1'b1;
  assign _zz_1493 = _zz_5746;
  assign _zz_1494 = _zz_5754;
  assign _zz_448 = ($signed(_zz_5762) * $signed(data_mid_2_53_real));
  assign _zz_1495 = _zz_5763;
  assign _zz_446 = _zz_5766[35 : 0];
  assign _zz_1496 = _zz_5767;
  assign _zz_447 = _zz_5770[35 : 0];
  assign _zz_449 = 1'b1;
  assign _zz_1497 = _zz_5771;
  assign _zz_1498 = _zz_5779;
  assign _zz_450 = 1'b1;
  assign _zz_1499 = _zz_5787;
  assign _zz_1500 = _zz_5795;
  assign _zz_453 = ($signed(_zz_5803) * $signed(data_mid_2_54_real));
  assign _zz_1501 = _zz_5804;
  assign _zz_451 = _zz_5807[35 : 0];
  assign _zz_1502 = _zz_5808;
  assign _zz_452 = _zz_5811[35 : 0];
  assign _zz_454 = 1'b1;
  assign _zz_1503 = _zz_5812;
  assign _zz_1504 = _zz_5820;
  assign _zz_455 = 1'b1;
  assign _zz_1505 = _zz_5828;
  assign _zz_1506 = _zz_5836;
  assign _zz_458 = ($signed(_zz_5844) * $signed(data_mid_2_55_real));
  assign _zz_1507 = _zz_5845;
  assign _zz_456 = _zz_5848[35 : 0];
  assign _zz_1508 = _zz_5849;
  assign _zz_457 = _zz_5852[35 : 0];
  assign _zz_459 = 1'b1;
  assign _zz_1509 = _zz_5853;
  assign _zz_1510 = _zz_5861;
  assign _zz_460 = 1'b1;
  assign _zz_1511 = _zz_5869;
  assign _zz_1512 = _zz_5877;
  assign _zz_463 = ($signed(_zz_5885) * $signed(data_mid_2_60_real));
  assign _zz_1513 = _zz_5886;
  assign _zz_461 = _zz_5889[35 : 0];
  assign _zz_1514 = _zz_5890;
  assign _zz_462 = _zz_5893[35 : 0];
  assign _zz_464 = 1'b1;
  assign _zz_1515 = _zz_5894;
  assign _zz_1516 = _zz_5902;
  assign _zz_465 = 1'b1;
  assign _zz_1517 = _zz_5910;
  assign _zz_1518 = _zz_5918;
  assign _zz_468 = ($signed(_zz_5926) * $signed(data_mid_2_61_real));
  assign _zz_1519 = _zz_5927;
  assign _zz_466 = _zz_5930[35 : 0];
  assign _zz_1520 = _zz_5931;
  assign _zz_467 = _zz_5934[35 : 0];
  assign _zz_469 = 1'b1;
  assign _zz_1521 = _zz_5935;
  assign _zz_1522 = _zz_5943;
  assign _zz_470 = 1'b1;
  assign _zz_1523 = _zz_5951;
  assign _zz_1524 = _zz_5959;
  assign _zz_473 = ($signed(_zz_5967) * $signed(data_mid_2_62_real));
  assign _zz_1525 = _zz_5968;
  assign _zz_471 = _zz_5971[35 : 0];
  assign _zz_1526 = _zz_5972;
  assign _zz_472 = _zz_5975[35 : 0];
  assign _zz_474 = 1'b1;
  assign _zz_1527 = _zz_5976;
  assign _zz_1528 = _zz_5984;
  assign _zz_475 = 1'b1;
  assign _zz_1529 = _zz_5992;
  assign _zz_1530 = _zz_6000;
  assign _zz_478 = ($signed(_zz_6008) * $signed(data_mid_2_63_real));
  assign _zz_1531 = _zz_6009;
  assign _zz_476 = _zz_6012[35 : 0];
  assign _zz_1532 = _zz_6013;
  assign _zz_477 = _zz_6016[35 : 0];
  assign _zz_479 = 1'b1;
  assign _zz_1533 = _zz_6017;
  assign _zz_1534 = _zz_6025;
  assign _zz_480 = 1'b1;
  assign _zz_1535 = _zz_6033;
  assign _zz_1536 = _zz_6041;
  assign _zz_483 = ($signed(_zz_6049) * $signed(data_mid_3_8_real));
  assign _zz_1537 = _zz_6050;
  assign _zz_481 = _zz_6053[35 : 0];
  assign _zz_1538 = _zz_6054;
  assign _zz_482 = _zz_6057[35 : 0];
  assign _zz_484 = 1'b1;
  assign _zz_1539 = _zz_6058;
  assign _zz_1540 = _zz_6066;
  assign _zz_485 = 1'b1;
  assign _zz_1541 = _zz_6074;
  assign _zz_1542 = _zz_6082;
  assign _zz_488 = ($signed(_zz_6090) * $signed(data_mid_3_9_real));
  assign _zz_1543 = _zz_6091;
  assign _zz_486 = _zz_6094[35 : 0];
  assign _zz_1544 = _zz_6095;
  assign _zz_487 = _zz_6098[35 : 0];
  assign _zz_489 = 1'b1;
  assign _zz_1545 = _zz_6099;
  assign _zz_1546 = _zz_6107;
  assign _zz_490 = 1'b1;
  assign _zz_1547 = _zz_6115;
  assign _zz_1548 = _zz_6123;
  assign _zz_493 = ($signed(_zz_6131) * $signed(data_mid_3_10_real));
  assign _zz_1549 = _zz_6132;
  assign _zz_491 = _zz_6135[35 : 0];
  assign _zz_1550 = _zz_6136;
  assign _zz_492 = _zz_6139[35 : 0];
  assign _zz_494 = 1'b1;
  assign _zz_1551 = _zz_6140;
  assign _zz_1552 = _zz_6148;
  assign _zz_495 = 1'b1;
  assign _zz_1553 = _zz_6156;
  assign _zz_1554 = _zz_6164;
  assign _zz_498 = ($signed(_zz_6172) * $signed(data_mid_3_11_real));
  assign _zz_1555 = _zz_6173;
  assign _zz_496 = _zz_6176[35 : 0];
  assign _zz_1556 = _zz_6177;
  assign _zz_497 = _zz_6180[35 : 0];
  assign _zz_499 = 1'b1;
  assign _zz_1557 = _zz_6181;
  assign _zz_1558 = _zz_6189;
  assign _zz_500 = 1'b1;
  assign _zz_1559 = _zz_6197;
  assign _zz_1560 = _zz_6205;
  assign _zz_503 = ($signed(_zz_6213) * $signed(data_mid_3_12_real));
  assign _zz_1561 = _zz_6214;
  assign _zz_501 = _zz_6217[35 : 0];
  assign _zz_1562 = _zz_6218;
  assign _zz_502 = _zz_6221[35 : 0];
  assign _zz_504 = 1'b1;
  assign _zz_1563 = _zz_6222;
  assign _zz_1564 = _zz_6230;
  assign _zz_505 = 1'b1;
  assign _zz_1565 = _zz_6238;
  assign _zz_1566 = _zz_6246;
  assign _zz_508 = ($signed(_zz_6254) * $signed(data_mid_3_13_real));
  assign _zz_1567 = _zz_6255;
  assign _zz_506 = _zz_6258[35 : 0];
  assign _zz_1568 = _zz_6259;
  assign _zz_507 = _zz_6262[35 : 0];
  assign _zz_509 = 1'b1;
  assign _zz_1569 = _zz_6263;
  assign _zz_1570 = _zz_6271;
  assign _zz_510 = 1'b1;
  assign _zz_1571 = _zz_6279;
  assign _zz_1572 = _zz_6287;
  assign _zz_513 = ($signed(_zz_6295) * $signed(data_mid_3_14_real));
  assign _zz_1573 = _zz_6296;
  assign _zz_511 = _zz_6299[35 : 0];
  assign _zz_1574 = _zz_6300;
  assign _zz_512 = _zz_6303[35 : 0];
  assign _zz_514 = 1'b1;
  assign _zz_1575 = _zz_6304;
  assign _zz_1576 = _zz_6312;
  assign _zz_515 = 1'b1;
  assign _zz_1577 = _zz_6320;
  assign _zz_1578 = _zz_6328;
  assign _zz_518 = ($signed(_zz_6336) * $signed(data_mid_3_15_real));
  assign _zz_1579 = _zz_6337;
  assign _zz_516 = _zz_6340[35 : 0];
  assign _zz_1580 = _zz_6341;
  assign _zz_517 = _zz_6344[35 : 0];
  assign _zz_519 = 1'b1;
  assign _zz_1581 = _zz_6345;
  assign _zz_1582 = _zz_6353;
  assign _zz_520 = 1'b1;
  assign _zz_1583 = _zz_6361;
  assign _zz_1584 = _zz_6369;
  assign _zz_523 = ($signed(_zz_6377) * $signed(data_mid_3_24_real));
  assign _zz_1585 = _zz_6378;
  assign _zz_521 = _zz_6381[35 : 0];
  assign _zz_1586 = _zz_6382;
  assign _zz_522 = _zz_6385[35 : 0];
  assign _zz_524 = 1'b1;
  assign _zz_1587 = _zz_6386;
  assign _zz_1588 = _zz_6394;
  assign _zz_525 = 1'b1;
  assign _zz_1589 = _zz_6402;
  assign _zz_1590 = _zz_6410;
  assign _zz_528 = ($signed(_zz_6418) * $signed(data_mid_3_25_real));
  assign _zz_1591 = _zz_6419;
  assign _zz_526 = _zz_6422[35 : 0];
  assign _zz_1592 = _zz_6423;
  assign _zz_527 = _zz_6426[35 : 0];
  assign _zz_529 = 1'b1;
  assign _zz_1593 = _zz_6427;
  assign _zz_1594 = _zz_6435;
  assign _zz_530 = 1'b1;
  assign _zz_1595 = _zz_6443;
  assign _zz_1596 = _zz_6451;
  assign _zz_533 = ($signed(_zz_6459) * $signed(data_mid_3_26_real));
  assign _zz_1597 = _zz_6460;
  assign _zz_531 = _zz_6463[35 : 0];
  assign _zz_1598 = _zz_6464;
  assign _zz_532 = _zz_6467[35 : 0];
  assign _zz_534 = 1'b1;
  assign _zz_1599 = _zz_6468;
  assign _zz_1600 = _zz_6476;
  assign _zz_535 = 1'b1;
  assign _zz_1601 = _zz_6484;
  assign _zz_1602 = _zz_6492;
  assign _zz_538 = ($signed(_zz_6500) * $signed(data_mid_3_27_real));
  assign _zz_1603 = _zz_6501;
  assign _zz_536 = _zz_6504[35 : 0];
  assign _zz_1604 = _zz_6505;
  assign _zz_537 = _zz_6508[35 : 0];
  assign _zz_539 = 1'b1;
  assign _zz_1605 = _zz_6509;
  assign _zz_1606 = _zz_6517;
  assign _zz_540 = 1'b1;
  assign _zz_1607 = _zz_6525;
  assign _zz_1608 = _zz_6533;
  assign _zz_543 = ($signed(_zz_6541) * $signed(data_mid_3_28_real));
  assign _zz_1609 = _zz_6542;
  assign _zz_541 = _zz_6545[35 : 0];
  assign _zz_1610 = _zz_6546;
  assign _zz_542 = _zz_6549[35 : 0];
  assign _zz_544 = 1'b1;
  assign _zz_1611 = _zz_6550;
  assign _zz_1612 = _zz_6558;
  assign _zz_545 = 1'b1;
  assign _zz_1613 = _zz_6566;
  assign _zz_1614 = _zz_6574;
  assign _zz_548 = ($signed(_zz_6582) * $signed(data_mid_3_29_real));
  assign _zz_1615 = _zz_6583;
  assign _zz_546 = _zz_6586[35 : 0];
  assign _zz_1616 = _zz_6587;
  assign _zz_547 = _zz_6590[35 : 0];
  assign _zz_549 = 1'b1;
  assign _zz_1617 = _zz_6591;
  assign _zz_1618 = _zz_6599;
  assign _zz_550 = 1'b1;
  assign _zz_1619 = _zz_6607;
  assign _zz_1620 = _zz_6615;
  assign _zz_553 = ($signed(_zz_6623) * $signed(data_mid_3_30_real));
  assign _zz_1621 = _zz_6624;
  assign _zz_551 = _zz_6627[35 : 0];
  assign _zz_1622 = _zz_6628;
  assign _zz_552 = _zz_6631[35 : 0];
  assign _zz_554 = 1'b1;
  assign _zz_1623 = _zz_6632;
  assign _zz_1624 = _zz_6640;
  assign _zz_555 = 1'b1;
  assign _zz_1625 = _zz_6648;
  assign _zz_1626 = _zz_6656;
  assign _zz_558 = ($signed(_zz_6664) * $signed(data_mid_3_31_real));
  assign _zz_1627 = _zz_6665;
  assign _zz_556 = _zz_6668[35 : 0];
  assign _zz_1628 = _zz_6669;
  assign _zz_557 = _zz_6672[35 : 0];
  assign _zz_559 = 1'b1;
  assign _zz_1629 = _zz_6673;
  assign _zz_1630 = _zz_6681;
  assign _zz_560 = 1'b1;
  assign _zz_1631 = _zz_6689;
  assign _zz_1632 = _zz_6697;
  assign _zz_563 = ($signed(_zz_6705) * $signed(data_mid_3_40_real));
  assign _zz_1633 = _zz_6706;
  assign _zz_561 = _zz_6709[35 : 0];
  assign _zz_1634 = _zz_6710;
  assign _zz_562 = _zz_6713[35 : 0];
  assign _zz_564 = 1'b1;
  assign _zz_1635 = _zz_6714;
  assign _zz_1636 = _zz_6722;
  assign _zz_565 = 1'b1;
  assign _zz_1637 = _zz_6730;
  assign _zz_1638 = _zz_6738;
  assign _zz_568 = ($signed(_zz_6746) * $signed(data_mid_3_41_real));
  assign _zz_1639 = _zz_6747;
  assign _zz_566 = _zz_6750[35 : 0];
  assign _zz_1640 = _zz_6751;
  assign _zz_567 = _zz_6754[35 : 0];
  assign _zz_569 = 1'b1;
  assign _zz_1641 = _zz_6755;
  assign _zz_1642 = _zz_6763;
  assign _zz_570 = 1'b1;
  assign _zz_1643 = _zz_6771;
  assign _zz_1644 = _zz_6779;
  assign _zz_573 = ($signed(_zz_6787) * $signed(data_mid_3_42_real));
  assign _zz_1645 = _zz_6788;
  assign _zz_571 = _zz_6791[35 : 0];
  assign _zz_1646 = _zz_6792;
  assign _zz_572 = _zz_6795[35 : 0];
  assign _zz_574 = 1'b1;
  assign _zz_1647 = _zz_6796;
  assign _zz_1648 = _zz_6804;
  assign _zz_575 = 1'b1;
  assign _zz_1649 = _zz_6812;
  assign _zz_1650 = _zz_6820;
  assign _zz_578 = ($signed(_zz_6828) * $signed(data_mid_3_43_real));
  assign _zz_1651 = _zz_6829;
  assign _zz_576 = _zz_6832[35 : 0];
  assign _zz_1652 = _zz_6833;
  assign _zz_577 = _zz_6836[35 : 0];
  assign _zz_579 = 1'b1;
  assign _zz_1653 = _zz_6837;
  assign _zz_1654 = _zz_6845;
  assign _zz_580 = 1'b1;
  assign _zz_1655 = _zz_6853;
  assign _zz_1656 = _zz_6861;
  assign _zz_583 = ($signed(_zz_6869) * $signed(data_mid_3_44_real));
  assign _zz_1657 = _zz_6870;
  assign _zz_581 = _zz_6873[35 : 0];
  assign _zz_1658 = _zz_6874;
  assign _zz_582 = _zz_6877[35 : 0];
  assign _zz_584 = 1'b1;
  assign _zz_1659 = _zz_6878;
  assign _zz_1660 = _zz_6886;
  assign _zz_585 = 1'b1;
  assign _zz_1661 = _zz_6894;
  assign _zz_1662 = _zz_6902;
  assign _zz_588 = ($signed(_zz_6910) * $signed(data_mid_3_45_real));
  assign _zz_1663 = _zz_6911;
  assign _zz_586 = _zz_6914[35 : 0];
  assign _zz_1664 = _zz_6915;
  assign _zz_587 = _zz_6918[35 : 0];
  assign _zz_589 = 1'b1;
  assign _zz_1665 = _zz_6919;
  assign _zz_1666 = _zz_6927;
  assign _zz_590 = 1'b1;
  assign _zz_1667 = _zz_6935;
  assign _zz_1668 = _zz_6943;
  assign _zz_593 = ($signed(_zz_6951) * $signed(data_mid_3_46_real));
  assign _zz_1669 = _zz_6952;
  assign _zz_591 = _zz_6955[35 : 0];
  assign _zz_1670 = _zz_6956;
  assign _zz_592 = _zz_6959[35 : 0];
  assign _zz_594 = 1'b1;
  assign _zz_1671 = _zz_6960;
  assign _zz_1672 = _zz_6968;
  assign _zz_595 = 1'b1;
  assign _zz_1673 = _zz_6976;
  assign _zz_1674 = _zz_6984;
  assign _zz_598 = ($signed(_zz_6992) * $signed(data_mid_3_47_real));
  assign _zz_1675 = _zz_6993;
  assign _zz_596 = _zz_6996[35 : 0];
  assign _zz_1676 = _zz_6997;
  assign _zz_597 = _zz_7000[35 : 0];
  assign _zz_599 = 1'b1;
  assign _zz_1677 = _zz_7001;
  assign _zz_1678 = _zz_7009;
  assign _zz_600 = 1'b1;
  assign _zz_1679 = _zz_7017;
  assign _zz_1680 = _zz_7025;
  assign _zz_603 = ($signed(_zz_7033) * $signed(data_mid_3_56_real));
  assign _zz_1681 = _zz_7034;
  assign _zz_601 = _zz_7037[35 : 0];
  assign _zz_1682 = _zz_7038;
  assign _zz_602 = _zz_7041[35 : 0];
  assign _zz_604 = 1'b1;
  assign _zz_1683 = _zz_7042;
  assign _zz_1684 = _zz_7050;
  assign _zz_605 = 1'b1;
  assign _zz_1685 = _zz_7058;
  assign _zz_1686 = _zz_7066;
  assign _zz_608 = ($signed(_zz_7074) * $signed(data_mid_3_57_real));
  assign _zz_1687 = _zz_7075;
  assign _zz_606 = _zz_7078[35 : 0];
  assign _zz_1688 = _zz_7079;
  assign _zz_607 = _zz_7082[35 : 0];
  assign _zz_609 = 1'b1;
  assign _zz_1689 = _zz_7083;
  assign _zz_1690 = _zz_7091;
  assign _zz_610 = 1'b1;
  assign _zz_1691 = _zz_7099;
  assign _zz_1692 = _zz_7107;
  assign _zz_613 = ($signed(_zz_7115) * $signed(data_mid_3_58_real));
  assign _zz_1693 = _zz_7116;
  assign _zz_611 = _zz_7119[35 : 0];
  assign _zz_1694 = _zz_7120;
  assign _zz_612 = _zz_7123[35 : 0];
  assign _zz_614 = 1'b1;
  assign _zz_1695 = _zz_7124;
  assign _zz_1696 = _zz_7132;
  assign _zz_615 = 1'b1;
  assign _zz_1697 = _zz_7140;
  assign _zz_1698 = _zz_7148;
  assign _zz_618 = ($signed(_zz_7156) * $signed(data_mid_3_59_real));
  assign _zz_1699 = _zz_7157;
  assign _zz_616 = _zz_7160[35 : 0];
  assign _zz_1700 = _zz_7161;
  assign _zz_617 = _zz_7164[35 : 0];
  assign _zz_619 = 1'b1;
  assign _zz_1701 = _zz_7165;
  assign _zz_1702 = _zz_7173;
  assign _zz_620 = 1'b1;
  assign _zz_1703 = _zz_7181;
  assign _zz_1704 = _zz_7189;
  assign _zz_623 = ($signed(_zz_7197) * $signed(data_mid_3_60_real));
  assign _zz_1705 = _zz_7198;
  assign _zz_621 = _zz_7201[35 : 0];
  assign _zz_1706 = _zz_7202;
  assign _zz_622 = _zz_7205[35 : 0];
  assign _zz_624 = 1'b1;
  assign _zz_1707 = _zz_7206;
  assign _zz_1708 = _zz_7214;
  assign _zz_625 = 1'b1;
  assign _zz_1709 = _zz_7222;
  assign _zz_1710 = _zz_7230;
  assign _zz_628 = ($signed(_zz_7238) * $signed(data_mid_3_61_real));
  assign _zz_1711 = _zz_7239;
  assign _zz_626 = _zz_7242[35 : 0];
  assign _zz_1712 = _zz_7243;
  assign _zz_627 = _zz_7246[35 : 0];
  assign _zz_629 = 1'b1;
  assign _zz_1713 = _zz_7247;
  assign _zz_1714 = _zz_7255;
  assign _zz_630 = 1'b1;
  assign _zz_1715 = _zz_7263;
  assign _zz_1716 = _zz_7271;
  assign _zz_633 = ($signed(_zz_7279) * $signed(data_mid_3_62_real));
  assign _zz_1717 = _zz_7280;
  assign _zz_631 = _zz_7283[35 : 0];
  assign _zz_1718 = _zz_7284;
  assign _zz_632 = _zz_7287[35 : 0];
  assign _zz_634 = 1'b1;
  assign _zz_1719 = _zz_7288;
  assign _zz_1720 = _zz_7296;
  assign _zz_635 = 1'b1;
  assign _zz_1721 = _zz_7304;
  assign _zz_1722 = _zz_7312;
  assign _zz_638 = ($signed(_zz_7320) * $signed(data_mid_3_63_real));
  assign _zz_1723 = _zz_7321;
  assign _zz_636 = _zz_7324[35 : 0];
  assign _zz_1724 = _zz_7325;
  assign _zz_637 = _zz_7328[35 : 0];
  assign _zz_639 = 1'b1;
  assign _zz_1725 = _zz_7329;
  assign _zz_1726 = _zz_7337;
  assign _zz_640 = 1'b1;
  assign _zz_1727 = _zz_7345;
  assign _zz_1728 = _zz_7353;
  assign _zz_643 = ($signed(_zz_7361) * $signed(data_mid_4_16_real));
  assign _zz_1729 = _zz_7362;
  assign _zz_641 = _zz_7365[35 : 0];
  assign _zz_1730 = _zz_7366;
  assign _zz_642 = _zz_7369[35 : 0];
  assign _zz_644 = 1'b1;
  assign _zz_1731 = _zz_7370;
  assign _zz_1732 = _zz_7378;
  assign _zz_645 = 1'b1;
  assign _zz_1733 = _zz_7386;
  assign _zz_1734 = _zz_7394;
  assign _zz_648 = ($signed(_zz_7402) * $signed(data_mid_4_17_real));
  assign _zz_1735 = _zz_7403;
  assign _zz_646 = _zz_7406[35 : 0];
  assign _zz_1736 = _zz_7407;
  assign _zz_647 = _zz_7410[35 : 0];
  assign _zz_649 = 1'b1;
  assign _zz_1737 = _zz_7411;
  assign _zz_1738 = _zz_7419;
  assign _zz_650 = 1'b1;
  assign _zz_1739 = _zz_7427;
  assign _zz_1740 = _zz_7435;
  assign _zz_653 = ($signed(_zz_7443) * $signed(data_mid_4_18_real));
  assign _zz_1741 = _zz_7444;
  assign _zz_651 = _zz_7447[35 : 0];
  assign _zz_1742 = _zz_7448;
  assign _zz_652 = _zz_7451[35 : 0];
  assign _zz_654 = 1'b1;
  assign _zz_1743 = _zz_7452;
  assign _zz_1744 = _zz_7460;
  assign _zz_655 = 1'b1;
  assign _zz_1745 = _zz_7468;
  assign _zz_1746 = _zz_7476;
  assign _zz_658 = ($signed(_zz_7484) * $signed(data_mid_4_19_real));
  assign _zz_1747 = _zz_7485;
  assign _zz_656 = _zz_7488[35 : 0];
  assign _zz_1748 = _zz_7489;
  assign _zz_657 = _zz_7492[35 : 0];
  assign _zz_659 = 1'b1;
  assign _zz_1749 = _zz_7493;
  assign _zz_1750 = _zz_7501;
  assign _zz_660 = 1'b1;
  assign _zz_1751 = _zz_7509;
  assign _zz_1752 = _zz_7517;
  assign _zz_663 = ($signed(_zz_7525) * $signed(data_mid_4_20_real));
  assign _zz_1753 = _zz_7526;
  assign _zz_661 = _zz_7529[35 : 0];
  assign _zz_1754 = _zz_7530;
  assign _zz_662 = _zz_7533[35 : 0];
  assign _zz_664 = 1'b1;
  assign _zz_1755 = _zz_7534;
  assign _zz_1756 = _zz_7542;
  assign _zz_665 = 1'b1;
  assign _zz_1757 = _zz_7550;
  assign _zz_1758 = _zz_7558;
  assign _zz_668 = ($signed(_zz_7566) * $signed(data_mid_4_21_real));
  assign _zz_1759 = _zz_7567;
  assign _zz_666 = _zz_7570[35 : 0];
  assign _zz_1760 = _zz_7571;
  assign _zz_667 = _zz_7574[35 : 0];
  assign _zz_669 = 1'b1;
  assign _zz_1761 = _zz_7575;
  assign _zz_1762 = _zz_7583;
  assign _zz_670 = 1'b1;
  assign _zz_1763 = _zz_7591;
  assign _zz_1764 = _zz_7599;
  assign _zz_673 = ($signed(_zz_7607) * $signed(data_mid_4_22_real));
  assign _zz_1765 = _zz_7608;
  assign _zz_671 = _zz_7611[35 : 0];
  assign _zz_1766 = _zz_7612;
  assign _zz_672 = _zz_7615[35 : 0];
  assign _zz_674 = 1'b1;
  assign _zz_1767 = _zz_7616;
  assign _zz_1768 = _zz_7624;
  assign _zz_675 = 1'b1;
  assign _zz_1769 = _zz_7632;
  assign _zz_1770 = _zz_7640;
  assign _zz_678 = ($signed(_zz_7648) * $signed(data_mid_4_23_real));
  assign _zz_1771 = _zz_7649;
  assign _zz_676 = _zz_7652[35 : 0];
  assign _zz_1772 = _zz_7653;
  assign _zz_677 = _zz_7656[35 : 0];
  assign _zz_679 = 1'b1;
  assign _zz_1773 = _zz_7657;
  assign _zz_1774 = _zz_7665;
  assign _zz_680 = 1'b1;
  assign _zz_1775 = _zz_7673;
  assign _zz_1776 = _zz_7681;
  assign _zz_683 = ($signed(_zz_7689) * $signed(data_mid_4_24_real));
  assign _zz_1777 = _zz_7690;
  assign _zz_681 = _zz_7693[35 : 0];
  assign _zz_1778 = _zz_7694;
  assign _zz_682 = _zz_7697[35 : 0];
  assign _zz_684 = 1'b1;
  assign _zz_1779 = _zz_7698;
  assign _zz_1780 = _zz_7706;
  assign _zz_685 = 1'b1;
  assign _zz_1781 = _zz_7714;
  assign _zz_1782 = _zz_7722;
  assign _zz_688 = ($signed(_zz_7730) * $signed(data_mid_4_25_real));
  assign _zz_1783 = _zz_7731;
  assign _zz_686 = _zz_7734[35 : 0];
  assign _zz_1784 = _zz_7735;
  assign _zz_687 = _zz_7738[35 : 0];
  assign _zz_689 = 1'b1;
  assign _zz_1785 = _zz_7739;
  assign _zz_1786 = _zz_7747;
  assign _zz_690 = 1'b1;
  assign _zz_1787 = _zz_7755;
  assign _zz_1788 = _zz_7763;
  assign _zz_693 = ($signed(_zz_7771) * $signed(data_mid_4_26_real));
  assign _zz_1789 = _zz_7772;
  assign _zz_691 = _zz_7775[35 : 0];
  assign _zz_1790 = _zz_7776;
  assign _zz_692 = _zz_7779[35 : 0];
  assign _zz_694 = 1'b1;
  assign _zz_1791 = _zz_7780;
  assign _zz_1792 = _zz_7788;
  assign _zz_695 = 1'b1;
  assign _zz_1793 = _zz_7796;
  assign _zz_1794 = _zz_7804;
  assign _zz_698 = ($signed(_zz_7812) * $signed(data_mid_4_27_real));
  assign _zz_1795 = _zz_7813;
  assign _zz_696 = _zz_7816[35 : 0];
  assign _zz_1796 = _zz_7817;
  assign _zz_697 = _zz_7820[35 : 0];
  assign _zz_699 = 1'b1;
  assign _zz_1797 = _zz_7821;
  assign _zz_1798 = _zz_7829;
  assign _zz_700 = 1'b1;
  assign _zz_1799 = _zz_7837;
  assign _zz_1800 = _zz_7845;
  assign _zz_703 = ($signed(_zz_7853) * $signed(data_mid_4_28_real));
  assign _zz_1801 = _zz_7854;
  assign _zz_701 = _zz_7857[35 : 0];
  assign _zz_1802 = _zz_7858;
  assign _zz_702 = _zz_7861[35 : 0];
  assign _zz_704 = 1'b1;
  assign _zz_1803 = _zz_7862;
  assign _zz_1804 = _zz_7870;
  assign _zz_705 = 1'b1;
  assign _zz_1805 = _zz_7878;
  assign _zz_1806 = _zz_7886;
  assign _zz_708 = ($signed(_zz_7894) * $signed(data_mid_4_29_real));
  assign _zz_1807 = _zz_7895;
  assign _zz_706 = _zz_7898[35 : 0];
  assign _zz_1808 = _zz_7899;
  assign _zz_707 = _zz_7902[35 : 0];
  assign _zz_709 = 1'b1;
  assign _zz_1809 = _zz_7903;
  assign _zz_1810 = _zz_7911;
  assign _zz_710 = 1'b1;
  assign _zz_1811 = _zz_7919;
  assign _zz_1812 = _zz_7927;
  assign _zz_713 = ($signed(_zz_7935) * $signed(data_mid_4_30_real));
  assign _zz_1813 = _zz_7936;
  assign _zz_711 = _zz_7939[35 : 0];
  assign _zz_1814 = _zz_7940;
  assign _zz_712 = _zz_7943[35 : 0];
  assign _zz_714 = 1'b1;
  assign _zz_1815 = _zz_7944;
  assign _zz_1816 = _zz_7952;
  assign _zz_715 = 1'b1;
  assign _zz_1817 = _zz_7960;
  assign _zz_1818 = _zz_7968;
  assign _zz_718 = ($signed(_zz_7976) * $signed(data_mid_4_31_real));
  assign _zz_1819 = _zz_7977;
  assign _zz_716 = _zz_7980[35 : 0];
  assign _zz_1820 = _zz_7981;
  assign _zz_717 = _zz_7984[35 : 0];
  assign _zz_719 = 1'b1;
  assign _zz_1821 = _zz_7985;
  assign _zz_1822 = _zz_7993;
  assign _zz_720 = 1'b1;
  assign _zz_1823 = _zz_8001;
  assign _zz_1824 = _zz_8009;
  assign _zz_723 = ($signed(_zz_8017) * $signed(data_mid_4_48_real));
  assign _zz_1825 = _zz_8018;
  assign _zz_721 = _zz_8021[35 : 0];
  assign _zz_1826 = _zz_8022;
  assign _zz_722 = _zz_8025[35 : 0];
  assign _zz_724 = 1'b1;
  assign _zz_1827 = _zz_8026;
  assign _zz_1828 = _zz_8034;
  assign _zz_725 = 1'b1;
  assign _zz_1829 = _zz_8042;
  assign _zz_1830 = _zz_8050;
  assign _zz_728 = ($signed(_zz_8058) * $signed(data_mid_4_49_real));
  assign _zz_1831 = _zz_8059;
  assign _zz_726 = _zz_8062[35 : 0];
  assign _zz_1832 = _zz_8063;
  assign _zz_727 = _zz_8066[35 : 0];
  assign _zz_729 = 1'b1;
  assign _zz_1833 = _zz_8067;
  assign _zz_1834 = _zz_8075;
  assign _zz_730 = 1'b1;
  assign _zz_1835 = _zz_8083;
  assign _zz_1836 = _zz_8091;
  assign _zz_733 = ($signed(_zz_8099) * $signed(data_mid_4_50_real));
  assign _zz_1837 = _zz_8100;
  assign _zz_731 = _zz_8103[35 : 0];
  assign _zz_1838 = _zz_8104;
  assign _zz_732 = _zz_8107[35 : 0];
  assign _zz_734 = 1'b1;
  assign _zz_1839 = _zz_8108;
  assign _zz_1840 = _zz_8116;
  assign _zz_735 = 1'b1;
  assign _zz_1841 = _zz_8124;
  assign _zz_1842 = _zz_8132;
  assign _zz_738 = ($signed(_zz_8140) * $signed(data_mid_4_51_real));
  assign _zz_1843 = _zz_8141;
  assign _zz_736 = _zz_8144[35 : 0];
  assign _zz_1844 = _zz_8145;
  assign _zz_737 = _zz_8148[35 : 0];
  assign _zz_739 = 1'b1;
  assign _zz_1845 = _zz_8149;
  assign _zz_1846 = _zz_8157;
  assign _zz_740 = 1'b1;
  assign _zz_1847 = _zz_8165;
  assign _zz_1848 = _zz_8173;
  assign _zz_743 = ($signed(_zz_8181) * $signed(data_mid_4_52_real));
  assign _zz_1849 = _zz_8182;
  assign _zz_741 = _zz_8185[35 : 0];
  assign _zz_1850 = _zz_8186;
  assign _zz_742 = _zz_8189[35 : 0];
  assign _zz_744 = 1'b1;
  assign _zz_1851 = _zz_8190;
  assign _zz_1852 = _zz_8198;
  assign _zz_745 = 1'b1;
  assign _zz_1853 = _zz_8206;
  assign _zz_1854 = _zz_8214;
  assign _zz_748 = ($signed(_zz_8222) * $signed(data_mid_4_53_real));
  assign _zz_1855 = _zz_8223;
  assign _zz_746 = _zz_8226[35 : 0];
  assign _zz_1856 = _zz_8227;
  assign _zz_747 = _zz_8230[35 : 0];
  assign _zz_749 = 1'b1;
  assign _zz_1857 = _zz_8231;
  assign _zz_1858 = _zz_8239;
  assign _zz_750 = 1'b1;
  assign _zz_1859 = _zz_8247;
  assign _zz_1860 = _zz_8255;
  assign _zz_753 = ($signed(_zz_8263) * $signed(data_mid_4_54_real));
  assign _zz_1861 = _zz_8264;
  assign _zz_751 = _zz_8267[35 : 0];
  assign _zz_1862 = _zz_8268;
  assign _zz_752 = _zz_8271[35 : 0];
  assign _zz_754 = 1'b1;
  assign _zz_1863 = _zz_8272;
  assign _zz_1864 = _zz_8280;
  assign _zz_755 = 1'b1;
  assign _zz_1865 = _zz_8288;
  assign _zz_1866 = _zz_8296;
  assign _zz_758 = ($signed(_zz_8304) * $signed(data_mid_4_55_real));
  assign _zz_1867 = _zz_8305;
  assign _zz_756 = _zz_8308[35 : 0];
  assign _zz_1868 = _zz_8309;
  assign _zz_757 = _zz_8312[35 : 0];
  assign _zz_759 = 1'b1;
  assign _zz_1869 = _zz_8313;
  assign _zz_1870 = _zz_8321;
  assign _zz_760 = 1'b1;
  assign _zz_1871 = _zz_8329;
  assign _zz_1872 = _zz_8337;
  assign _zz_763 = ($signed(_zz_8345) * $signed(data_mid_4_56_real));
  assign _zz_1873 = _zz_8346;
  assign _zz_761 = _zz_8349[35 : 0];
  assign _zz_1874 = _zz_8350;
  assign _zz_762 = _zz_8353[35 : 0];
  assign _zz_764 = 1'b1;
  assign _zz_1875 = _zz_8354;
  assign _zz_1876 = _zz_8362;
  assign _zz_765 = 1'b1;
  assign _zz_1877 = _zz_8370;
  assign _zz_1878 = _zz_8378;
  assign _zz_768 = ($signed(_zz_8386) * $signed(data_mid_4_57_real));
  assign _zz_1879 = _zz_8387;
  assign _zz_766 = _zz_8390[35 : 0];
  assign _zz_1880 = _zz_8391;
  assign _zz_767 = _zz_8394[35 : 0];
  assign _zz_769 = 1'b1;
  assign _zz_1881 = _zz_8395;
  assign _zz_1882 = _zz_8403;
  assign _zz_770 = 1'b1;
  assign _zz_1883 = _zz_8411;
  assign _zz_1884 = _zz_8419;
  assign _zz_773 = ($signed(_zz_8427) * $signed(data_mid_4_58_real));
  assign _zz_1885 = _zz_8428;
  assign _zz_771 = _zz_8431[35 : 0];
  assign _zz_1886 = _zz_8432;
  assign _zz_772 = _zz_8435[35 : 0];
  assign _zz_774 = 1'b1;
  assign _zz_1887 = _zz_8436;
  assign _zz_1888 = _zz_8444;
  assign _zz_775 = 1'b1;
  assign _zz_1889 = _zz_8452;
  assign _zz_1890 = _zz_8460;
  assign _zz_778 = ($signed(_zz_8468) * $signed(data_mid_4_59_real));
  assign _zz_1891 = _zz_8469;
  assign _zz_776 = _zz_8472[35 : 0];
  assign _zz_1892 = _zz_8473;
  assign _zz_777 = _zz_8476[35 : 0];
  assign _zz_779 = 1'b1;
  assign _zz_1893 = _zz_8477;
  assign _zz_1894 = _zz_8485;
  assign _zz_780 = 1'b1;
  assign _zz_1895 = _zz_8493;
  assign _zz_1896 = _zz_8501;
  assign _zz_783 = ($signed(_zz_8509) * $signed(data_mid_4_60_real));
  assign _zz_1897 = _zz_8510;
  assign _zz_781 = _zz_8513[35 : 0];
  assign _zz_1898 = _zz_8514;
  assign _zz_782 = _zz_8517[35 : 0];
  assign _zz_784 = 1'b1;
  assign _zz_1899 = _zz_8518;
  assign _zz_1900 = _zz_8526;
  assign _zz_785 = 1'b1;
  assign _zz_1901 = _zz_8534;
  assign _zz_1902 = _zz_8542;
  assign _zz_788 = ($signed(_zz_8550) * $signed(data_mid_4_61_real));
  assign _zz_1903 = _zz_8551;
  assign _zz_786 = _zz_8554[35 : 0];
  assign _zz_1904 = _zz_8555;
  assign _zz_787 = _zz_8558[35 : 0];
  assign _zz_789 = 1'b1;
  assign _zz_1905 = _zz_8559;
  assign _zz_1906 = _zz_8567;
  assign _zz_790 = 1'b1;
  assign _zz_1907 = _zz_8575;
  assign _zz_1908 = _zz_8583;
  assign _zz_793 = ($signed(_zz_8591) * $signed(data_mid_4_62_real));
  assign _zz_1909 = _zz_8592;
  assign _zz_791 = _zz_8595[35 : 0];
  assign _zz_1910 = _zz_8596;
  assign _zz_792 = _zz_8599[35 : 0];
  assign _zz_794 = 1'b1;
  assign _zz_1911 = _zz_8600;
  assign _zz_1912 = _zz_8608;
  assign _zz_795 = 1'b1;
  assign _zz_1913 = _zz_8616;
  assign _zz_1914 = _zz_8624;
  assign _zz_798 = ($signed(_zz_8632) * $signed(data_mid_4_63_real));
  assign _zz_1915 = _zz_8633;
  assign _zz_796 = _zz_8636[35 : 0];
  assign _zz_1916 = _zz_8637;
  assign _zz_797 = _zz_8640[35 : 0];
  assign _zz_799 = 1'b1;
  assign _zz_1917 = _zz_8641;
  assign _zz_1918 = _zz_8649;
  assign _zz_800 = 1'b1;
  assign _zz_1919 = _zz_8657;
  assign _zz_1920 = _zz_8665;
  assign _zz_803 = ($signed(_zz_8673) * $signed(data_mid_5_32_real));
  assign _zz_1921 = _zz_8674;
  assign _zz_801 = _zz_8677[35 : 0];
  assign _zz_1922 = _zz_8678;
  assign _zz_802 = _zz_8681[35 : 0];
  assign _zz_804 = 1'b1;
  assign _zz_1923 = _zz_8682;
  assign _zz_1924 = _zz_8690;
  assign _zz_805 = 1'b1;
  assign _zz_1925 = _zz_8698;
  assign _zz_1926 = _zz_8706;
  assign _zz_808 = ($signed(_zz_8714) * $signed(data_mid_5_33_real));
  assign _zz_1927 = _zz_8715;
  assign _zz_806 = _zz_8718[35 : 0];
  assign _zz_1928 = _zz_8719;
  assign _zz_807 = _zz_8722[35 : 0];
  assign _zz_809 = 1'b1;
  assign _zz_1929 = _zz_8723;
  assign _zz_1930 = _zz_8731;
  assign _zz_810 = 1'b1;
  assign _zz_1931 = _zz_8739;
  assign _zz_1932 = _zz_8747;
  assign _zz_813 = ($signed(_zz_8755) * $signed(data_mid_5_34_real));
  assign _zz_1933 = _zz_8756;
  assign _zz_811 = _zz_8759[35 : 0];
  assign _zz_1934 = _zz_8760;
  assign _zz_812 = _zz_8763[35 : 0];
  assign _zz_814 = 1'b1;
  assign _zz_1935 = _zz_8764;
  assign _zz_1936 = _zz_8772;
  assign _zz_815 = 1'b1;
  assign _zz_1937 = _zz_8780;
  assign _zz_1938 = _zz_8788;
  assign _zz_818 = ($signed(_zz_8796) * $signed(data_mid_5_35_real));
  assign _zz_1939 = _zz_8797;
  assign _zz_816 = _zz_8800[35 : 0];
  assign _zz_1940 = _zz_8801;
  assign _zz_817 = _zz_8804[35 : 0];
  assign _zz_819 = 1'b1;
  assign _zz_1941 = _zz_8805;
  assign _zz_1942 = _zz_8813;
  assign _zz_820 = 1'b1;
  assign _zz_1943 = _zz_8821;
  assign _zz_1944 = _zz_8829;
  assign _zz_823 = ($signed(_zz_8837) * $signed(data_mid_5_36_real));
  assign _zz_1945 = _zz_8838;
  assign _zz_821 = _zz_8841[35 : 0];
  assign _zz_1946 = _zz_8842;
  assign _zz_822 = _zz_8845[35 : 0];
  assign _zz_824 = 1'b1;
  assign _zz_1947 = _zz_8846;
  assign _zz_1948 = _zz_8854;
  assign _zz_825 = 1'b1;
  assign _zz_1949 = _zz_8862;
  assign _zz_1950 = _zz_8870;
  assign _zz_828 = ($signed(_zz_8878) * $signed(data_mid_5_37_real));
  assign _zz_1951 = _zz_8879;
  assign _zz_826 = _zz_8882[35 : 0];
  assign _zz_1952 = _zz_8883;
  assign _zz_827 = _zz_8886[35 : 0];
  assign _zz_829 = 1'b1;
  assign _zz_1953 = _zz_8887;
  assign _zz_1954 = _zz_8895;
  assign _zz_830 = 1'b1;
  assign _zz_1955 = _zz_8903;
  assign _zz_1956 = _zz_8911;
  assign _zz_833 = ($signed(_zz_8919) * $signed(data_mid_5_38_real));
  assign _zz_1957 = _zz_8920;
  assign _zz_831 = _zz_8923[35 : 0];
  assign _zz_1958 = _zz_8924;
  assign _zz_832 = _zz_8927[35 : 0];
  assign _zz_834 = 1'b1;
  assign _zz_1959 = _zz_8928;
  assign _zz_1960 = _zz_8936;
  assign _zz_835 = 1'b1;
  assign _zz_1961 = _zz_8944;
  assign _zz_1962 = _zz_8952;
  assign _zz_838 = ($signed(_zz_8960) * $signed(data_mid_5_39_real));
  assign _zz_1963 = _zz_8961;
  assign _zz_836 = _zz_8964[35 : 0];
  assign _zz_1964 = _zz_8965;
  assign _zz_837 = _zz_8968[35 : 0];
  assign _zz_839 = 1'b1;
  assign _zz_1965 = _zz_8969;
  assign _zz_1966 = _zz_8977;
  assign _zz_840 = 1'b1;
  assign _zz_1967 = _zz_8985;
  assign _zz_1968 = _zz_8993;
  assign _zz_843 = ($signed(_zz_9001) * $signed(data_mid_5_40_real));
  assign _zz_1969 = _zz_9002;
  assign _zz_841 = _zz_9005[35 : 0];
  assign _zz_1970 = _zz_9006;
  assign _zz_842 = _zz_9009[35 : 0];
  assign _zz_844 = 1'b1;
  assign _zz_1971 = _zz_9010;
  assign _zz_1972 = _zz_9018;
  assign _zz_845 = 1'b1;
  assign _zz_1973 = _zz_9026;
  assign _zz_1974 = _zz_9034;
  assign _zz_848 = ($signed(_zz_9042) * $signed(data_mid_5_41_real));
  assign _zz_1975 = _zz_9043;
  assign _zz_846 = _zz_9046[35 : 0];
  assign _zz_1976 = _zz_9047;
  assign _zz_847 = _zz_9050[35 : 0];
  assign _zz_849 = 1'b1;
  assign _zz_1977 = _zz_9051;
  assign _zz_1978 = _zz_9059;
  assign _zz_850 = 1'b1;
  assign _zz_1979 = _zz_9067;
  assign _zz_1980 = _zz_9075;
  assign _zz_853 = ($signed(_zz_9083) * $signed(data_mid_5_42_real));
  assign _zz_1981 = _zz_9084;
  assign _zz_851 = _zz_9087[35 : 0];
  assign _zz_1982 = _zz_9088;
  assign _zz_852 = _zz_9091[35 : 0];
  assign _zz_854 = 1'b1;
  assign _zz_1983 = _zz_9092;
  assign _zz_1984 = _zz_9100;
  assign _zz_855 = 1'b1;
  assign _zz_1985 = _zz_9108;
  assign _zz_1986 = _zz_9116;
  assign _zz_858 = ($signed(_zz_9124) * $signed(data_mid_5_43_real));
  assign _zz_1987 = _zz_9125;
  assign _zz_856 = _zz_9128[35 : 0];
  assign _zz_1988 = _zz_9129;
  assign _zz_857 = _zz_9132[35 : 0];
  assign _zz_859 = 1'b1;
  assign _zz_1989 = _zz_9133;
  assign _zz_1990 = _zz_9141;
  assign _zz_860 = 1'b1;
  assign _zz_1991 = _zz_9149;
  assign _zz_1992 = _zz_9157;
  assign _zz_863 = ($signed(_zz_9165) * $signed(data_mid_5_44_real));
  assign _zz_1993 = _zz_9166;
  assign _zz_861 = _zz_9169[35 : 0];
  assign _zz_1994 = _zz_9170;
  assign _zz_862 = _zz_9173[35 : 0];
  assign _zz_864 = 1'b1;
  assign _zz_1995 = _zz_9174;
  assign _zz_1996 = _zz_9182;
  assign _zz_865 = 1'b1;
  assign _zz_1997 = _zz_9190;
  assign _zz_1998 = _zz_9198;
  assign _zz_868 = ($signed(_zz_9206) * $signed(data_mid_5_45_real));
  assign _zz_1999 = _zz_9207;
  assign _zz_866 = _zz_9210[35 : 0];
  assign _zz_2000 = _zz_9211;
  assign _zz_867 = _zz_9214[35 : 0];
  assign _zz_869 = 1'b1;
  assign _zz_2001 = _zz_9215;
  assign _zz_2002 = _zz_9223;
  assign _zz_870 = 1'b1;
  assign _zz_2003 = _zz_9231;
  assign _zz_2004 = _zz_9239;
  assign _zz_873 = ($signed(_zz_9247) * $signed(data_mid_5_46_real));
  assign _zz_2005 = _zz_9248;
  assign _zz_871 = _zz_9251[35 : 0];
  assign _zz_2006 = _zz_9252;
  assign _zz_872 = _zz_9255[35 : 0];
  assign _zz_874 = 1'b1;
  assign _zz_2007 = _zz_9256;
  assign _zz_2008 = _zz_9264;
  assign _zz_875 = 1'b1;
  assign _zz_2009 = _zz_9272;
  assign _zz_2010 = _zz_9280;
  assign _zz_878 = ($signed(_zz_9288) * $signed(data_mid_5_47_real));
  assign _zz_2011 = _zz_9289;
  assign _zz_876 = _zz_9292[35 : 0];
  assign _zz_2012 = _zz_9293;
  assign _zz_877 = _zz_9296[35 : 0];
  assign _zz_879 = 1'b1;
  assign _zz_2013 = _zz_9297;
  assign _zz_2014 = _zz_9305;
  assign _zz_880 = 1'b1;
  assign _zz_2015 = _zz_9313;
  assign _zz_2016 = _zz_9321;
  assign _zz_883 = ($signed(_zz_9329) * $signed(data_mid_5_48_real));
  assign _zz_2017 = _zz_9330;
  assign _zz_881 = _zz_9333[35 : 0];
  assign _zz_2018 = _zz_9334;
  assign _zz_882 = _zz_9337[35 : 0];
  assign _zz_884 = 1'b1;
  assign _zz_2019 = _zz_9338;
  assign _zz_2020 = _zz_9346;
  assign _zz_885 = 1'b1;
  assign _zz_2021 = _zz_9354;
  assign _zz_2022 = _zz_9362;
  assign _zz_888 = ($signed(_zz_9370) * $signed(data_mid_5_49_real));
  assign _zz_2023 = _zz_9371;
  assign _zz_886 = _zz_9374[35 : 0];
  assign _zz_2024 = _zz_9375;
  assign _zz_887 = _zz_9378[35 : 0];
  assign _zz_889 = 1'b1;
  assign _zz_2025 = _zz_9379;
  assign _zz_2026 = _zz_9387;
  assign _zz_890 = 1'b1;
  assign _zz_2027 = _zz_9395;
  assign _zz_2028 = _zz_9403;
  assign _zz_893 = ($signed(_zz_9411) * $signed(data_mid_5_50_real));
  assign _zz_2029 = _zz_9412;
  assign _zz_891 = _zz_9415[35 : 0];
  assign _zz_2030 = _zz_9416;
  assign _zz_892 = _zz_9419[35 : 0];
  assign _zz_894 = 1'b1;
  assign _zz_2031 = _zz_9420;
  assign _zz_2032 = _zz_9428;
  assign _zz_895 = 1'b1;
  assign _zz_2033 = _zz_9436;
  assign _zz_2034 = _zz_9444;
  assign _zz_898 = ($signed(_zz_9452) * $signed(data_mid_5_51_real));
  assign _zz_2035 = _zz_9453;
  assign _zz_896 = _zz_9456[35 : 0];
  assign _zz_2036 = _zz_9457;
  assign _zz_897 = _zz_9460[35 : 0];
  assign _zz_899 = 1'b1;
  assign _zz_2037 = _zz_9461;
  assign _zz_2038 = _zz_9469;
  assign _zz_900 = 1'b1;
  assign _zz_2039 = _zz_9477;
  assign _zz_2040 = _zz_9485;
  assign _zz_903 = ($signed(_zz_9493) * $signed(data_mid_5_52_real));
  assign _zz_2041 = _zz_9494;
  assign _zz_901 = _zz_9497[35 : 0];
  assign _zz_2042 = _zz_9498;
  assign _zz_902 = _zz_9501[35 : 0];
  assign _zz_904 = 1'b1;
  assign _zz_2043 = _zz_9502;
  assign _zz_2044 = _zz_9510;
  assign _zz_905 = 1'b1;
  assign _zz_2045 = _zz_9518;
  assign _zz_2046 = _zz_9526;
  assign _zz_908 = ($signed(_zz_9534) * $signed(data_mid_5_53_real));
  assign _zz_2047 = _zz_9535;
  assign _zz_906 = _zz_9538[35 : 0];
  assign _zz_2048 = _zz_9539;
  assign _zz_907 = _zz_9542[35 : 0];
  assign _zz_909 = 1'b1;
  assign _zz_2049 = _zz_9543;
  assign _zz_2050 = _zz_9551;
  assign _zz_910 = 1'b1;
  assign _zz_2051 = _zz_9559;
  assign _zz_2052 = _zz_9567;
  assign _zz_913 = ($signed(_zz_9575) * $signed(data_mid_5_54_real));
  assign _zz_2053 = _zz_9576;
  assign _zz_911 = _zz_9579[35 : 0];
  assign _zz_2054 = _zz_9580;
  assign _zz_912 = _zz_9583[35 : 0];
  assign _zz_914 = 1'b1;
  assign _zz_2055 = _zz_9584;
  assign _zz_2056 = _zz_9592;
  assign _zz_915 = 1'b1;
  assign _zz_2057 = _zz_9600;
  assign _zz_2058 = _zz_9608;
  assign _zz_918 = ($signed(_zz_9616) * $signed(data_mid_5_55_real));
  assign _zz_2059 = _zz_9617;
  assign _zz_916 = _zz_9620[35 : 0];
  assign _zz_2060 = _zz_9621;
  assign _zz_917 = _zz_9624[35 : 0];
  assign _zz_919 = 1'b1;
  assign _zz_2061 = _zz_9625;
  assign _zz_2062 = _zz_9633;
  assign _zz_920 = 1'b1;
  assign _zz_2063 = _zz_9641;
  assign _zz_2064 = _zz_9649;
  assign _zz_923 = ($signed(_zz_9657) * $signed(data_mid_5_56_real));
  assign _zz_2065 = _zz_9658;
  assign _zz_921 = _zz_9661[35 : 0];
  assign _zz_2066 = _zz_9662;
  assign _zz_922 = _zz_9665[35 : 0];
  assign _zz_924 = 1'b1;
  assign _zz_2067 = _zz_9666;
  assign _zz_2068 = _zz_9674;
  assign _zz_925 = 1'b1;
  assign _zz_2069 = _zz_9682;
  assign _zz_2070 = _zz_9690;
  assign _zz_928 = ($signed(_zz_9698) * $signed(data_mid_5_57_real));
  assign _zz_2071 = _zz_9699;
  assign _zz_926 = _zz_9702[35 : 0];
  assign _zz_2072 = _zz_9703;
  assign _zz_927 = _zz_9706[35 : 0];
  assign _zz_929 = 1'b1;
  assign _zz_2073 = _zz_9707;
  assign _zz_2074 = _zz_9715;
  assign _zz_930 = 1'b1;
  assign _zz_2075 = _zz_9723;
  assign _zz_2076 = _zz_9731;
  assign _zz_933 = ($signed(_zz_9739) * $signed(data_mid_5_58_real));
  assign _zz_2077 = _zz_9740;
  assign _zz_931 = _zz_9743[35 : 0];
  assign _zz_2078 = _zz_9744;
  assign _zz_932 = _zz_9747[35 : 0];
  assign _zz_934 = 1'b1;
  assign _zz_2079 = _zz_9748;
  assign _zz_2080 = _zz_9756;
  assign _zz_935 = 1'b1;
  assign _zz_2081 = _zz_9764;
  assign _zz_2082 = _zz_9772;
  assign _zz_938 = ($signed(_zz_9780) * $signed(data_mid_5_59_real));
  assign _zz_2083 = _zz_9781;
  assign _zz_936 = _zz_9784[35 : 0];
  assign _zz_2084 = _zz_9785;
  assign _zz_937 = _zz_9788[35 : 0];
  assign _zz_939 = 1'b1;
  assign _zz_2085 = _zz_9789;
  assign _zz_2086 = _zz_9797;
  assign _zz_940 = 1'b1;
  assign _zz_2087 = _zz_9805;
  assign _zz_2088 = _zz_9813;
  assign _zz_943 = ($signed(_zz_9821) * $signed(data_mid_5_60_real));
  assign _zz_2089 = _zz_9822;
  assign _zz_941 = _zz_9825[35 : 0];
  assign _zz_2090 = _zz_9826;
  assign _zz_942 = _zz_9829[35 : 0];
  assign _zz_944 = 1'b1;
  assign _zz_2091 = _zz_9830;
  assign _zz_2092 = _zz_9838;
  assign _zz_945 = 1'b1;
  assign _zz_2093 = _zz_9846;
  assign _zz_2094 = _zz_9854;
  assign _zz_948 = ($signed(_zz_9862) * $signed(data_mid_5_61_real));
  assign _zz_2095 = _zz_9863;
  assign _zz_946 = _zz_9866[35 : 0];
  assign _zz_2096 = _zz_9867;
  assign _zz_947 = _zz_9870[35 : 0];
  assign _zz_949 = 1'b1;
  assign _zz_2097 = _zz_9871;
  assign _zz_2098 = _zz_9879;
  assign _zz_950 = 1'b1;
  assign _zz_2099 = _zz_9887;
  assign _zz_2100 = _zz_9895;
  assign _zz_953 = ($signed(_zz_9903) * $signed(data_mid_5_62_real));
  assign _zz_2101 = _zz_9904;
  assign _zz_951 = _zz_9907[35 : 0];
  assign _zz_2102 = _zz_9908;
  assign _zz_952 = _zz_9911[35 : 0];
  assign _zz_954 = 1'b1;
  assign _zz_2103 = _zz_9912;
  assign _zz_2104 = _zz_9920;
  assign _zz_955 = 1'b1;
  assign _zz_2105 = _zz_9928;
  assign _zz_2106 = _zz_9936;
  assign _zz_958 = ($signed(_zz_9944) * $signed(data_mid_5_63_real));
  assign _zz_2107 = _zz_9945;
  assign _zz_956 = _zz_9948[35 : 0];
  assign _zz_2108 = _zz_9949;
  assign _zz_957 = _zz_9952[35 : 0];
  assign _zz_959 = 1'b1;
  assign _zz_2109 = _zz_9953;
  assign _zz_2110 = _zz_9961;
  assign _zz_960 = 1'b1;
  assign _zz_2111 = _zz_9969;
  assign _zz_2112 = _zz_9977;
  assign fft_row_valid = io_data_in_valid_delay_8;
  assign fft_row_payload_0_real = data_mid_6_0_real;
  assign fft_row_payload_0_imag = data_mid_6_0_imag;
  assign fft_row_payload_1_real = data_mid_6_1_real;
  assign fft_row_payload_1_imag = data_mid_6_1_imag;
  assign fft_row_payload_2_real = data_mid_6_2_real;
  assign fft_row_payload_2_imag = data_mid_6_2_imag;
  assign fft_row_payload_3_real = data_mid_6_3_real;
  assign fft_row_payload_3_imag = data_mid_6_3_imag;
  assign fft_row_payload_4_real = data_mid_6_4_real;
  assign fft_row_payload_4_imag = data_mid_6_4_imag;
  assign fft_row_payload_5_real = data_mid_6_5_real;
  assign fft_row_payload_5_imag = data_mid_6_5_imag;
  assign fft_row_payload_6_real = data_mid_6_6_real;
  assign fft_row_payload_6_imag = data_mid_6_6_imag;
  assign fft_row_payload_7_real = data_mid_6_7_real;
  assign fft_row_payload_7_imag = data_mid_6_7_imag;
  assign fft_row_payload_8_real = data_mid_6_8_real;
  assign fft_row_payload_8_imag = data_mid_6_8_imag;
  assign fft_row_payload_9_real = data_mid_6_9_real;
  assign fft_row_payload_9_imag = data_mid_6_9_imag;
  assign fft_row_payload_10_real = data_mid_6_10_real;
  assign fft_row_payload_10_imag = data_mid_6_10_imag;
  assign fft_row_payload_11_real = data_mid_6_11_real;
  assign fft_row_payload_11_imag = data_mid_6_11_imag;
  assign fft_row_payload_12_real = data_mid_6_12_real;
  assign fft_row_payload_12_imag = data_mid_6_12_imag;
  assign fft_row_payload_13_real = data_mid_6_13_real;
  assign fft_row_payload_13_imag = data_mid_6_13_imag;
  assign fft_row_payload_14_real = data_mid_6_14_real;
  assign fft_row_payload_14_imag = data_mid_6_14_imag;
  assign fft_row_payload_15_real = data_mid_6_15_real;
  assign fft_row_payload_15_imag = data_mid_6_15_imag;
  assign fft_row_payload_16_real = data_mid_6_16_real;
  assign fft_row_payload_16_imag = data_mid_6_16_imag;
  assign fft_row_payload_17_real = data_mid_6_17_real;
  assign fft_row_payload_17_imag = data_mid_6_17_imag;
  assign fft_row_payload_18_real = data_mid_6_18_real;
  assign fft_row_payload_18_imag = data_mid_6_18_imag;
  assign fft_row_payload_19_real = data_mid_6_19_real;
  assign fft_row_payload_19_imag = data_mid_6_19_imag;
  assign fft_row_payload_20_real = data_mid_6_20_real;
  assign fft_row_payload_20_imag = data_mid_6_20_imag;
  assign fft_row_payload_21_real = data_mid_6_21_real;
  assign fft_row_payload_21_imag = data_mid_6_21_imag;
  assign fft_row_payload_22_real = data_mid_6_22_real;
  assign fft_row_payload_22_imag = data_mid_6_22_imag;
  assign fft_row_payload_23_real = data_mid_6_23_real;
  assign fft_row_payload_23_imag = data_mid_6_23_imag;
  assign fft_row_payload_24_real = data_mid_6_24_real;
  assign fft_row_payload_24_imag = data_mid_6_24_imag;
  assign fft_row_payload_25_real = data_mid_6_25_real;
  assign fft_row_payload_25_imag = data_mid_6_25_imag;
  assign fft_row_payload_26_real = data_mid_6_26_real;
  assign fft_row_payload_26_imag = data_mid_6_26_imag;
  assign fft_row_payload_27_real = data_mid_6_27_real;
  assign fft_row_payload_27_imag = data_mid_6_27_imag;
  assign fft_row_payload_28_real = data_mid_6_28_real;
  assign fft_row_payload_28_imag = data_mid_6_28_imag;
  assign fft_row_payload_29_real = data_mid_6_29_real;
  assign fft_row_payload_29_imag = data_mid_6_29_imag;
  assign fft_row_payload_30_real = data_mid_6_30_real;
  assign fft_row_payload_30_imag = data_mid_6_30_imag;
  assign fft_row_payload_31_real = data_mid_6_31_real;
  assign fft_row_payload_31_imag = data_mid_6_31_imag;
  assign fft_row_payload_32_real = data_mid_6_32_real;
  assign fft_row_payload_32_imag = data_mid_6_32_imag;
  assign fft_row_payload_33_real = data_mid_6_33_real;
  assign fft_row_payload_33_imag = data_mid_6_33_imag;
  assign fft_row_payload_34_real = data_mid_6_34_real;
  assign fft_row_payload_34_imag = data_mid_6_34_imag;
  assign fft_row_payload_35_real = data_mid_6_35_real;
  assign fft_row_payload_35_imag = data_mid_6_35_imag;
  assign fft_row_payload_36_real = data_mid_6_36_real;
  assign fft_row_payload_36_imag = data_mid_6_36_imag;
  assign fft_row_payload_37_real = data_mid_6_37_real;
  assign fft_row_payload_37_imag = data_mid_6_37_imag;
  assign fft_row_payload_38_real = data_mid_6_38_real;
  assign fft_row_payload_38_imag = data_mid_6_38_imag;
  assign fft_row_payload_39_real = data_mid_6_39_real;
  assign fft_row_payload_39_imag = data_mid_6_39_imag;
  assign fft_row_payload_40_real = data_mid_6_40_real;
  assign fft_row_payload_40_imag = data_mid_6_40_imag;
  assign fft_row_payload_41_real = data_mid_6_41_real;
  assign fft_row_payload_41_imag = data_mid_6_41_imag;
  assign fft_row_payload_42_real = data_mid_6_42_real;
  assign fft_row_payload_42_imag = data_mid_6_42_imag;
  assign fft_row_payload_43_real = data_mid_6_43_real;
  assign fft_row_payload_43_imag = data_mid_6_43_imag;
  assign fft_row_payload_44_real = data_mid_6_44_real;
  assign fft_row_payload_44_imag = data_mid_6_44_imag;
  assign fft_row_payload_45_real = data_mid_6_45_real;
  assign fft_row_payload_45_imag = data_mid_6_45_imag;
  assign fft_row_payload_46_real = data_mid_6_46_real;
  assign fft_row_payload_46_imag = data_mid_6_46_imag;
  assign fft_row_payload_47_real = data_mid_6_47_real;
  assign fft_row_payload_47_imag = data_mid_6_47_imag;
  assign fft_row_payload_48_real = data_mid_6_48_real;
  assign fft_row_payload_48_imag = data_mid_6_48_imag;
  assign fft_row_payload_49_real = data_mid_6_49_real;
  assign fft_row_payload_49_imag = data_mid_6_49_imag;
  assign fft_row_payload_50_real = data_mid_6_50_real;
  assign fft_row_payload_50_imag = data_mid_6_50_imag;
  assign fft_row_payload_51_real = data_mid_6_51_real;
  assign fft_row_payload_51_imag = data_mid_6_51_imag;
  assign fft_row_payload_52_real = data_mid_6_52_real;
  assign fft_row_payload_52_imag = data_mid_6_52_imag;
  assign fft_row_payload_53_real = data_mid_6_53_real;
  assign fft_row_payload_53_imag = data_mid_6_53_imag;
  assign fft_row_payload_54_real = data_mid_6_54_real;
  assign fft_row_payload_54_imag = data_mid_6_54_imag;
  assign fft_row_payload_55_real = data_mid_6_55_real;
  assign fft_row_payload_55_imag = data_mid_6_55_imag;
  assign fft_row_payload_56_real = data_mid_6_56_real;
  assign fft_row_payload_56_imag = data_mid_6_56_imag;
  assign fft_row_payload_57_real = data_mid_6_57_real;
  assign fft_row_payload_57_imag = data_mid_6_57_imag;
  assign fft_row_payload_58_real = data_mid_6_58_real;
  assign fft_row_payload_58_imag = data_mid_6_58_imag;
  assign fft_row_payload_59_real = data_mid_6_59_real;
  assign fft_row_payload_59_imag = data_mid_6_59_imag;
  assign fft_row_payload_60_real = data_mid_6_60_real;
  assign fft_row_payload_60_imag = data_mid_6_60_imag;
  assign fft_row_payload_61_real = data_mid_6_61_real;
  assign fft_row_payload_61_imag = data_mid_6_61_imag;
  assign fft_row_payload_62_real = data_mid_6_62_real;
  assign fft_row_payload_62_imag = data_mid_6_62_imag;
  assign fft_row_payload_63_real = data_mid_6_63_real;
  assign fft_row_payload_63_imag = data_mid_6_63_imag;
  always @ (posedge clk) begin
    if(io_data_in_valid)begin
      data_in_0_real <= io_data_in_payload_0_real;
      data_in_0_imag <= io_data_in_payload_0_imag;
      data_in_1_real <= io_data_in_payload_1_real;
      data_in_1_imag <= io_data_in_payload_1_imag;
      data_in_2_real <= io_data_in_payload_2_real;
      data_in_2_imag <= io_data_in_payload_2_imag;
      data_in_3_real <= io_data_in_payload_3_real;
      data_in_3_imag <= io_data_in_payload_3_imag;
      data_in_4_real <= io_data_in_payload_4_real;
      data_in_4_imag <= io_data_in_payload_4_imag;
      data_in_5_real <= io_data_in_payload_5_real;
      data_in_5_imag <= io_data_in_payload_5_imag;
      data_in_6_real <= io_data_in_payload_6_real;
      data_in_6_imag <= io_data_in_payload_6_imag;
      data_in_7_real <= io_data_in_payload_7_real;
      data_in_7_imag <= io_data_in_payload_7_imag;
      data_in_8_real <= io_data_in_payload_8_real;
      data_in_8_imag <= io_data_in_payload_8_imag;
      data_in_9_real <= io_data_in_payload_9_real;
      data_in_9_imag <= io_data_in_payload_9_imag;
      data_in_10_real <= io_data_in_payload_10_real;
      data_in_10_imag <= io_data_in_payload_10_imag;
      data_in_11_real <= io_data_in_payload_11_real;
      data_in_11_imag <= io_data_in_payload_11_imag;
      data_in_12_real <= io_data_in_payload_12_real;
      data_in_12_imag <= io_data_in_payload_12_imag;
      data_in_13_real <= io_data_in_payload_13_real;
      data_in_13_imag <= io_data_in_payload_13_imag;
      data_in_14_real <= io_data_in_payload_14_real;
      data_in_14_imag <= io_data_in_payload_14_imag;
      data_in_15_real <= io_data_in_payload_15_real;
      data_in_15_imag <= io_data_in_payload_15_imag;
      data_in_16_real <= io_data_in_payload_16_real;
      data_in_16_imag <= io_data_in_payload_16_imag;
      data_in_17_real <= io_data_in_payload_17_real;
      data_in_17_imag <= io_data_in_payload_17_imag;
      data_in_18_real <= io_data_in_payload_18_real;
      data_in_18_imag <= io_data_in_payload_18_imag;
      data_in_19_real <= io_data_in_payload_19_real;
      data_in_19_imag <= io_data_in_payload_19_imag;
      data_in_20_real <= io_data_in_payload_20_real;
      data_in_20_imag <= io_data_in_payload_20_imag;
      data_in_21_real <= io_data_in_payload_21_real;
      data_in_21_imag <= io_data_in_payload_21_imag;
      data_in_22_real <= io_data_in_payload_22_real;
      data_in_22_imag <= io_data_in_payload_22_imag;
      data_in_23_real <= io_data_in_payload_23_real;
      data_in_23_imag <= io_data_in_payload_23_imag;
      data_in_24_real <= io_data_in_payload_24_real;
      data_in_24_imag <= io_data_in_payload_24_imag;
      data_in_25_real <= io_data_in_payload_25_real;
      data_in_25_imag <= io_data_in_payload_25_imag;
      data_in_26_real <= io_data_in_payload_26_real;
      data_in_26_imag <= io_data_in_payload_26_imag;
      data_in_27_real <= io_data_in_payload_27_real;
      data_in_27_imag <= io_data_in_payload_27_imag;
      data_in_28_real <= io_data_in_payload_28_real;
      data_in_28_imag <= io_data_in_payload_28_imag;
      data_in_29_real <= io_data_in_payload_29_real;
      data_in_29_imag <= io_data_in_payload_29_imag;
      data_in_30_real <= io_data_in_payload_30_real;
      data_in_30_imag <= io_data_in_payload_30_imag;
      data_in_31_real <= io_data_in_payload_31_real;
      data_in_31_imag <= io_data_in_payload_31_imag;
      data_in_32_real <= io_data_in_payload_32_real;
      data_in_32_imag <= io_data_in_payload_32_imag;
      data_in_33_real <= io_data_in_payload_33_real;
      data_in_33_imag <= io_data_in_payload_33_imag;
      data_in_34_real <= io_data_in_payload_34_real;
      data_in_34_imag <= io_data_in_payload_34_imag;
      data_in_35_real <= io_data_in_payload_35_real;
      data_in_35_imag <= io_data_in_payload_35_imag;
      data_in_36_real <= io_data_in_payload_36_real;
      data_in_36_imag <= io_data_in_payload_36_imag;
      data_in_37_real <= io_data_in_payload_37_real;
      data_in_37_imag <= io_data_in_payload_37_imag;
      data_in_38_real <= io_data_in_payload_38_real;
      data_in_38_imag <= io_data_in_payload_38_imag;
      data_in_39_real <= io_data_in_payload_39_real;
      data_in_39_imag <= io_data_in_payload_39_imag;
      data_in_40_real <= io_data_in_payload_40_real;
      data_in_40_imag <= io_data_in_payload_40_imag;
      data_in_41_real <= io_data_in_payload_41_real;
      data_in_41_imag <= io_data_in_payload_41_imag;
      data_in_42_real <= io_data_in_payload_42_real;
      data_in_42_imag <= io_data_in_payload_42_imag;
      data_in_43_real <= io_data_in_payload_43_real;
      data_in_43_imag <= io_data_in_payload_43_imag;
      data_in_44_real <= io_data_in_payload_44_real;
      data_in_44_imag <= io_data_in_payload_44_imag;
      data_in_45_real <= io_data_in_payload_45_real;
      data_in_45_imag <= io_data_in_payload_45_imag;
      data_in_46_real <= io_data_in_payload_46_real;
      data_in_46_imag <= io_data_in_payload_46_imag;
      data_in_47_real <= io_data_in_payload_47_real;
      data_in_47_imag <= io_data_in_payload_47_imag;
      data_in_48_real <= io_data_in_payload_48_real;
      data_in_48_imag <= io_data_in_payload_48_imag;
      data_in_49_real <= io_data_in_payload_49_real;
      data_in_49_imag <= io_data_in_payload_49_imag;
      data_in_50_real <= io_data_in_payload_50_real;
      data_in_50_imag <= io_data_in_payload_50_imag;
      data_in_51_real <= io_data_in_payload_51_real;
      data_in_51_imag <= io_data_in_payload_51_imag;
      data_in_52_real <= io_data_in_payload_52_real;
      data_in_52_imag <= io_data_in_payload_52_imag;
      data_in_53_real <= io_data_in_payload_53_real;
      data_in_53_imag <= io_data_in_payload_53_imag;
      data_in_54_real <= io_data_in_payload_54_real;
      data_in_54_imag <= io_data_in_payload_54_imag;
      data_in_55_real <= io_data_in_payload_55_real;
      data_in_55_imag <= io_data_in_payload_55_imag;
      data_in_56_real <= io_data_in_payload_56_real;
      data_in_56_imag <= io_data_in_payload_56_imag;
      data_in_57_real <= io_data_in_payload_57_real;
      data_in_57_imag <= io_data_in_payload_57_imag;
      data_in_58_real <= io_data_in_payload_58_real;
      data_in_58_imag <= io_data_in_payload_58_imag;
      data_in_59_real <= io_data_in_payload_59_real;
      data_in_59_imag <= io_data_in_payload_59_imag;
      data_in_60_real <= io_data_in_payload_60_real;
      data_in_60_imag <= io_data_in_payload_60_imag;
      data_in_61_real <= io_data_in_payload_61_real;
      data_in_61_imag <= io_data_in_payload_61_imag;
      data_in_62_real <= io_data_in_payload_62_real;
      data_in_62_imag <= io_data_in_payload_62_imag;
      data_in_63_real <= io_data_in_payload_63_real;
      data_in_63_imag <= io_data_in_payload_63_imag;
    end
    data_mid_0_0_real <= data_reorder_0_real;
    data_mid_0_0_imag <= data_reorder_0_imag;
    data_mid_0_1_real <= data_reorder_1_real;
    data_mid_0_1_imag <= data_reorder_1_imag;
    data_mid_0_2_real <= data_reorder_2_real;
    data_mid_0_2_imag <= data_reorder_2_imag;
    data_mid_0_3_real <= data_reorder_3_real;
    data_mid_0_3_imag <= data_reorder_3_imag;
    data_mid_0_4_real <= data_reorder_4_real;
    data_mid_0_4_imag <= data_reorder_4_imag;
    data_mid_0_5_real <= data_reorder_5_real;
    data_mid_0_5_imag <= data_reorder_5_imag;
    data_mid_0_6_real <= data_reorder_6_real;
    data_mid_0_6_imag <= data_reorder_6_imag;
    data_mid_0_7_real <= data_reorder_7_real;
    data_mid_0_7_imag <= data_reorder_7_imag;
    data_mid_0_8_real <= data_reorder_8_real;
    data_mid_0_8_imag <= data_reorder_8_imag;
    data_mid_0_9_real <= data_reorder_9_real;
    data_mid_0_9_imag <= data_reorder_9_imag;
    data_mid_0_10_real <= data_reorder_10_real;
    data_mid_0_10_imag <= data_reorder_10_imag;
    data_mid_0_11_real <= data_reorder_11_real;
    data_mid_0_11_imag <= data_reorder_11_imag;
    data_mid_0_12_real <= data_reorder_12_real;
    data_mid_0_12_imag <= data_reorder_12_imag;
    data_mid_0_13_real <= data_reorder_13_real;
    data_mid_0_13_imag <= data_reorder_13_imag;
    data_mid_0_14_real <= data_reorder_14_real;
    data_mid_0_14_imag <= data_reorder_14_imag;
    data_mid_0_15_real <= data_reorder_15_real;
    data_mid_0_15_imag <= data_reorder_15_imag;
    data_mid_0_16_real <= data_reorder_16_real;
    data_mid_0_16_imag <= data_reorder_16_imag;
    data_mid_0_17_real <= data_reorder_17_real;
    data_mid_0_17_imag <= data_reorder_17_imag;
    data_mid_0_18_real <= data_reorder_18_real;
    data_mid_0_18_imag <= data_reorder_18_imag;
    data_mid_0_19_real <= data_reorder_19_real;
    data_mid_0_19_imag <= data_reorder_19_imag;
    data_mid_0_20_real <= data_reorder_20_real;
    data_mid_0_20_imag <= data_reorder_20_imag;
    data_mid_0_21_real <= data_reorder_21_real;
    data_mid_0_21_imag <= data_reorder_21_imag;
    data_mid_0_22_real <= data_reorder_22_real;
    data_mid_0_22_imag <= data_reorder_22_imag;
    data_mid_0_23_real <= data_reorder_23_real;
    data_mid_0_23_imag <= data_reorder_23_imag;
    data_mid_0_24_real <= data_reorder_24_real;
    data_mid_0_24_imag <= data_reorder_24_imag;
    data_mid_0_25_real <= data_reorder_25_real;
    data_mid_0_25_imag <= data_reorder_25_imag;
    data_mid_0_26_real <= data_reorder_26_real;
    data_mid_0_26_imag <= data_reorder_26_imag;
    data_mid_0_27_real <= data_reorder_27_real;
    data_mid_0_27_imag <= data_reorder_27_imag;
    data_mid_0_28_real <= data_reorder_28_real;
    data_mid_0_28_imag <= data_reorder_28_imag;
    data_mid_0_29_real <= data_reorder_29_real;
    data_mid_0_29_imag <= data_reorder_29_imag;
    data_mid_0_30_real <= data_reorder_30_real;
    data_mid_0_30_imag <= data_reorder_30_imag;
    data_mid_0_31_real <= data_reorder_31_real;
    data_mid_0_31_imag <= data_reorder_31_imag;
    data_mid_0_32_real <= data_reorder_32_real;
    data_mid_0_32_imag <= data_reorder_32_imag;
    data_mid_0_33_real <= data_reorder_33_real;
    data_mid_0_33_imag <= data_reorder_33_imag;
    data_mid_0_34_real <= data_reorder_34_real;
    data_mid_0_34_imag <= data_reorder_34_imag;
    data_mid_0_35_real <= data_reorder_35_real;
    data_mid_0_35_imag <= data_reorder_35_imag;
    data_mid_0_36_real <= data_reorder_36_real;
    data_mid_0_36_imag <= data_reorder_36_imag;
    data_mid_0_37_real <= data_reorder_37_real;
    data_mid_0_37_imag <= data_reorder_37_imag;
    data_mid_0_38_real <= data_reorder_38_real;
    data_mid_0_38_imag <= data_reorder_38_imag;
    data_mid_0_39_real <= data_reorder_39_real;
    data_mid_0_39_imag <= data_reorder_39_imag;
    data_mid_0_40_real <= data_reorder_40_real;
    data_mid_0_40_imag <= data_reorder_40_imag;
    data_mid_0_41_real <= data_reorder_41_real;
    data_mid_0_41_imag <= data_reorder_41_imag;
    data_mid_0_42_real <= data_reorder_42_real;
    data_mid_0_42_imag <= data_reorder_42_imag;
    data_mid_0_43_real <= data_reorder_43_real;
    data_mid_0_43_imag <= data_reorder_43_imag;
    data_mid_0_44_real <= data_reorder_44_real;
    data_mid_0_44_imag <= data_reorder_44_imag;
    data_mid_0_45_real <= data_reorder_45_real;
    data_mid_0_45_imag <= data_reorder_45_imag;
    data_mid_0_46_real <= data_reorder_46_real;
    data_mid_0_46_imag <= data_reorder_46_imag;
    data_mid_0_47_real <= data_reorder_47_real;
    data_mid_0_47_imag <= data_reorder_47_imag;
    data_mid_0_48_real <= data_reorder_48_real;
    data_mid_0_48_imag <= data_reorder_48_imag;
    data_mid_0_49_real <= data_reorder_49_real;
    data_mid_0_49_imag <= data_reorder_49_imag;
    data_mid_0_50_real <= data_reorder_50_real;
    data_mid_0_50_imag <= data_reorder_50_imag;
    data_mid_0_51_real <= data_reorder_51_real;
    data_mid_0_51_imag <= data_reorder_51_imag;
    data_mid_0_52_real <= data_reorder_52_real;
    data_mid_0_52_imag <= data_reorder_52_imag;
    data_mid_0_53_real <= data_reorder_53_real;
    data_mid_0_53_imag <= data_reorder_53_imag;
    data_mid_0_54_real <= data_reorder_54_real;
    data_mid_0_54_imag <= data_reorder_54_imag;
    data_mid_0_55_real <= data_reorder_55_real;
    data_mid_0_55_imag <= data_reorder_55_imag;
    data_mid_0_56_real <= data_reorder_56_real;
    data_mid_0_56_imag <= data_reorder_56_imag;
    data_mid_0_57_real <= data_reorder_57_real;
    data_mid_0_57_imag <= data_reorder_57_imag;
    data_mid_0_58_real <= data_reorder_58_real;
    data_mid_0_58_imag <= data_reorder_58_imag;
    data_mid_0_59_real <= data_reorder_59_real;
    data_mid_0_59_imag <= data_reorder_59_imag;
    data_mid_0_60_real <= data_reorder_60_real;
    data_mid_0_60_imag <= data_reorder_60_imag;
    data_mid_0_61_real <= data_reorder_61_real;
    data_mid_0_61_imag <= data_reorder_61_imag;
    data_mid_0_62_real <= data_reorder_62_real;
    data_mid_0_62_imag <= data_reorder_62_imag;
    data_mid_0_63_real <= data_reorder_63_real;
    data_mid_0_63_imag <= data_reorder_63_imag;
    data_mid_1_1_real <= _zz_2129[17 : 0];
    data_mid_1_1_imag <= _zz_2137[17 : 0];
    data_mid_1_0_real <= _zz_2145[17 : 0];
    data_mid_1_0_imag <= _zz_2153[17 : 0];
    data_mid_1_3_real <= _zz_2170[17 : 0];
    data_mid_1_3_imag <= _zz_2178[17 : 0];
    data_mid_1_2_real <= _zz_2186[17 : 0];
    data_mid_1_2_imag <= _zz_2194[17 : 0];
    data_mid_1_5_real <= _zz_2211[17 : 0];
    data_mid_1_5_imag <= _zz_2219[17 : 0];
    data_mid_1_4_real <= _zz_2227[17 : 0];
    data_mid_1_4_imag <= _zz_2235[17 : 0];
    data_mid_1_7_real <= _zz_2252[17 : 0];
    data_mid_1_7_imag <= _zz_2260[17 : 0];
    data_mid_1_6_real <= _zz_2268[17 : 0];
    data_mid_1_6_imag <= _zz_2276[17 : 0];
    data_mid_1_9_real <= _zz_2293[17 : 0];
    data_mid_1_9_imag <= _zz_2301[17 : 0];
    data_mid_1_8_real <= _zz_2309[17 : 0];
    data_mid_1_8_imag <= _zz_2317[17 : 0];
    data_mid_1_11_real <= _zz_2334[17 : 0];
    data_mid_1_11_imag <= _zz_2342[17 : 0];
    data_mid_1_10_real <= _zz_2350[17 : 0];
    data_mid_1_10_imag <= _zz_2358[17 : 0];
    data_mid_1_13_real <= _zz_2375[17 : 0];
    data_mid_1_13_imag <= _zz_2383[17 : 0];
    data_mid_1_12_real <= _zz_2391[17 : 0];
    data_mid_1_12_imag <= _zz_2399[17 : 0];
    data_mid_1_15_real <= _zz_2416[17 : 0];
    data_mid_1_15_imag <= _zz_2424[17 : 0];
    data_mid_1_14_real <= _zz_2432[17 : 0];
    data_mid_1_14_imag <= _zz_2440[17 : 0];
    data_mid_1_17_real <= _zz_2457[17 : 0];
    data_mid_1_17_imag <= _zz_2465[17 : 0];
    data_mid_1_16_real <= _zz_2473[17 : 0];
    data_mid_1_16_imag <= _zz_2481[17 : 0];
    data_mid_1_19_real <= _zz_2498[17 : 0];
    data_mid_1_19_imag <= _zz_2506[17 : 0];
    data_mid_1_18_real <= _zz_2514[17 : 0];
    data_mid_1_18_imag <= _zz_2522[17 : 0];
    data_mid_1_21_real <= _zz_2539[17 : 0];
    data_mid_1_21_imag <= _zz_2547[17 : 0];
    data_mid_1_20_real <= _zz_2555[17 : 0];
    data_mid_1_20_imag <= _zz_2563[17 : 0];
    data_mid_1_23_real <= _zz_2580[17 : 0];
    data_mid_1_23_imag <= _zz_2588[17 : 0];
    data_mid_1_22_real <= _zz_2596[17 : 0];
    data_mid_1_22_imag <= _zz_2604[17 : 0];
    data_mid_1_25_real <= _zz_2621[17 : 0];
    data_mid_1_25_imag <= _zz_2629[17 : 0];
    data_mid_1_24_real <= _zz_2637[17 : 0];
    data_mid_1_24_imag <= _zz_2645[17 : 0];
    data_mid_1_27_real <= _zz_2662[17 : 0];
    data_mid_1_27_imag <= _zz_2670[17 : 0];
    data_mid_1_26_real <= _zz_2678[17 : 0];
    data_mid_1_26_imag <= _zz_2686[17 : 0];
    data_mid_1_29_real <= _zz_2703[17 : 0];
    data_mid_1_29_imag <= _zz_2711[17 : 0];
    data_mid_1_28_real <= _zz_2719[17 : 0];
    data_mid_1_28_imag <= _zz_2727[17 : 0];
    data_mid_1_31_real <= _zz_2744[17 : 0];
    data_mid_1_31_imag <= _zz_2752[17 : 0];
    data_mid_1_30_real <= _zz_2760[17 : 0];
    data_mid_1_30_imag <= _zz_2768[17 : 0];
    data_mid_1_33_real <= _zz_2785[17 : 0];
    data_mid_1_33_imag <= _zz_2793[17 : 0];
    data_mid_1_32_real <= _zz_2801[17 : 0];
    data_mid_1_32_imag <= _zz_2809[17 : 0];
    data_mid_1_35_real <= _zz_2826[17 : 0];
    data_mid_1_35_imag <= _zz_2834[17 : 0];
    data_mid_1_34_real <= _zz_2842[17 : 0];
    data_mid_1_34_imag <= _zz_2850[17 : 0];
    data_mid_1_37_real <= _zz_2867[17 : 0];
    data_mid_1_37_imag <= _zz_2875[17 : 0];
    data_mid_1_36_real <= _zz_2883[17 : 0];
    data_mid_1_36_imag <= _zz_2891[17 : 0];
    data_mid_1_39_real <= _zz_2908[17 : 0];
    data_mid_1_39_imag <= _zz_2916[17 : 0];
    data_mid_1_38_real <= _zz_2924[17 : 0];
    data_mid_1_38_imag <= _zz_2932[17 : 0];
    data_mid_1_41_real <= _zz_2949[17 : 0];
    data_mid_1_41_imag <= _zz_2957[17 : 0];
    data_mid_1_40_real <= _zz_2965[17 : 0];
    data_mid_1_40_imag <= _zz_2973[17 : 0];
    data_mid_1_43_real <= _zz_2990[17 : 0];
    data_mid_1_43_imag <= _zz_2998[17 : 0];
    data_mid_1_42_real <= _zz_3006[17 : 0];
    data_mid_1_42_imag <= _zz_3014[17 : 0];
    data_mid_1_45_real <= _zz_3031[17 : 0];
    data_mid_1_45_imag <= _zz_3039[17 : 0];
    data_mid_1_44_real <= _zz_3047[17 : 0];
    data_mid_1_44_imag <= _zz_3055[17 : 0];
    data_mid_1_47_real <= _zz_3072[17 : 0];
    data_mid_1_47_imag <= _zz_3080[17 : 0];
    data_mid_1_46_real <= _zz_3088[17 : 0];
    data_mid_1_46_imag <= _zz_3096[17 : 0];
    data_mid_1_49_real <= _zz_3113[17 : 0];
    data_mid_1_49_imag <= _zz_3121[17 : 0];
    data_mid_1_48_real <= _zz_3129[17 : 0];
    data_mid_1_48_imag <= _zz_3137[17 : 0];
    data_mid_1_51_real <= _zz_3154[17 : 0];
    data_mid_1_51_imag <= _zz_3162[17 : 0];
    data_mid_1_50_real <= _zz_3170[17 : 0];
    data_mid_1_50_imag <= _zz_3178[17 : 0];
    data_mid_1_53_real <= _zz_3195[17 : 0];
    data_mid_1_53_imag <= _zz_3203[17 : 0];
    data_mid_1_52_real <= _zz_3211[17 : 0];
    data_mid_1_52_imag <= _zz_3219[17 : 0];
    data_mid_1_55_real <= _zz_3236[17 : 0];
    data_mid_1_55_imag <= _zz_3244[17 : 0];
    data_mid_1_54_real <= _zz_3252[17 : 0];
    data_mid_1_54_imag <= _zz_3260[17 : 0];
    data_mid_1_57_real <= _zz_3277[17 : 0];
    data_mid_1_57_imag <= _zz_3285[17 : 0];
    data_mid_1_56_real <= _zz_3293[17 : 0];
    data_mid_1_56_imag <= _zz_3301[17 : 0];
    data_mid_1_59_real <= _zz_3318[17 : 0];
    data_mid_1_59_imag <= _zz_3326[17 : 0];
    data_mid_1_58_real <= _zz_3334[17 : 0];
    data_mid_1_58_imag <= _zz_3342[17 : 0];
    data_mid_1_61_real <= _zz_3359[17 : 0];
    data_mid_1_61_imag <= _zz_3367[17 : 0];
    data_mid_1_60_real <= _zz_3375[17 : 0];
    data_mid_1_60_imag <= _zz_3383[17 : 0];
    data_mid_1_63_real <= _zz_3400[17 : 0];
    data_mid_1_63_imag <= _zz_3408[17 : 0];
    data_mid_1_62_real <= _zz_3416[17 : 0];
    data_mid_1_62_imag <= _zz_3424[17 : 0];
    data_mid_2_2_real <= _zz_3441[17 : 0];
    data_mid_2_2_imag <= _zz_3449[17 : 0];
    data_mid_2_0_real <= _zz_3457[17 : 0];
    data_mid_2_0_imag <= _zz_3465[17 : 0];
    data_mid_2_3_real <= _zz_3482[17 : 0];
    data_mid_2_3_imag <= _zz_3490[17 : 0];
    data_mid_2_1_real <= _zz_3498[17 : 0];
    data_mid_2_1_imag <= _zz_3506[17 : 0];
    data_mid_2_6_real <= _zz_3523[17 : 0];
    data_mid_2_6_imag <= _zz_3531[17 : 0];
    data_mid_2_4_real <= _zz_3539[17 : 0];
    data_mid_2_4_imag <= _zz_3547[17 : 0];
    data_mid_2_7_real <= _zz_3564[17 : 0];
    data_mid_2_7_imag <= _zz_3572[17 : 0];
    data_mid_2_5_real <= _zz_3580[17 : 0];
    data_mid_2_5_imag <= _zz_3588[17 : 0];
    data_mid_2_10_real <= _zz_3605[17 : 0];
    data_mid_2_10_imag <= _zz_3613[17 : 0];
    data_mid_2_8_real <= _zz_3621[17 : 0];
    data_mid_2_8_imag <= _zz_3629[17 : 0];
    data_mid_2_11_real <= _zz_3646[17 : 0];
    data_mid_2_11_imag <= _zz_3654[17 : 0];
    data_mid_2_9_real <= _zz_3662[17 : 0];
    data_mid_2_9_imag <= _zz_3670[17 : 0];
    data_mid_2_14_real <= _zz_3687[17 : 0];
    data_mid_2_14_imag <= _zz_3695[17 : 0];
    data_mid_2_12_real <= _zz_3703[17 : 0];
    data_mid_2_12_imag <= _zz_3711[17 : 0];
    data_mid_2_15_real <= _zz_3728[17 : 0];
    data_mid_2_15_imag <= _zz_3736[17 : 0];
    data_mid_2_13_real <= _zz_3744[17 : 0];
    data_mid_2_13_imag <= _zz_3752[17 : 0];
    data_mid_2_18_real <= _zz_3769[17 : 0];
    data_mid_2_18_imag <= _zz_3777[17 : 0];
    data_mid_2_16_real <= _zz_3785[17 : 0];
    data_mid_2_16_imag <= _zz_3793[17 : 0];
    data_mid_2_19_real <= _zz_3810[17 : 0];
    data_mid_2_19_imag <= _zz_3818[17 : 0];
    data_mid_2_17_real <= _zz_3826[17 : 0];
    data_mid_2_17_imag <= _zz_3834[17 : 0];
    data_mid_2_22_real <= _zz_3851[17 : 0];
    data_mid_2_22_imag <= _zz_3859[17 : 0];
    data_mid_2_20_real <= _zz_3867[17 : 0];
    data_mid_2_20_imag <= _zz_3875[17 : 0];
    data_mid_2_23_real <= _zz_3892[17 : 0];
    data_mid_2_23_imag <= _zz_3900[17 : 0];
    data_mid_2_21_real <= _zz_3908[17 : 0];
    data_mid_2_21_imag <= _zz_3916[17 : 0];
    data_mid_2_26_real <= _zz_3933[17 : 0];
    data_mid_2_26_imag <= _zz_3941[17 : 0];
    data_mid_2_24_real <= _zz_3949[17 : 0];
    data_mid_2_24_imag <= _zz_3957[17 : 0];
    data_mid_2_27_real <= _zz_3974[17 : 0];
    data_mid_2_27_imag <= _zz_3982[17 : 0];
    data_mid_2_25_real <= _zz_3990[17 : 0];
    data_mid_2_25_imag <= _zz_3998[17 : 0];
    data_mid_2_30_real <= _zz_4015[17 : 0];
    data_mid_2_30_imag <= _zz_4023[17 : 0];
    data_mid_2_28_real <= _zz_4031[17 : 0];
    data_mid_2_28_imag <= _zz_4039[17 : 0];
    data_mid_2_31_real <= _zz_4056[17 : 0];
    data_mid_2_31_imag <= _zz_4064[17 : 0];
    data_mid_2_29_real <= _zz_4072[17 : 0];
    data_mid_2_29_imag <= _zz_4080[17 : 0];
    data_mid_2_34_real <= _zz_4097[17 : 0];
    data_mid_2_34_imag <= _zz_4105[17 : 0];
    data_mid_2_32_real <= _zz_4113[17 : 0];
    data_mid_2_32_imag <= _zz_4121[17 : 0];
    data_mid_2_35_real <= _zz_4138[17 : 0];
    data_mid_2_35_imag <= _zz_4146[17 : 0];
    data_mid_2_33_real <= _zz_4154[17 : 0];
    data_mid_2_33_imag <= _zz_4162[17 : 0];
    data_mid_2_38_real <= _zz_4179[17 : 0];
    data_mid_2_38_imag <= _zz_4187[17 : 0];
    data_mid_2_36_real <= _zz_4195[17 : 0];
    data_mid_2_36_imag <= _zz_4203[17 : 0];
    data_mid_2_39_real <= _zz_4220[17 : 0];
    data_mid_2_39_imag <= _zz_4228[17 : 0];
    data_mid_2_37_real <= _zz_4236[17 : 0];
    data_mid_2_37_imag <= _zz_4244[17 : 0];
    data_mid_2_42_real <= _zz_4261[17 : 0];
    data_mid_2_42_imag <= _zz_4269[17 : 0];
    data_mid_2_40_real <= _zz_4277[17 : 0];
    data_mid_2_40_imag <= _zz_4285[17 : 0];
    data_mid_2_43_real <= _zz_4302[17 : 0];
    data_mid_2_43_imag <= _zz_4310[17 : 0];
    data_mid_2_41_real <= _zz_4318[17 : 0];
    data_mid_2_41_imag <= _zz_4326[17 : 0];
    data_mid_2_46_real <= _zz_4343[17 : 0];
    data_mid_2_46_imag <= _zz_4351[17 : 0];
    data_mid_2_44_real <= _zz_4359[17 : 0];
    data_mid_2_44_imag <= _zz_4367[17 : 0];
    data_mid_2_47_real <= _zz_4384[17 : 0];
    data_mid_2_47_imag <= _zz_4392[17 : 0];
    data_mid_2_45_real <= _zz_4400[17 : 0];
    data_mid_2_45_imag <= _zz_4408[17 : 0];
    data_mid_2_50_real <= _zz_4425[17 : 0];
    data_mid_2_50_imag <= _zz_4433[17 : 0];
    data_mid_2_48_real <= _zz_4441[17 : 0];
    data_mid_2_48_imag <= _zz_4449[17 : 0];
    data_mid_2_51_real <= _zz_4466[17 : 0];
    data_mid_2_51_imag <= _zz_4474[17 : 0];
    data_mid_2_49_real <= _zz_4482[17 : 0];
    data_mid_2_49_imag <= _zz_4490[17 : 0];
    data_mid_2_54_real <= _zz_4507[17 : 0];
    data_mid_2_54_imag <= _zz_4515[17 : 0];
    data_mid_2_52_real <= _zz_4523[17 : 0];
    data_mid_2_52_imag <= _zz_4531[17 : 0];
    data_mid_2_55_real <= _zz_4548[17 : 0];
    data_mid_2_55_imag <= _zz_4556[17 : 0];
    data_mid_2_53_real <= _zz_4564[17 : 0];
    data_mid_2_53_imag <= _zz_4572[17 : 0];
    data_mid_2_58_real <= _zz_4589[17 : 0];
    data_mid_2_58_imag <= _zz_4597[17 : 0];
    data_mid_2_56_real <= _zz_4605[17 : 0];
    data_mid_2_56_imag <= _zz_4613[17 : 0];
    data_mid_2_59_real <= _zz_4630[17 : 0];
    data_mid_2_59_imag <= _zz_4638[17 : 0];
    data_mid_2_57_real <= _zz_4646[17 : 0];
    data_mid_2_57_imag <= _zz_4654[17 : 0];
    data_mid_2_62_real <= _zz_4671[17 : 0];
    data_mid_2_62_imag <= _zz_4679[17 : 0];
    data_mid_2_60_real <= _zz_4687[17 : 0];
    data_mid_2_60_imag <= _zz_4695[17 : 0];
    data_mid_2_63_real <= _zz_4712[17 : 0];
    data_mid_2_63_imag <= _zz_4720[17 : 0];
    data_mid_2_61_real <= _zz_4728[17 : 0];
    data_mid_2_61_imag <= _zz_4736[17 : 0];
    data_mid_3_4_real <= _zz_4753[17 : 0];
    data_mid_3_4_imag <= _zz_4761[17 : 0];
    data_mid_3_0_real <= _zz_4769[17 : 0];
    data_mid_3_0_imag <= _zz_4777[17 : 0];
    data_mid_3_5_real <= _zz_4794[17 : 0];
    data_mid_3_5_imag <= _zz_4802[17 : 0];
    data_mid_3_1_real <= _zz_4810[17 : 0];
    data_mid_3_1_imag <= _zz_4818[17 : 0];
    data_mid_3_6_real <= _zz_4835[17 : 0];
    data_mid_3_6_imag <= _zz_4843[17 : 0];
    data_mid_3_2_real <= _zz_4851[17 : 0];
    data_mid_3_2_imag <= _zz_4859[17 : 0];
    data_mid_3_7_real <= _zz_4876[17 : 0];
    data_mid_3_7_imag <= _zz_4884[17 : 0];
    data_mid_3_3_real <= _zz_4892[17 : 0];
    data_mid_3_3_imag <= _zz_4900[17 : 0];
    data_mid_3_12_real <= _zz_4917[17 : 0];
    data_mid_3_12_imag <= _zz_4925[17 : 0];
    data_mid_3_8_real <= _zz_4933[17 : 0];
    data_mid_3_8_imag <= _zz_4941[17 : 0];
    data_mid_3_13_real <= _zz_4958[17 : 0];
    data_mid_3_13_imag <= _zz_4966[17 : 0];
    data_mid_3_9_real <= _zz_4974[17 : 0];
    data_mid_3_9_imag <= _zz_4982[17 : 0];
    data_mid_3_14_real <= _zz_4999[17 : 0];
    data_mid_3_14_imag <= _zz_5007[17 : 0];
    data_mid_3_10_real <= _zz_5015[17 : 0];
    data_mid_3_10_imag <= _zz_5023[17 : 0];
    data_mid_3_15_real <= _zz_5040[17 : 0];
    data_mid_3_15_imag <= _zz_5048[17 : 0];
    data_mid_3_11_real <= _zz_5056[17 : 0];
    data_mid_3_11_imag <= _zz_5064[17 : 0];
    data_mid_3_20_real <= _zz_5081[17 : 0];
    data_mid_3_20_imag <= _zz_5089[17 : 0];
    data_mid_3_16_real <= _zz_5097[17 : 0];
    data_mid_3_16_imag <= _zz_5105[17 : 0];
    data_mid_3_21_real <= _zz_5122[17 : 0];
    data_mid_3_21_imag <= _zz_5130[17 : 0];
    data_mid_3_17_real <= _zz_5138[17 : 0];
    data_mid_3_17_imag <= _zz_5146[17 : 0];
    data_mid_3_22_real <= _zz_5163[17 : 0];
    data_mid_3_22_imag <= _zz_5171[17 : 0];
    data_mid_3_18_real <= _zz_5179[17 : 0];
    data_mid_3_18_imag <= _zz_5187[17 : 0];
    data_mid_3_23_real <= _zz_5204[17 : 0];
    data_mid_3_23_imag <= _zz_5212[17 : 0];
    data_mid_3_19_real <= _zz_5220[17 : 0];
    data_mid_3_19_imag <= _zz_5228[17 : 0];
    data_mid_3_28_real <= _zz_5245[17 : 0];
    data_mid_3_28_imag <= _zz_5253[17 : 0];
    data_mid_3_24_real <= _zz_5261[17 : 0];
    data_mid_3_24_imag <= _zz_5269[17 : 0];
    data_mid_3_29_real <= _zz_5286[17 : 0];
    data_mid_3_29_imag <= _zz_5294[17 : 0];
    data_mid_3_25_real <= _zz_5302[17 : 0];
    data_mid_3_25_imag <= _zz_5310[17 : 0];
    data_mid_3_30_real <= _zz_5327[17 : 0];
    data_mid_3_30_imag <= _zz_5335[17 : 0];
    data_mid_3_26_real <= _zz_5343[17 : 0];
    data_mid_3_26_imag <= _zz_5351[17 : 0];
    data_mid_3_31_real <= _zz_5368[17 : 0];
    data_mid_3_31_imag <= _zz_5376[17 : 0];
    data_mid_3_27_real <= _zz_5384[17 : 0];
    data_mid_3_27_imag <= _zz_5392[17 : 0];
    data_mid_3_36_real <= _zz_5409[17 : 0];
    data_mid_3_36_imag <= _zz_5417[17 : 0];
    data_mid_3_32_real <= _zz_5425[17 : 0];
    data_mid_3_32_imag <= _zz_5433[17 : 0];
    data_mid_3_37_real <= _zz_5450[17 : 0];
    data_mid_3_37_imag <= _zz_5458[17 : 0];
    data_mid_3_33_real <= _zz_5466[17 : 0];
    data_mid_3_33_imag <= _zz_5474[17 : 0];
    data_mid_3_38_real <= _zz_5491[17 : 0];
    data_mid_3_38_imag <= _zz_5499[17 : 0];
    data_mid_3_34_real <= _zz_5507[17 : 0];
    data_mid_3_34_imag <= _zz_5515[17 : 0];
    data_mid_3_39_real <= _zz_5532[17 : 0];
    data_mid_3_39_imag <= _zz_5540[17 : 0];
    data_mid_3_35_real <= _zz_5548[17 : 0];
    data_mid_3_35_imag <= _zz_5556[17 : 0];
    data_mid_3_44_real <= _zz_5573[17 : 0];
    data_mid_3_44_imag <= _zz_5581[17 : 0];
    data_mid_3_40_real <= _zz_5589[17 : 0];
    data_mid_3_40_imag <= _zz_5597[17 : 0];
    data_mid_3_45_real <= _zz_5614[17 : 0];
    data_mid_3_45_imag <= _zz_5622[17 : 0];
    data_mid_3_41_real <= _zz_5630[17 : 0];
    data_mid_3_41_imag <= _zz_5638[17 : 0];
    data_mid_3_46_real <= _zz_5655[17 : 0];
    data_mid_3_46_imag <= _zz_5663[17 : 0];
    data_mid_3_42_real <= _zz_5671[17 : 0];
    data_mid_3_42_imag <= _zz_5679[17 : 0];
    data_mid_3_47_real <= _zz_5696[17 : 0];
    data_mid_3_47_imag <= _zz_5704[17 : 0];
    data_mid_3_43_real <= _zz_5712[17 : 0];
    data_mid_3_43_imag <= _zz_5720[17 : 0];
    data_mid_3_52_real <= _zz_5737[17 : 0];
    data_mid_3_52_imag <= _zz_5745[17 : 0];
    data_mid_3_48_real <= _zz_5753[17 : 0];
    data_mid_3_48_imag <= _zz_5761[17 : 0];
    data_mid_3_53_real <= _zz_5778[17 : 0];
    data_mid_3_53_imag <= _zz_5786[17 : 0];
    data_mid_3_49_real <= _zz_5794[17 : 0];
    data_mid_3_49_imag <= _zz_5802[17 : 0];
    data_mid_3_54_real <= _zz_5819[17 : 0];
    data_mid_3_54_imag <= _zz_5827[17 : 0];
    data_mid_3_50_real <= _zz_5835[17 : 0];
    data_mid_3_50_imag <= _zz_5843[17 : 0];
    data_mid_3_55_real <= _zz_5860[17 : 0];
    data_mid_3_55_imag <= _zz_5868[17 : 0];
    data_mid_3_51_real <= _zz_5876[17 : 0];
    data_mid_3_51_imag <= _zz_5884[17 : 0];
    data_mid_3_60_real <= _zz_5901[17 : 0];
    data_mid_3_60_imag <= _zz_5909[17 : 0];
    data_mid_3_56_real <= _zz_5917[17 : 0];
    data_mid_3_56_imag <= _zz_5925[17 : 0];
    data_mid_3_61_real <= _zz_5942[17 : 0];
    data_mid_3_61_imag <= _zz_5950[17 : 0];
    data_mid_3_57_real <= _zz_5958[17 : 0];
    data_mid_3_57_imag <= _zz_5966[17 : 0];
    data_mid_3_62_real <= _zz_5983[17 : 0];
    data_mid_3_62_imag <= _zz_5991[17 : 0];
    data_mid_3_58_real <= _zz_5999[17 : 0];
    data_mid_3_58_imag <= _zz_6007[17 : 0];
    data_mid_3_63_real <= _zz_6024[17 : 0];
    data_mid_3_63_imag <= _zz_6032[17 : 0];
    data_mid_3_59_real <= _zz_6040[17 : 0];
    data_mid_3_59_imag <= _zz_6048[17 : 0];
    data_mid_4_8_real <= _zz_6065[17 : 0];
    data_mid_4_8_imag <= _zz_6073[17 : 0];
    data_mid_4_0_real <= _zz_6081[17 : 0];
    data_mid_4_0_imag <= _zz_6089[17 : 0];
    data_mid_4_9_real <= _zz_6106[17 : 0];
    data_mid_4_9_imag <= _zz_6114[17 : 0];
    data_mid_4_1_real <= _zz_6122[17 : 0];
    data_mid_4_1_imag <= _zz_6130[17 : 0];
    data_mid_4_10_real <= _zz_6147[17 : 0];
    data_mid_4_10_imag <= _zz_6155[17 : 0];
    data_mid_4_2_real <= _zz_6163[17 : 0];
    data_mid_4_2_imag <= _zz_6171[17 : 0];
    data_mid_4_11_real <= _zz_6188[17 : 0];
    data_mid_4_11_imag <= _zz_6196[17 : 0];
    data_mid_4_3_real <= _zz_6204[17 : 0];
    data_mid_4_3_imag <= _zz_6212[17 : 0];
    data_mid_4_12_real <= _zz_6229[17 : 0];
    data_mid_4_12_imag <= _zz_6237[17 : 0];
    data_mid_4_4_real <= _zz_6245[17 : 0];
    data_mid_4_4_imag <= _zz_6253[17 : 0];
    data_mid_4_13_real <= _zz_6270[17 : 0];
    data_mid_4_13_imag <= _zz_6278[17 : 0];
    data_mid_4_5_real <= _zz_6286[17 : 0];
    data_mid_4_5_imag <= _zz_6294[17 : 0];
    data_mid_4_14_real <= _zz_6311[17 : 0];
    data_mid_4_14_imag <= _zz_6319[17 : 0];
    data_mid_4_6_real <= _zz_6327[17 : 0];
    data_mid_4_6_imag <= _zz_6335[17 : 0];
    data_mid_4_15_real <= _zz_6352[17 : 0];
    data_mid_4_15_imag <= _zz_6360[17 : 0];
    data_mid_4_7_real <= _zz_6368[17 : 0];
    data_mid_4_7_imag <= _zz_6376[17 : 0];
    data_mid_4_24_real <= _zz_6393[17 : 0];
    data_mid_4_24_imag <= _zz_6401[17 : 0];
    data_mid_4_16_real <= _zz_6409[17 : 0];
    data_mid_4_16_imag <= _zz_6417[17 : 0];
    data_mid_4_25_real <= _zz_6434[17 : 0];
    data_mid_4_25_imag <= _zz_6442[17 : 0];
    data_mid_4_17_real <= _zz_6450[17 : 0];
    data_mid_4_17_imag <= _zz_6458[17 : 0];
    data_mid_4_26_real <= _zz_6475[17 : 0];
    data_mid_4_26_imag <= _zz_6483[17 : 0];
    data_mid_4_18_real <= _zz_6491[17 : 0];
    data_mid_4_18_imag <= _zz_6499[17 : 0];
    data_mid_4_27_real <= _zz_6516[17 : 0];
    data_mid_4_27_imag <= _zz_6524[17 : 0];
    data_mid_4_19_real <= _zz_6532[17 : 0];
    data_mid_4_19_imag <= _zz_6540[17 : 0];
    data_mid_4_28_real <= _zz_6557[17 : 0];
    data_mid_4_28_imag <= _zz_6565[17 : 0];
    data_mid_4_20_real <= _zz_6573[17 : 0];
    data_mid_4_20_imag <= _zz_6581[17 : 0];
    data_mid_4_29_real <= _zz_6598[17 : 0];
    data_mid_4_29_imag <= _zz_6606[17 : 0];
    data_mid_4_21_real <= _zz_6614[17 : 0];
    data_mid_4_21_imag <= _zz_6622[17 : 0];
    data_mid_4_30_real <= _zz_6639[17 : 0];
    data_mid_4_30_imag <= _zz_6647[17 : 0];
    data_mid_4_22_real <= _zz_6655[17 : 0];
    data_mid_4_22_imag <= _zz_6663[17 : 0];
    data_mid_4_31_real <= _zz_6680[17 : 0];
    data_mid_4_31_imag <= _zz_6688[17 : 0];
    data_mid_4_23_real <= _zz_6696[17 : 0];
    data_mid_4_23_imag <= _zz_6704[17 : 0];
    data_mid_4_40_real <= _zz_6721[17 : 0];
    data_mid_4_40_imag <= _zz_6729[17 : 0];
    data_mid_4_32_real <= _zz_6737[17 : 0];
    data_mid_4_32_imag <= _zz_6745[17 : 0];
    data_mid_4_41_real <= _zz_6762[17 : 0];
    data_mid_4_41_imag <= _zz_6770[17 : 0];
    data_mid_4_33_real <= _zz_6778[17 : 0];
    data_mid_4_33_imag <= _zz_6786[17 : 0];
    data_mid_4_42_real <= _zz_6803[17 : 0];
    data_mid_4_42_imag <= _zz_6811[17 : 0];
    data_mid_4_34_real <= _zz_6819[17 : 0];
    data_mid_4_34_imag <= _zz_6827[17 : 0];
    data_mid_4_43_real <= _zz_6844[17 : 0];
    data_mid_4_43_imag <= _zz_6852[17 : 0];
    data_mid_4_35_real <= _zz_6860[17 : 0];
    data_mid_4_35_imag <= _zz_6868[17 : 0];
    data_mid_4_44_real <= _zz_6885[17 : 0];
    data_mid_4_44_imag <= _zz_6893[17 : 0];
    data_mid_4_36_real <= _zz_6901[17 : 0];
    data_mid_4_36_imag <= _zz_6909[17 : 0];
    data_mid_4_45_real <= _zz_6926[17 : 0];
    data_mid_4_45_imag <= _zz_6934[17 : 0];
    data_mid_4_37_real <= _zz_6942[17 : 0];
    data_mid_4_37_imag <= _zz_6950[17 : 0];
    data_mid_4_46_real <= _zz_6967[17 : 0];
    data_mid_4_46_imag <= _zz_6975[17 : 0];
    data_mid_4_38_real <= _zz_6983[17 : 0];
    data_mid_4_38_imag <= _zz_6991[17 : 0];
    data_mid_4_47_real <= _zz_7008[17 : 0];
    data_mid_4_47_imag <= _zz_7016[17 : 0];
    data_mid_4_39_real <= _zz_7024[17 : 0];
    data_mid_4_39_imag <= _zz_7032[17 : 0];
    data_mid_4_56_real <= _zz_7049[17 : 0];
    data_mid_4_56_imag <= _zz_7057[17 : 0];
    data_mid_4_48_real <= _zz_7065[17 : 0];
    data_mid_4_48_imag <= _zz_7073[17 : 0];
    data_mid_4_57_real <= _zz_7090[17 : 0];
    data_mid_4_57_imag <= _zz_7098[17 : 0];
    data_mid_4_49_real <= _zz_7106[17 : 0];
    data_mid_4_49_imag <= _zz_7114[17 : 0];
    data_mid_4_58_real <= _zz_7131[17 : 0];
    data_mid_4_58_imag <= _zz_7139[17 : 0];
    data_mid_4_50_real <= _zz_7147[17 : 0];
    data_mid_4_50_imag <= _zz_7155[17 : 0];
    data_mid_4_59_real <= _zz_7172[17 : 0];
    data_mid_4_59_imag <= _zz_7180[17 : 0];
    data_mid_4_51_real <= _zz_7188[17 : 0];
    data_mid_4_51_imag <= _zz_7196[17 : 0];
    data_mid_4_60_real <= _zz_7213[17 : 0];
    data_mid_4_60_imag <= _zz_7221[17 : 0];
    data_mid_4_52_real <= _zz_7229[17 : 0];
    data_mid_4_52_imag <= _zz_7237[17 : 0];
    data_mid_4_61_real <= _zz_7254[17 : 0];
    data_mid_4_61_imag <= _zz_7262[17 : 0];
    data_mid_4_53_real <= _zz_7270[17 : 0];
    data_mid_4_53_imag <= _zz_7278[17 : 0];
    data_mid_4_62_real <= _zz_7295[17 : 0];
    data_mid_4_62_imag <= _zz_7303[17 : 0];
    data_mid_4_54_real <= _zz_7311[17 : 0];
    data_mid_4_54_imag <= _zz_7319[17 : 0];
    data_mid_4_63_real <= _zz_7336[17 : 0];
    data_mid_4_63_imag <= _zz_7344[17 : 0];
    data_mid_4_55_real <= _zz_7352[17 : 0];
    data_mid_4_55_imag <= _zz_7360[17 : 0];
    data_mid_5_16_real <= _zz_7377[17 : 0];
    data_mid_5_16_imag <= _zz_7385[17 : 0];
    data_mid_5_0_real <= _zz_7393[17 : 0];
    data_mid_5_0_imag <= _zz_7401[17 : 0];
    data_mid_5_17_real <= _zz_7418[17 : 0];
    data_mid_5_17_imag <= _zz_7426[17 : 0];
    data_mid_5_1_real <= _zz_7434[17 : 0];
    data_mid_5_1_imag <= _zz_7442[17 : 0];
    data_mid_5_18_real <= _zz_7459[17 : 0];
    data_mid_5_18_imag <= _zz_7467[17 : 0];
    data_mid_5_2_real <= _zz_7475[17 : 0];
    data_mid_5_2_imag <= _zz_7483[17 : 0];
    data_mid_5_19_real <= _zz_7500[17 : 0];
    data_mid_5_19_imag <= _zz_7508[17 : 0];
    data_mid_5_3_real <= _zz_7516[17 : 0];
    data_mid_5_3_imag <= _zz_7524[17 : 0];
    data_mid_5_20_real <= _zz_7541[17 : 0];
    data_mid_5_20_imag <= _zz_7549[17 : 0];
    data_mid_5_4_real <= _zz_7557[17 : 0];
    data_mid_5_4_imag <= _zz_7565[17 : 0];
    data_mid_5_21_real <= _zz_7582[17 : 0];
    data_mid_5_21_imag <= _zz_7590[17 : 0];
    data_mid_5_5_real <= _zz_7598[17 : 0];
    data_mid_5_5_imag <= _zz_7606[17 : 0];
    data_mid_5_22_real <= _zz_7623[17 : 0];
    data_mid_5_22_imag <= _zz_7631[17 : 0];
    data_mid_5_6_real <= _zz_7639[17 : 0];
    data_mid_5_6_imag <= _zz_7647[17 : 0];
    data_mid_5_23_real <= _zz_7664[17 : 0];
    data_mid_5_23_imag <= _zz_7672[17 : 0];
    data_mid_5_7_real <= _zz_7680[17 : 0];
    data_mid_5_7_imag <= _zz_7688[17 : 0];
    data_mid_5_24_real <= _zz_7705[17 : 0];
    data_mid_5_24_imag <= _zz_7713[17 : 0];
    data_mid_5_8_real <= _zz_7721[17 : 0];
    data_mid_5_8_imag <= _zz_7729[17 : 0];
    data_mid_5_25_real <= _zz_7746[17 : 0];
    data_mid_5_25_imag <= _zz_7754[17 : 0];
    data_mid_5_9_real <= _zz_7762[17 : 0];
    data_mid_5_9_imag <= _zz_7770[17 : 0];
    data_mid_5_26_real <= _zz_7787[17 : 0];
    data_mid_5_26_imag <= _zz_7795[17 : 0];
    data_mid_5_10_real <= _zz_7803[17 : 0];
    data_mid_5_10_imag <= _zz_7811[17 : 0];
    data_mid_5_27_real <= _zz_7828[17 : 0];
    data_mid_5_27_imag <= _zz_7836[17 : 0];
    data_mid_5_11_real <= _zz_7844[17 : 0];
    data_mid_5_11_imag <= _zz_7852[17 : 0];
    data_mid_5_28_real <= _zz_7869[17 : 0];
    data_mid_5_28_imag <= _zz_7877[17 : 0];
    data_mid_5_12_real <= _zz_7885[17 : 0];
    data_mid_5_12_imag <= _zz_7893[17 : 0];
    data_mid_5_29_real <= _zz_7910[17 : 0];
    data_mid_5_29_imag <= _zz_7918[17 : 0];
    data_mid_5_13_real <= _zz_7926[17 : 0];
    data_mid_5_13_imag <= _zz_7934[17 : 0];
    data_mid_5_30_real <= _zz_7951[17 : 0];
    data_mid_5_30_imag <= _zz_7959[17 : 0];
    data_mid_5_14_real <= _zz_7967[17 : 0];
    data_mid_5_14_imag <= _zz_7975[17 : 0];
    data_mid_5_31_real <= _zz_7992[17 : 0];
    data_mid_5_31_imag <= _zz_8000[17 : 0];
    data_mid_5_15_real <= _zz_8008[17 : 0];
    data_mid_5_15_imag <= _zz_8016[17 : 0];
    data_mid_5_48_real <= _zz_8033[17 : 0];
    data_mid_5_48_imag <= _zz_8041[17 : 0];
    data_mid_5_32_real <= _zz_8049[17 : 0];
    data_mid_5_32_imag <= _zz_8057[17 : 0];
    data_mid_5_49_real <= _zz_8074[17 : 0];
    data_mid_5_49_imag <= _zz_8082[17 : 0];
    data_mid_5_33_real <= _zz_8090[17 : 0];
    data_mid_5_33_imag <= _zz_8098[17 : 0];
    data_mid_5_50_real <= _zz_8115[17 : 0];
    data_mid_5_50_imag <= _zz_8123[17 : 0];
    data_mid_5_34_real <= _zz_8131[17 : 0];
    data_mid_5_34_imag <= _zz_8139[17 : 0];
    data_mid_5_51_real <= _zz_8156[17 : 0];
    data_mid_5_51_imag <= _zz_8164[17 : 0];
    data_mid_5_35_real <= _zz_8172[17 : 0];
    data_mid_5_35_imag <= _zz_8180[17 : 0];
    data_mid_5_52_real <= _zz_8197[17 : 0];
    data_mid_5_52_imag <= _zz_8205[17 : 0];
    data_mid_5_36_real <= _zz_8213[17 : 0];
    data_mid_5_36_imag <= _zz_8221[17 : 0];
    data_mid_5_53_real <= _zz_8238[17 : 0];
    data_mid_5_53_imag <= _zz_8246[17 : 0];
    data_mid_5_37_real <= _zz_8254[17 : 0];
    data_mid_5_37_imag <= _zz_8262[17 : 0];
    data_mid_5_54_real <= _zz_8279[17 : 0];
    data_mid_5_54_imag <= _zz_8287[17 : 0];
    data_mid_5_38_real <= _zz_8295[17 : 0];
    data_mid_5_38_imag <= _zz_8303[17 : 0];
    data_mid_5_55_real <= _zz_8320[17 : 0];
    data_mid_5_55_imag <= _zz_8328[17 : 0];
    data_mid_5_39_real <= _zz_8336[17 : 0];
    data_mid_5_39_imag <= _zz_8344[17 : 0];
    data_mid_5_56_real <= _zz_8361[17 : 0];
    data_mid_5_56_imag <= _zz_8369[17 : 0];
    data_mid_5_40_real <= _zz_8377[17 : 0];
    data_mid_5_40_imag <= _zz_8385[17 : 0];
    data_mid_5_57_real <= _zz_8402[17 : 0];
    data_mid_5_57_imag <= _zz_8410[17 : 0];
    data_mid_5_41_real <= _zz_8418[17 : 0];
    data_mid_5_41_imag <= _zz_8426[17 : 0];
    data_mid_5_58_real <= _zz_8443[17 : 0];
    data_mid_5_58_imag <= _zz_8451[17 : 0];
    data_mid_5_42_real <= _zz_8459[17 : 0];
    data_mid_5_42_imag <= _zz_8467[17 : 0];
    data_mid_5_59_real <= _zz_8484[17 : 0];
    data_mid_5_59_imag <= _zz_8492[17 : 0];
    data_mid_5_43_real <= _zz_8500[17 : 0];
    data_mid_5_43_imag <= _zz_8508[17 : 0];
    data_mid_5_60_real <= _zz_8525[17 : 0];
    data_mid_5_60_imag <= _zz_8533[17 : 0];
    data_mid_5_44_real <= _zz_8541[17 : 0];
    data_mid_5_44_imag <= _zz_8549[17 : 0];
    data_mid_5_61_real <= _zz_8566[17 : 0];
    data_mid_5_61_imag <= _zz_8574[17 : 0];
    data_mid_5_45_real <= _zz_8582[17 : 0];
    data_mid_5_45_imag <= _zz_8590[17 : 0];
    data_mid_5_62_real <= _zz_8607[17 : 0];
    data_mid_5_62_imag <= _zz_8615[17 : 0];
    data_mid_5_46_real <= _zz_8623[17 : 0];
    data_mid_5_46_imag <= _zz_8631[17 : 0];
    data_mid_5_63_real <= _zz_8648[17 : 0];
    data_mid_5_63_imag <= _zz_8656[17 : 0];
    data_mid_5_47_real <= _zz_8664[17 : 0];
    data_mid_5_47_imag <= _zz_8672[17 : 0];
    data_mid_6_32_real <= _zz_8689[17 : 0];
    data_mid_6_32_imag <= _zz_8697[17 : 0];
    data_mid_6_0_real <= _zz_8705[17 : 0];
    data_mid_6_0_imag <= _zz_8713[17 : 0];
    data_mid_6_33_real <= _zz_8730[17 : 0];
    data_mid_6_33_imag <= _zz_8738[17 : 0];
    data_mid_6_1_real <= _zz_8746[17 : 0];
    data_mid_6_1_imag <= _zz_8754[17 : 0];
    data_mid_6_34_real <= _zz_8771[17 : 0];
    data_mid_6_34_imag <= _zz_8779[17 : 0];
    data_mid_6_2_real <= _zz_8787[17 : 0];
    data_mid_6_2_imag <= _zz_8795[17 : 0];
    data_mid_6_35_real <= _zz_8812[17 : 0];
    data_mid_6_35_imag <= _zz_8820[17 : 0];
    data_mid_6_3_real <= _zz_8828[17 : 0];
    data_mid_6_3_imag <= _zz_8836[17 : 0];
    data_mid_6_36_real <= _zz_8853[17 : 0];
    data_mid_6_36_imag <= _zz_8861[17 : 0];
    data_mid_6_4_real <= _zz_8869[17 : 0];
    data_mid_6_4_imag <= _zz_8877[17 : 0];
    data_mid_6_37_real <= _zz_8894[17 : 0];
    data_mid_6_37_imag <= _zz_8902[17 : 0];
    data_mid_6_5_real <= _zz_8910[17 : 0];
    data_mid_6_5_imag <= _zz_8918[17 : 0];
    data_mid_6_38_real <= _zz_8935[17 : 0];
    data_mid_6_38_imag <= _zz_8943[17 : 0];
    data_mid_6_6_real <= _zz_8951[17 : 0];
    data_mid_6_6_imag <= _zz_8959[17 : 0];
    data_mid_6_39_real <= _zz_8976[17 : 0];
    data_mid_6_39_imag <= _zz_8984[17 : 0];
    data_mid_6_7_real <= _zz_8992[17 : 0];
    data_mid_6_7_imag <= _zz_9000[17 : 0];
    data_mid_6_40_real <= _zz_9017[17 : 0];
    data_mid_6_40_imag <= _zz_9025[17 : 0];
    data_mid_6_8_real <= _zz_9033[17 : 0];
    data_mid_6_8_imag <= _zz_9041[17 : 0];
    data_mid_6_41_real <= _zz_9058[17 : 0];
    data_mid_6_41_imag <= _zz_9066[17 : 0];
    data_mid_6_9_real <= _zz_9074[17 : 0];
    data_mid_6_9_imag <= _zz_9082[17 : 0];
    data_mid_6_42_real <= _zz_9099[17 : 0];
    data_mid_6_42_imag <= _zz_9107[17 : 0];
    data_mid_6_10_real <= _zz_9115[17 : 0];
    data_mid_6_10_imag <= _zz_9123[17 : 0];
    data_mid_6_43_real <= _zz_9140[17 : 0];
    data_mid_6_43_imag <= _zz_9148[17 : 0];
    data_mid_6_11_real <= _zz_9156[17 : 0];
    data_mid_6_11_imag <= _zz_9164[17 : 0];
    data_mid_6_44_real <= _zz_9181[17 : 0];
    data_mid_6_44_imag <= _zz_9189[17 : 0];
    data_mid_6_12_real <= _zz_9197[17 : 0];
    data_mid_6_12_imag <= _zz_9205[17 : 0];
    data_mid_6_45_real <= _zz_9222[17 : 0];
    data_mid_6_45_imag <= _zz_9230[17 : 0];
    data_mid_6_13_real <= _zz_9238[17 : 0];
    data_mid_6_13_imag <= _zz_9246[17 : 0];
    data_mid_6_46_real <= _zz_9263[17 : 0];
    data_mid_6_46_imag <= _zz_9271[17 : 0];
    data_mid_6_14_real <= _zz_9279[17 : 0];
    data_mid_6_14_imag <= _zz_9287[17 : 0];
    data_mid_6_47_real <= _zz_9304[17 : 0];
    data_mid_6_47_imag <= _zz_9312[17 : 0];
    data_mid_6_15_real <= _zz_9320[17 : 0];
    data_mid_6_15_imag <= _zz_9328[17 : 0];
    data_mid_6_48_real <= _zz_9345[17 : 0];
    data_mid_6_48_imag <= _zz_9353[17 : 0];
    data_mid_6_16_real <= _zz_9361[17 : 0];
    data_mid_6_16_imag <= _zz_9369[17 : 0];
    data_mid_6_49_real <= _zz_9386[17 : 0];
    data_mid_6_49_imag <= _zz_9394[17 : 0];
    data_mid_6_17_real <= _zz_9402[17 : 0];
    data_mid_6_17_imag <= _zz_9410[17 : 0];
    data_mid_6_50_real <= _zz_9427[17 : 0];
    data_mid_6_50_imag <= _zz_9435[17 : 0];
    data_mid_6_18_real <= _zz_9443[17 : 0];
    data_mid_6_18_imag <= _zz_9451[17 : 0];
    data_mid_6_51_real <= _zz_9468[17 : 0];
    data_mid_6_51_imag <= _zz_9476[17 : 0];
    data_mid_6_19_real <= _zz_9484[17 : 0];
    data_mid_6_19_imag <= _zz_9492[17 : 0];
    data_mid_6_52_real <= _zz_9509[17 : 0];
    data_mid_6_52_imag <= _zz_9517[17 : 0];
    data_mid_6_20_real <= _zz_9525[17 : 0];
    data_mid_6_20_imag <= _zz_9533[17 : 0];
    data_mid_6_53_real <= _zz_9550[17 : 0];
    data_mid_6_53_imag <= _zz_9558[17 : 0];
    data_mid_6_21_real <= _zz_9566[17 : 0];
    data_mid_6_21_imag <= _zz_9574[17 : 0];
    data_mid_6_54_real <= _zz_9591[17 : 0];
    data_mid_6_54_imag <= _zz_9599[17 : 0];
    data_mid_6_22_real <= _zz_9607[17 : 0];
    data_mid_6_22_imag <= _zz_9615[17 : 0];
    data_mid_6_55_real <= _zz_9632[17 : 0];
    data_mid_6_55_imag <= _zz_9640[17 : 0];
    data_mid_6_23_real <= _zz_9648[17 : 0];
    data_mid_6_23_imag <= _zz_9656[17 : 0];
    data_mid_6_56_real <= _zz_9673[17 : 0];
    data_mid_6_56_imag <= _zz_9681[17 : 0];
    data_mid_6_24_real <= _zz_9689[17 : 0];
    data_mid_6_24_imag <= _zz_9697[17 : 0];
    data_mid_6_57_real <= _zz_9714[17 : 0];
    data_mid_6_57_imag <= _zz_9722[17 : 0];
    data_mid_6_25_real <= _zz_9730[17 : 0];
    data_mid_6_25_imag <= _zz_9738[17 : 0];
    data_mid_6_58_real <= _zz_9755[17 : 0];
    data_mid_6_58_imag <= _zz_9763[17 : 0];
    data_mid_6_26_real <= _zz_9771[17 : 0];
    data_mid_6_26_imag <= _zz_9779[17 : 0];
    data_mid_6_59_real <= _zz_9796[17 : 0];
    data_mid_6_59_imag <= _zz_9804[17 : 0];
    data_mid_6_27_real <= _zz_9812[17 : 0];
    data_mid_6_27_imag <= _zz_9820[17 : 0];
    data_mid_6_60_real <= _zz_9837[17 : 0];
    data_mid_6_60_imag <= _zz_9845[17 : 0];
    data_mid_6_28_real <= _zz_9853[17 : 0];
    data_mid_6_28_imag <= _zz_9861[17 : 0];
    data_mid_6_61_real <= _zz_9878[17 : 0];
    data_mid_6_61_imag <= _zz_9886[17 : 0];
    data_mid_6_29_real <= _zz_9894[17 : 0];
    data_mid_6_29_imag <= _zz_9902[17 : 0];
    data_mid_6_62_real <= _zz_9919[17 : 0];
    data_mid_6_62_imag <= _zz_9927[17 : 0];
    data_mid_6_30_real <= _zz_9935[17 : 0];
    data_mid_6_30_imag <= _zz_9943[17 : 0];
    data_mid_6_63_real <= _zz_9960[17 : 0];
    data_mid_6_63_imag <= _zz_9968[17 : 0];
    data_mid_6_31_real <= _zz_9976[17 : 0];
    data_mid_6_31_imag <= _zz_9984[17 : 0];
  end

  always @ (posedge clk or posedge reset) begin
    if (reset) begin
      io_data_in_valid_delay_1 <= 1'b0;
      io_data_in_valid_delay_2 <= 1'b0;
      io_data_in_valid_delay_3 <= 1'b0;
      io_data_in_valid_delay_4 <= 1'b0;
      io_data_in_valid_delay_5 <= 1'b0;
      io_data_in_valid_delay_6 <= 1'b0;
      io_data_in_valid_delay_7 <= 1'b0;
      io_data_in_valid_delay_8 <= 1'b0;
    end else begin
      io_data_in_valid_delay_1 <= io_data_in_valid;
      io_data_in_valid_delay_2 <= io_data_in_valid_delay_1;
      io_data_in_valid_delay_3 <= io_data_in_valid_delay_2;
      io_data_in_valid_delay_4 <= io_data_in_valid_delay_3;
      io_data_in_valid_delay_5 <= io_data_in_valid_delay_4;
      io_data_in_valid_delay_6 <= io_data_in_valid_delay_5;
      io_data_in_valid_delay_7 <= io_data_in_valid_delay_6;
      io_data_in_valid_delay_8 <= io_data_in_valid_delay_7;
    end
  end


endmodule

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

//SInt36fixTo26_9_ROUNDTOINF replaced by SInt36fixTo26_9_ROUNDTOINF

module SInt36fixTo26_9_ROUNDTOINF (
  input      [35:0]   din,
  output     [17:0]   dout
);
  wire       [36:0]   _zz_9;
  wire       [36:0]   _zz_10;
  wire       [8:0]    _zz_11;
  wire       [27:0]   _zz_12;
  wire       [27:0]   _zz_13;
  wire       [36:0]   _zz_14;
  wire       [36:0]   _zz_15;
  wire       [36:0]   _zz_16;
  wire       [10:0]   _zz_17;
  wire       [9:0]    _zz_18;
  reg        [27:0]   _zz_1;
  wire       [35:0]   _zz_2;
  wire       [35:0]   _zz_3;
  wire       [35:0]   _zz_4;
  wire       [36:0]   _zz_5;
  wire       [35:0]   _zz_6;
  reg        [27:0]   _zz_7;
  reg        [17:0]   _zz_8;

  assign _zz_9 = {_zz_4[35],_zz_4};
  assign _zz_10 = {_zz_3[35],_zz_3};
  assign _zz_11 = _zz_5[8 : 0];
  assign _zz_12 = _zz_5[36 : 9];
  assign _zz_13 = 28'h0000001;
  assign _zz_14 = ($signed(_zz_15) + $signed(_zz_16));
  assign _zz_15 = {_zz_6[35],_zz_6};
  assign _zz_16 = {_zz_2[35],_zz_2};
  assign _zz_17 = _zz_1[27 : 17];
  assign _zz_18 = _zz_1[26 : 17];
  assign _zz_2 = {{27'h0,1'b1},8'h0};
  assign _zz_3 = {28'hfffffff,8'h0};
  assign _zz_4 = din[35 : 0];
  assign _zz_5 = ($signed(_zz_9) + $signed(_zz_10));
  assign _zz_6 = din[35 : 0];
  always @ (*) begin
    if((_zz_11 != 9'h0))begin
      _zz_7 = ($signed(_zz_12) + $signed(_zz_13));
    end else begin
      _zz_7 = _zz_5[36 : 9];
    end
  end

  always @ (*) begin
    if(_zz_5[36])begin
      _zz_1 = _zz_7;
    end else begin
      _zz_1 = (_zz_14 >>> 9);
    end
  end

  always @ (*) begin
    if(_zz_1[27])begin
      if((! (_zz_17 == 11'h7ff)))begin
        _zz_8 = 18'h20000;
      end else begin
        _zz_8 = _zz_1[17 : 0];
      end
    end else begin
      if((_zz_18 != 10'h0))begin
        _zz_8 = 18'h1ffff;
      end else begin
        _zz_8 = _zz_1[17 : 0];
      end
    end
  end

  assign dout = _zz_8;

endmodule

//SInt36fixTo35_0_ROUNDTOINF replaced by SInt36fixTo35_0_ROUNDTOINF

module SInt36fixTo35_0_ROUNDTOINF (
  input      [35:0]   din,
  output     [35:0]   dout
);

  assign dout = din;

endmodule
