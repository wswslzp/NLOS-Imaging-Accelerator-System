//[info] running main -n 4 -hw complex fixedpoint 8 8 dft
module product(input clk,
  input reset,
  input next,
  input [31:0] i0,
  input [31:0] i1,
  input [31:0] i2,
  input [31:0] i3,
  input [31:0] i4,
  input [31:0] i5,
  input [31:0] i6,
  input [31:0] i7,
  input [31:0] i8,
  input [31:0] i9,
  input [31:0] i10,
  input [31:0] i11,
  input [31:0] i12,
  input [31:0] i13,
  input [31:0] i14,
  input [31:0] i15,
  output next_out,
  output [31:0] o0,
  output [31:0] o1,
  output [31:0] o2,
  output [31:0] o3,
  output [31:0] o4,
  output [31:0] o5,
  output [31:0] o6,
  output [31:0] o7,
  output [31:0] o8,
  output [31:0] o9,
  output [31:0] o10,
  output [31:0] o11,
  output [31:0] o12,
  output [31:0] o13,
  output [31:0] o14,
  output [31:0] o15);

  wire [31:0] s1;
  wire [31:0] s2;
  wire [31:0] s3;
  wire [31:0] s4;
  wire [31:0] s5;
  wire [31:0] s6;
  wire [31:0] s7;
  wire [31:0] s8;
  wire [31:0] s9;
  wire [31:0] s10;
  wire [31:0] s11;
  wire [31:0] s12;
  wire [31:0] s13;
  wire [31:0] s14;
  wire [31:0] s15;
  wire [31:0] s16;
  reg [15:0] s17;
  reg [15:0] s18;
  reg [15:0] s19;
  reg [15:0] s20;
  reg [15:0] s21;
  reg [15:0] s22;
  reg [15:0] s23;
  reg [15:0] s24;
  reg [15:0] s25;
  reg [15:0] s26;
  reg [15:0] s27;
  reg [15:0] s28;
  reg [15:0] s29;
  reg [15:0] s30;
  reg [15:0] s31;
  reg [15:0] s32;
  reg [15:0] s33;
  reg [15:0] s34;
  reg [15:0] s35;
  reg [15:0] s36;
  reg [15:0] s37;
  reg [15:0] s38;
  reg [15:0] s39;
  reg [15:0] s40;
  reg [15:0] s41;
  reg [15:0] s42;
  reg [15:0] s43;
  reg [15:0] s44;
  reg [15:0] s45;
  reg [15:0] s46;
  reg [15:0] s47;
  wire [15:0] s48;
  wire [15:0] s49;
  wire [15:0] s50;
  wire [15:0] s51;
  wire [15:0] s52;
  wire [15:0] s53;
  wire [15:0] s54;
  wire [15:0] s55;
  wire [15:0] s56;
  wire [15:0] s57;
  wire [15:0] s58;
  wire [15:0] s59;
  wire [15:0] s60;
  wire [15:0] s61;
  wire [15:0] s62;
  wire [15:0] s63;
  wire [15:0] s64;
  wire [15:0] s65;
  wire [15:0] s66;
  wire [15:0] s67;
  wire [15:0] s68;
  wire [15:0] s69;
  wire [15:0] s70;
  wire [15:0] s71;
  wire [15:0] s72;
  wire [15:0] s73;
  wire [15:0] s74;
  wire [15:0] s75;
  wire [15:0] s76;
  wire [15:0] s77;
  wire [15:0] s78;
  reg [15:0] s79;
  reg [15:0] s80;
  reg [15:0] s81;
  reg [15:0] s82;
  reg [15:0] s83;
  reg [15:0] s84;
  reg [15:0] s85;
  reg [15:0] s86;
  reg [15:0] s87;
  reg [15:0] s88;
  reg [15:0] s89;
  reg [15:0] s90;
  reg [15:0] s91;
  reg [15:0] s92;
  reg [15:0] s93;
  reg [15:0] s94;
  reg [15:0] s95;
  reg [15:0] s96;
  reg [15:0] s97;
  reg [15:0] s98;
  reg [15:0] s99;
  reg [15:0] s100;
  reg [15:0] s101;
  reg [15:0] s102;
  reg [15:0] s103;
  reg [15:0] s104;
  reg [15:0] s105;
  reg [15:0] s106;
  reg [15:0] s107;
  reg [15:0] s108;
  reg [15:0] s109;
  wire [15:0] s110;
  wire [15:0] s111;
  wire [15:0] s112;
  wire [15:0] s113;
  wire [15:0] s114;
  wire [15:0] s115;
  wire [15:0] s116;
  wire [15:0] s117;
  wire [15:0] s118;
  wire [15:0] s119;
  wire [15:0] s120;
  wire [15:0] s121;
  wire [15:0] s122;
  wire [15:0] s123;
  wire [15:0] s124;
  wire [15:0] s125;
  wire [15:0] s126;
  wire [15:0] s127;
  reg [15:0] s128;
  reg [15:0] s129;
  wire [15:0] s130;
  wire [15:0] s131;
  wire [15:0] s132;
  wire [15:0] s133;
  wire [15:0] s134;
  wire [15:0] s135;
  wire [15:0] s136;
  wire [15:0] s137;
  wire [15:0] s138;
  wire [15:0] s139;
  wire [15:0] s140;
  reg [15:0] s141;
  reg [15:0] s142;
  reg [15:0] s143;
  reg [15:0] s144;
  reg [15:0] s145;
  reg [15:0] s146;
  reg [15:0] s147;
  reg [15:0] s148;
  reg [15:0] s149;
  reg [15:0] s150;
  reg [15:0] s151;
  reg [15:0] s152;
  reg [15:0] s153;
  reg [15:0] s154;
  reg [15:0] s155;
  reg [15:0] s156;
  reg [15:0] s157;
  reg [15:0] s158;
  reg [15:0] s159;
  reg [15:0] s160;
  reg [15:0] s161;
  reg [15:0] s162;
  reg [15:0] s163;
  reg [15:0] s164;
  reg [15:0] s165;
  reg [15:0] s166;
  reg [15:0] s167;
  reg [15:0] s168;
  reg [15:0] s169;
  wire [15:0] s170;
  wire [15:0] s171;
  reg [15:0] s172;
  reg [15:0] s173;
  reg [15:0] s174;
  reg [15:0] s175;
  reg [15:0] s176;
  reg [15:0] s177;
  reg [15:0] s178;
  reg [15:0] s179;
  reg [15:0] s180;
  wire [15:0] s181;
  wire [15:0] s182;
  wire [15:0] s183;
  wire [15:0] s184;
  wire [15:0] s185;
  wire [15:0] s186;
  wire [15:0] s187;
  wire [15:0] s188;
  reg [15:0] s189;
  reg [15:0] s190;
  wire [15:0] s191;
  wire [15:0] s192;
  reg [15:0] s193;
  reg [15:0] s194;
  wire [15:0] s195;
  wire [15:0] s196;
  reg [15:0] s197;
  reg [15:0] s198;
  reg [15:0] s199;
  reg [15:0] s200;
  reg [15:0] s201;
  reg [15:0] s202;
  wire [15:0] s203;
  wire [15:0] s204;
  reg [15:0] s205;
  reg [15:0] s206;
  wire [15:0] s207;
  reg [15:0] s208;
  reg [15:0] s209;
  reg [15:0] s210;
  reg [15:0] s211;
  reg [15:0] s212;
  reg [15:0] s213;
  reg [15:0] s214;
  reg [15:0] s215;
  reg [15:0] s216;
  reg [15:0] s217;
  reg [15:0] s218;
  reg [15:0] s219;
  reg [15:0] s220;
  reg [15:0] s221;
  reg [15:0] s222;
  reg [15:0] s223;
  reg [15:0] s224;
  reg [15:0] s225;
  reg [15:0] s226;
  reg [15:0] s227;
  reg [15:0] s228;
  reg [15:0] s229;
  reg [15:0] s230;
  reg [15:0] s231;
  reg [15:0] s232;
  reg [15:0] s233;
  reg [15:0] s234;
  reg [15:0] s235;
  reg [15:0] s236;
  reg [15:0] s237;
  reg [15:0] s238;
  reg [15:0] s239;
  reg [15:0] s240;
  reg [15:0] s241;
  reg [15:0] s242;
  reg [15:0] s243;
  reg [15:0] s244;
  reg [15:0] s245;
  reg [15:0] s246;
  wire [15:0] s247;
  wire [15:0] s248;
  reg [15:0] s249;
  reg [15:0] s250;
  reg [15:0] s251;
  reg [15:0] s252;
  reg [15:0] s253;
  reg [15:0] s254;
  reg [15:0] s255;
  wire [15:0] s256;
  wire [15:0] s257;
  reg [15:0] s258;
  reg [15:0] s259;
  reg [15:0] s260;
  reg [15:0] s261;
  reg [15:0] s262;
  reg [15:0] s263;
  reg [15:0] s264;
  reg [15:0] s265;
  reg [15:0] s266;
  wire [15:0] s267;
  wire [15:0] s268;
  wire [15:0] s269;
  wire [15:0] s270;
  reg [15:0] s271;
  reg [15:0] s272;
  wire [15:0] s273;
  wire [15:0] s274;
  reg [15:0] s275;
  reg [15:0] s276;
  reg [15:0] s277;
  reg [15:0] s278;
  wire [15:0] s279;
  wire [15:0] s280;
  reg [15:0] s281;
  reg [15:0] s282;
  wire [15:0] s283;
  wire [15:0] s284;
  wire [15:0] s285;
  wire [15:0] s286;
  reg [15:0] s287;
  reg [15:0] s288;
  wire [15:0] s289;
  wire [15:0] s290;
  wire [15:0] s291;
  wire [15:0] s292;
  wire [15:0] s293;
  wire [15:0] s294;
  wire [15:0] s295;
  wire [15:0] s296;
  reg [15:0] s297;
  wire [15:0] s298;
  wire [15:0] s299;
  wire [15:0] s300;
  wire [15:0] s301;
  reg [15:0] s302;
  reg [15:0] s303;
  reg [15:0] s304;
  reg [15:0] s305;
  wire [15:0] s306;
  wire [15:0] s307;
  wire [15:0] s308;
  wire [15:0] s309;
  wire [15:0] s310;
  wire [15:0] s311;
  wire [15:0] s312;
  wire [15:0] s313;
  wire [15:0] s314;
  wire [15:0] s315;
  wire [15:0] s316;
  wire [15:0] s317;
  wire [15:0] s318;
  reg [15:0] s319;
  reg [15:0] s320;
  wire [15:0] s321;
  wire [15:0] s322;
  reg [15:0] s323;
  reg [15:0] s324;
  reg [15:0] s325;
  reg [15:0] s326;
  wire [15:0] s327;
  wire [15:0] s328;
  reg [15:0] s329;
  reg [15:0] s330;
  reg [15:0] s331;
  reg [15:0] s332;
  reg [15:0] s333;
  reg [15:0] s334;
  wire [31:0] s335;
  wire [31:0] s336;
  reg [31:0] s337;
  reg [31:0] s338;
  reg [15:0] s339;
  reg [15:0] s340;
  wire [31:0] s341;
  wire [31:0] s342;
  wire [31:0] s343;
  wire [31:0] s344;
  reg [31:0] s345;
  reg [31:0] s346;
  wire [31:0] s347;
  wire [31:0] s348;
  reg [15:0] s349;
  wire [31:0] s350;
  wire [31:0] s351;
  wire [31:0] s352;
  wire [31:0] s353;
  reg [15:0] s354;
  reg [15:0] s355;
  reg [15:0] s356;
  reg [15:0] s357;
  wire [31:0] s358;
  wire [31:0] s359;
  wire [31:0] s360;
  wire [31:0] s361;
  wire [31:0] s362;
  wire [31:0] s363;
  wire [31:0] s364;
  wire [31:0] s365;
  wire [31:0] s366;
  reg [15:0] s367;
  reg [15:0] s368;
  reg [31:0] s369;
  reg [31:0] s370;
  reg [15:0] s371;
  reg [15:0] s372;
  reg [15:0] s373;
  reg [15:0] s374;
  reg [31:0] s375;
  reg [31:0] s376;
  reg [15:0] s377;
  reg [15:0] s378;
  reg [15:0] s379;
  reg [15:0] s380;
  wire [15:0] s381;
  wire [15:0] s382;
  reg [15:0] s383;
  reg [15:0] s384;
  reg [31:0] s385;
  reg [31:0] s386;
  wire [15:0] s387;
  wire [15:0] s388;
  reg [15:0] s389;
  reg [15:0] s390;
  reg [31:0] s391;
  reg [31:0] s392;
  wire [15:0] s393;
  reg [15:0] s394;
  reg [15:0] s395;
  reg [15:0] s396;
  reg [15:0] s397;
  reg [15:0] s398;
  reg [15:0] s399;
  reg [15:0] s400;
  reg [15:0] s401;
  reg [15:0] s402;
  reg [15:0] s403;
  reg [15:0] s404;
  reg [15:0] s405;
  reg [15:0] s406;
  reg [31:0] s407;
  reg [31:0] s408;
  reg [15:0] s409;
  reg [15:0] s410;
  reg [15:0] s411;
  reg [15:0] s412;
  reg [31:0] s413;
  reg [31:0] s414;
  wire [15:0] s415;
  wire [15:0] s416;
  reg [15:0] s417;
  reg [15:0] s418;
  wire [31:0] s419;
  wire [31:0] s420;
  wire [15:0] s421;
  wire [15:0] s422;
  reg [31:0] s423;
  reg [31:0] s424;
  wire [31:0] s425;
  wire [31:0] s426;
  wire [15:0] s427;
  wire [15:0] s428;
  reg [31:0] s429;
  reg [31:0] s430;
  wire [31:0] s431;
  wire [15:0] s432;
  wire [15:0] s433;
  wire [15:0] s434;
  wire [15:0] s435;
  reg [15:0] s436;
  reg [15:0] s437;
  wire [15:0] s438;
  wire [15:0] s439;
  wire [15:0] s440;
  wire [15:0] s441;
  wire [15:0] s442;
  reg [15:0] s443;
  reg [15:0] s444;
  reg [31:0] s445;
  reg [31:0] s446;
  wire [15:0] s447;
  wire [15:0] s448;
  reg [15:0] s449;
  reg [15:0] s450;
  reg [31:0] s451;
  reg [31:0] s452;
  wire [15:0] s453;
  wire [15:0] s454;
  reg [15:0] s455;
  reg [15:0] s456;
  wire [15:0] s457;
  wire [15:0] s458;
  reg [15:0] s459;
  reg [15:0] s460;
  reg [15:0] s461;
  reg [15:0] s462;
  reg [15:0] s463;
  reg [15:0] s464;
  reg [31:0] s465;
  reg [31:0] s466;
  reg [15:0] s467;
  reg [15:0] s468;
  reg [31:0] s469;
  reg [31:0] s470;
  reg [15:0] s471;
  reg [15:0] s472;
  reg [15:0] s473;
  reg [15:0] s474;
  reg [31:0] s475;
  reg [31:0] s476;
  wire [15:0] s477;
  wire [15:0] s478;
  wire [15:0] s479;
  wire [15:0] s480;
  reg [31:0] s481;
  reg [31:0] s482;
  wire [15:0] s483;
  wire [15:0] s484;
  wire [15:0] s485;
  wire [15:0] s486;
  reg [15:0] s487;
  reg [15:0] s488;
  reg [31:0] s489;
  reg [31:0] s490;
  reg [31:0] s491;
  reg [31:0] s492;
  wire [15:0] s493;
  wire [15:0] s494;
  reg [15:0] s495;
  reg [15:0] s496;
  reg [15:0] s497;
  reg [15:0] s498;
  wire [15:0] s499;
  wire [15:0] s500;
  wire [15:0] s501;
  wire [15:0] s502;
  wire [15:0] s503;
  wire [15:0] s504;
  reg [31:0] s505;
  reg [31:0] s506;
  wire [15:0] s507;
  wire [15:0] s508;
  reg [31:0] s509;
  reg [31:0] s510;
  wire [15:0] s511;
  wire [15:0] s512;
  wire [15:0] s513;
  wire [15:0] s514;
  reg [31:0] s515;
  reg [31:0] s516;
  reg [31:0] s517;
  reg [31:0] s518;
  reg [31:0] s519;
  reg [31:0] s520;
  reg [31:0] s521;
  reg [31:0] s522;
  reg [15:0] s523;
  reg [15:0] s524;
  reg [31:0] s525;
  reg [31:0] s526;
  reg [15:0] s527;
  reg [15:0] s528;
  reg [15:0] s529;
  reg [15:0] s530;
  reg [15:0] s531;
  reg [15:0] s532;
  reg [15:0] s533;
  reg [15:0] s534;
  reg [15:0] s535;
  reg [15:0] s536;
  reg [15:0] s537;
  reg [15:0] s538;
  reg [31:0] s539;
  reg [31:0] s540;
  reg [31:0] s541;
  reg [31:0] s542;
  reg [15:0] s543;
  reg [31:0] s544;
  reg [31:0] s545;
  reg [31:0] s546;
  reg [31:0] s547;
  reg [31:0] s548;
  reg [31:0] s549;
  reg [31:0] s550;
  reg [31:0] s551;
  reg [15:0] s552;
  reg [15:0] s553;
  reg [31:0] s554;
  reg [31:0] s555;
  reg [15:0] s556;
  reg [15:0] s557;
  reg [15:0] s558;
  reg [15:0] s559;
  wire [15:0] s560;
  wire [15:0] s561;
  reg [15:0] s562;
  reg [15:0] s563;
  wire [15:0] s564;
  wire [15:0] s565;
  reg [15:0] s566;
  reg [15:0] s567;
  reg [31:0] s568;
  reg [31:0] s569;
  reg [31:0] s570;
  reg [31:0] s571;
  reg [15:0] s572;
  reg [31:0] s573;
  reg [31:0] s574;
  reg [31:0] s575;
  reg [31:0] s576;
  reg [31:0] s577;
  reg [31:0] s578;
  reg [31:0] s579;
  reg [31:0] s580;
  reg [15:0] s581;
  reg [15:0] s582;
  reg [31:0] s583;
  reg [31:0] s584;
  wire [15:0] s585;
  wire [15:0] s586;
  reg [15:0] s587;
  reg [15:0] s588;
  reg [15:0] s589;
  reg [15:0] s590;
  reg [15:0] s591;
  reg [15:0] s592;
  reg [31:0] s593;
  reg [31:0] s594;
  reg [31:0] s595;
  reg [31:0] s596;
  reg [15:0] s597;
  reg [31:0] s598;
  reg [31:0] s599;
  reg [31:0] s600;
  reg [31:0] s601;
  reg [31:0] s602;
  reg [31:0] s603;
  reg [31:0] s604;
  reg [31:0] s605;
  wire [15:0] s606;
  wire [15:0] s607;
  reg [31:0] s608;
  reg [31:0] s609;
  reg [31:0] s610;
  reg [31:0] s611;
  wire [15:0] s612;
  wire [15:0] s613;
  wire [15:0] s614;
  wire [15:0] s615;
  wire [15:0] s616;
  wire [15:0] s617;
  wire [15:0] s618;
  wire [31:0] s619;
  wire [31:0] s620;
  wire [31:0] s621;
  wire [31:0] s622;
  wire [31:0] s623;
  reg [15:0] s624;
  reg [15:0] s625;
  reg [15:0] s626;
  wire [15:0] s627;
  wire [15:0] s628;
  wire [15:0] s629;
  reg [15:0] s630;
  reg [15:0] s631;
  wire [15:0] s632;
  wire [15:0] s633;
  assign next_out = next;
  assign o0 = s1;
  assign o1 = s2;
  assign o2 = s3;
  assign o3 = s4;
  assign o4 = s5;
  assign o5 = s6;
  assign o6 = s7;
  assign o7 = s8;
  assign o8 = s9;
  assign o9 = s10;
  assign o10 = s11;
  assign o11 = s12;
  assign o12 = s13;
  assign o13 = s14;
  assign o14 = s15;
  assign o15 = s16;
  // Cpx(FixPlus(FixPlus(FixPlus(S20, S28), FixPlus(S36, S44)), FixPlus(FixPlus(S52, S60), FixPlus(S68, S76))), FixPlus(FixPlus(FixPlus(S21, S29), FixPlus(S37, S45)), FixPlus(FixPlus(S53, S61), FixPlus(S69, S77))))
  assign s1 = {s17, s18};
  // Cpx(FixPlus(FixPlus(FixMinus(S16, S17), FixMinus(S111, S112)), FixMinus(FixTimes(S149, S159), FixTimes(S150, S160))), FixPlus(FixPlus(FixMinus(S23, S30), FixPlus(S113, S114)), FixPlus(FixTimes(S149, S160), FixTimes(S150, S159))))
  assign s2 = {s19, s20};
  // Cpx(FixPlus(FixMinus(FixPlus(S16, S17), FixPlus(S24, S25)), FixMinus(FixTimes(S99, S109), FixTimes(S153, S110))), FixPlus(FixMinus(FixMinus(S21, S29), FixMinus(S36, S44)), FixPlus(FixTimes(S99, S110), FixTimes(S153, S109))))
  assign s3 = {s21, s22};
  // Cpx(FixPlus(FixPlus(FixMinus(S16, S17), FixMinus(S113, S118)), FixMinus(FixTimes(S155, S173), FixTimes(S156, S174))), FixPlus(FixPlus(FixPlus(S23, S30), FixPlus(S113, S118)), FixPlus(FixTimes(S155, S174), FixTimes(S156, S173))))
  assign s4 = {s23, s24};
  // Cpx(FixMinus(FixPlus(FixPlus(S16, S17), FixPlus(S24, S25)), FixPlus(FixPlus(S32, S33), FixPlus(S40, S41))), FixMinus(FixMinus(FixPlus(S21, S29), FixPlus(S37, S45)), FixMinus(FixPlus(S52, S60), FixPlus(S68, S76))))
  assign s5 = {s25, s26};
  // Cpx(FixPlus(FixMinus(FixMinus(S16, S17), FixMinus(S111, S112)), FixMinus(FixTimes(S151, S160), FixTimes(S152, S174))), FixPlus(FixMinus(FixMinus(S23, S30), FixPlus(S113, S114)), FixPlus(FixTimes(S151, S174), FixTimes(S152, S160))))
  assign s6 = {s27, s28};
  // Cpx(FixPlus(FixMinus(FixPlus(S16, S17), FixPlus(S24, S25)), FixMinus(FixTimes(S99, S110), FixTimes(S154, S110))), FixPlus(FixPlus(FixMinus(S21, S29), FixMinus(S36, S44)), FixPlus(FixTimes(S99, S110), FixTimes(S154, S110))))
  assign s7 = {s29, s30};
  // Cpx(FixPlus(FixMinus(FixMinus(S16, S17), FixMinus(S113, S118)), FixMinus(FixTimes(S157, S174), FixTimes(S158, S160))), FixPlus(FixMinus(FixPlus(S23, S30), FixPlus(S113, S118)), FixPlus(FixTimes(S157, S160), FixTimes(S158, S174))))
  assign s8 = {s31, s32};
  // Cpx(FixMinus(FixPlus(FixPlus(S20, S28), FixPlus(S36, S44)), FixPlus(FixPlus(S52, S60), FixPlus(S68, S76))), FixMinus(FixPlus(FixPlus(S21, S29), FixPlus(S37, S45)), FixPlus(FixPlus(S53, S61), FixPlus(S69, S77))))
  assign s9 = {s33, s34};
  // Cpx(FixMinus(FixPlus(FixMinus(S16, S17), FixMinus(S111, S112)), FixMinus(FixTimes(S149, S159), FixTimes(S150, S160))), FixMinus(FixPlus(FixMinus(S23, S30), FixPlus(S113, S114)), FixPlus(FixTimes(S149, S160), FixTimes(S150, S159))))
  assign s10 = {s35, s36};
  // Cpx(FixMinus(FixMinus(FixPlus(S16, S17), FixPlus(S24, S25)), FixMinus(FixTimes(S99, S109), FixTimes(S153, S110))), FixMinus(FixMinus(FixMinus(S21, S29), FixMinus(S36, S44)), FixPlus(FixTimes(S99, S110), FixTimes(S153, S109))))
  assign s11 = {s37, s38};
  // Cpx(FixMinus(FixPlus(FixMinus(S16, S17), FixMinus(S113, S118)), FixMinus(FixTimes(S155, S173), FixTimes(S156, S174))), FixMinus(FixPlus(FixPlus(S23, S30), FixPlus(S113, S118)), FixPlus(FixTimes(S155, S174), FixTimes(S156, S173))))
  assign s12 = {s39, s40};
  // Cpx(FixMinus(FixPlus(FixPlus(S16, S17), FixPlus(S24, S25)), FixPlus(FixPlus(S32, S33), FixPlus(S40, S41))), FixPlus(FixMinus(FixPlus(S21, S29), FixPlus(S37, S45)), FixMinus(FixPlus(S52, S60), FixPlus(S68, S76))))
  assign s13 = {s41, s26};
  // Cpx(FixMinus(FixMinus(FixMinus(S16, S17), FixMinus(S111, S112)), FixMinus(FixTimes(S151, S160), FixTimes(S152, S174))), FixMinus(FixMinus(FixMinus(S23, S30), FixPlus(S113, S114)), FixPlus(FixTimes(S151, S174), FixTimes(S152, S160))))
  assign s14 = {s42, s43};
  // Cpx(FixMinus(FixMinus(FixPlus(S16, S17), FixPlus(S24, S25)), FixMinus(FixTimes(S99, S110), FixTimes(S154, S110))), FixMinus(FixPlus(FixMinus(S21, S29), FixMinus(S36, S44)), FixPlus(FixTimes(S99, S110), FixTimes(S154, S110))))
  assign s15 = {s44, s45};
  // Cpx(FixMinus(FixMinus(FixMinus(S16, S17), FixMinus(S113, S118)), FixMinus(FixTimes(S157, S174), FixTimes(S158, S160))), FixMinus(FixMinus(FixPlus(S23, S30), FixPlus(S113, S118)), FixPlus(FixTimes(S157, S160), FixTimes(S158, S174))))
  assign s16 = {s46, s47};
  // FixPlus(FixPlus(FixPlus(FixPlus(S18, S19), FixPlus(S26, S27)), FixPlus(FixPlus(S34, S35), FixPlus(S42, S43))), FixPlus(FixPlus(FixPlus(S50, S51), FixPlus(S58, S59)), FixPlus(FixPlus(S66, S67), FixPlus(S74, S75))))
  assign s48 = s79 + s80;
  // FixPlus(FixPlus(FixPlus(FixPlus(S16, S17), FixPlus(S24, S25)), FixPlus(FixPlus(S32, S33), FixPlus(S40, S41))), FixPlus(FixPlus(FixPlus(S48, S49), FixPlus(S56, S57)), FixPlus(FixPlus(S64, S65), FixPlus(S72, S73))))
  assign s49 = s81 + s82;
  // FixPlus(FixPlus(FixMinus(FixMinus(S18, S19), FixMinus(S24, S25)), FixPlus(FixTimes(S38, S110), FixTimes(S95, S109))), FixPlus(FixTimes(FixPlus(S54, S125), -0.3826834323650898), FixTimes(FixPlus(S101, S126), 0.9238795325112867)))
  assign s50 = s83 + s84;
  // FixPlus(FixPlus(FixMinus(Re(S0), Re(S8)), FixMinus(FixTimes(S38, S109), FixTimes(S95, S110))), FixMinus(FixTimes(FixPlus(S54, S125), 0.9238795325112867), FixTimes(FixPlus(S101, S126), -0.3826834323650898)))
  assign s51 = s85 + s86;
  // FixPlus(FixMinus(FixMinus(FixPlus(S18, S19), FixPlus(S26, S27)), FixMinus(FixPlus(S32, S33), FixPlus(S40, S41))), FixPlus(FixTimes(FixMinus(S52, S60), -0.7071067811865475), FixTimes(FixMinus(S100, S105), 0.7071067811865476)))
  assign s52 = s87 + s88;
  // FixPlus(FixMinus(FixPlus(Re(S0), Re(S8)), FixPlus(Re(S4), Re(S12))), FixMinus(FixTimes(FixMinus(S52, S60), 0.7071067811865476), FixTimes(FixMinus(S100, S105), -0.7071067811865475)))
  assign s53 = s89 + s90;
  // FixPlus(FixPlus(FixPlus(FixMinus(S18, S19), FixMinus(S24, S25)), FixPlus(FixTimes(S38, S110), FixTimes(S96, S110))), FixPlus(FixTimes(FixPlus(S54, S129), -0.9238795325112867), FixTimes(FixPlus(S102, S130), 0.38268343236508984)))
  assign s54 = s91 + s92;
  // FixPlus(FixPlus(FixMinus(Re(S0), Re(S8)), FixMinus(FixTimes(S38, S110), FixTimes(S96, S110))), FixMinus(FixTimes(FixPlus(S54, S129), 0.38268343236508984), FixTimes(FixPlus(S102, S130), -0.9238795325112867)))
  assign s55 = s93 + s94;
  // FixMinus(FixMinus(FixPlus(FixPlus(S18, S19), FixPlus(S26, S27)), FixPlus(FixPlus(S34, S35), FixPlus(S42, S43))), FixMinus(FixPlus(FixPlus(S48, S49), FixPlus(S56, S57)), FixPlus(FixPlus(S64, S65), FixPlus(S72, S73))))
  assign s56 = s95 - s96;
  // FixMinus(FixPlus(FixPlus(Re(S0), Re(S8)), FixPlus(Re(S4), Re(S12))), FixPlus(FixPlus(Re(S2), Re(S10)), FixPlus(Re(S6), Re(S14))))
  assign s57 = s97 - s98;
  // FixPlus(FixMinus(FixMinus(FixMinus(S18, S19), FixMinus(S24, S25)), FixPlus(FixTimes(S38, S110), FixTimes(S95, S109))), FixPlus(FixTimes(FixMinus(S54, S125), -0.9238795325112867), FixTimes(FixMinus(S101, S126), -0.3826834323650898)))
  assign s58 = s99 + s100;
  // FixPlus(FixMinus(FixMinus(Re(S0), Re(S8)), FixMinus(FixTimes(S38, S109), FixTimes(S95, S110))), FixMinus(FixTimes(FixMinus(S54, S125), -0.3826834323650898), FixTimes(FixMinus(S101, S126), -0.9238795325112867)))
  assign s59 = s101 + s102;
  // FixPlus(FixPlus(FixMinus(FixPlus(S18, S19), FixPlus(S26, S27)), FixMinus(FixPlus(S32, S33), FixPlus(S40, S41))), FixPlus(FixTimes(FixMinus(S52, S60), -0.7071067811865475), FixTimes(FixPlus(S100, S105), -0.7071067811865475)))
  assign s60 = s103 + s104;
  // FixPlus(FixMinus(FixPlus(Re(S0), Re(S8)), FixPlus(Re(S4), Re(S12))), FixMinus(FixTimes(FixMinus(S52, S60), -0.7071067811865475), FixTimes(FixPlus(S100, S105), -0.7071067811865475)))
  assign s61 = s89 + s105;
  // FixPlus(FixMinus(FixPlus(FixMinus(S18, S19), FixMinus(S24, S25)), FixPlus(FixTimes(S38, S110), FixTimes(S96, S110))), FixPlus(FixTimes(FixMinus(S54, S129), -0.3826834323650898), FixTimes(FixMinus(S102, S130), -0.9238795325112867)))
  assign s62 = s106 + s107;
  // FixPlus(FixMinus(FixMinus(Re(S0), Re(S8)), FixMinus(FixTimes(S38, S110), FixTimes(S96, S110))), FixMinus(FixTimes(FixMinus(S54, S129), -0.9238795325112867), FixTimes(FixMinus(S102, S130), -0.3826834323650898)))
  assign s63 = s108 + s109;
  // FixMinus(FixPlus(FixPlus(FixPlus(S18, S19), FixPlus(S26, S27)), FixPlus(FixPlus(S34, S35), FixPlus(S42, S43))), FixPlus(FixPlus(FixPlus(S50, S51), FixPlus(S58, S59)), FixPlus(FixPlus(S66, S67), FixPlus(S74, S75))))
  assign s64 = s79 - s80;
  // FixMinus(FixPlus(FixPlus(FixPlus(S16, S17), FixPlus(S24, S25)), FixPlus(FixPlus(S32, S33), FixPlus(S40, S41))), FixPlus(FixPlus(FixPlus(S48, S49), FixPlus(S56, S57)), FixPlus(FixPlus(S64, S65), FixPlus(S72, S73))))
  assign s65 = s81 - s82;
  // FixMinus(FixPlus(FixMinus(FixMinus(S18, S19), FixMinus(S24, S25)), FixPlus(FixTimes(S38, S110), FixTimes(S95, S109))), FixPlus(FixTimes(FixPlus(S54, S125), -0.3826834323650898), FixTimes(FixPlus(S101, S126), 0.9238795325112867)))
  assign s66 = s83 - s84;
  // FixMinus(FixPlus(FixMinus(Re(S0), Re(S8)), FixMinus(FixTimes(S38, S109), FixTimes(S95, S110))), FixMinus(FixTimes(FixPlus(S54, S125), 0.9238795325112867), FixTimes(FixPlus(S101, S126), -0.3826834323650898)))
  assign s67 = s85 - s86;
  // FixMinus(FixMinus(FixMinus(FixPlus(S18, S19), FixPlus(S26, S27)), FixMinus(FixPlus(S32, S33), FixPlus(S40, S41))), FixPlus(FixTimes(FixMinus(S52, S60), -0.7071067811865475), FixTimes(FixMinus(S100, S105), 0.7071067811865476)))
  assign s68 = s87 - s88;
  // FixMinus(FixMinus(FixPlus(Re(S0), Re(S8)), FixPlus(Re(S4), Re(S12))), FixMinus(FixTimes(FixMinus(S52, S60), 0.7071067811865476), FixTimes(FixMinus(S100, S105), -0.7071067811865475)))
  assign s69 = s89 - s90;
  // FixMinus(FixPlus(FixPlus(FixMinus(S18, S19), FixMinus(S24, S25)), FixPlus(FixTimes(S38, S110), FixTimes(S96, S110))), FixPlus(FixTimes(FixPlus(S54, S129), -0.9238795325112867), FixTimes(FixPlus(S102, S130), 0.38268343236508984)))
  assign s70 = s91 - s92;
  // FixMinus(FixPlus(FixMinus(Re(S0), Re(S8)), FixMinus(FixTimes(S38, S110), FixTimes(S96, S110))), FixMinus(FixTimes(FixPlus(S54, S129), 0.38268343236508984), FixTimes(FixPlus(S102, S130), -0.9238795325112867)))
  assign s71 = s93 - s94;
  // FixPlus(FixMinus(FixPlus(FixPlus(S18, S19), FixPlus(S26, S27)), FixPlus(FixPlus(S34, S35), FixPlus(S42, S43))), FixMinus(FixPlus(FixPlus(S48, S49), FixPlus(S56, S57)), FixPlus(FixPlus(S64, S65), FixPlus(S72, S73))))
  assign s72 = s95 + s96;
  // FixMinus(FixMinus(FixMinus(FixMinus(S18, S19), FixMinus(S24, S25)), FixPlus(FixTimes(S38, S110), FixTimes(S95, S109))), FixPlus(FixTimes(FixMinus(S54, S125), -0.9238795325112867), FixTimes(FixMinus(S101, S126), -0.3826834323650898)))
  assign s73 = s99 - s100;
  // FixMinus(FixMinus(FixMinus(Re(S0), Re(S8)), FixMinus(FixTimes(S38, S109), FixTimes(S95, S110))), FixMinus(FixTimes(FixMinus(S54, S125), -0.3826834323650898), FixTimes(FixMinus(S101, S126), -0.9238795325112867)))
  assign s74 = s101 - s102;
  // FixMinus(FixPlus(FixMinus(FixPlus(S18, S19), FixPlus(S26, S27)), FixMinus(FixPlus(S32, S33), FixPlus(S40, S41))), FixPlus(FixTimes(FixMinus(S52, S60), -0.7071067811865475), FixTimes(FixPlus(S100, S105), -0.7071067811865475)))
  assign s75 = s103 - s104;
  // FixMinus(FixMinus(FixPlus(Re(S0), Re(S8)), FixPlus(Re(S4), Re(S12))), FixMinus(FixTimes(FixMinus(S52, S60), -0.7071067811865475), FixTimes(FixPlus(S100, S105), -0.7071067811865475)))
  assign s76 = s89 - s105;
  // FixMinus(FixMinus(FixPlus(FixMinus(S18, S19), FixMinus(S24, S25)), FixPlus(FixTimes(S38, S110), FixTimes(S96, S110))), FixPlus(FixTimes(FixMinus(S54, S129), -0.3826834323650898), FixTimes(FixMinus(S102, S130), -0.9238795325112867)))
  assign s77 = s106 - s107;
  // FixMinus(FixMinus(FixMinus(Re(S0), Re(S8)), FixMinus(FixTimes(S38, S110), FixTimes(S96, S110))), FixMinus(FixTimes(FixMinus(S54, S129), -0.9238795325112867), FixTimes(FixMinus(S102, S130), -0.3826834323650898)))
  assign s78 = s108 - s109;
  // FixPlus(FixPlus(FixPlus(Im(S0), Im(S8)), FixPlus(Im(S4), Im(S12))), FixPlus(FixPlus(Im(S2), Im(S10)), FixPlus(Im(S6), Im(S14))))
  assign s110 = s141 + s142;
  // FixPlus(FixPlus(FixPlus(Im(S1), Im(S9)), FixPlus(Im(S5), Im(S13))), FixPlus(FixPlus(Im(S3), Im(S11)), FixPlus(Im(S7), Im(S15))))
  assign s111 = s143 + s144;
  // FixPlus(FixPlus(FixPlus(Re(S0), Re(S8)), FixPlus(Re(S4), Re(S12))), FixPlus(FixPlus(Re(S2), Re(S10)), FixPlus(Re(S6), Re(S14))))
  assign s112 = s128 + s129;
  // FixPlus(FixPlus(FixPlus(Re(S1), Re(S9)), FixPlus(Re(S5), Re(S13))), FixPlus(FixPlus(Re(S3), Re(S11)), FixPlus(Re(S7), Re(S15))))
  assign s113 = s145 + s146;
  // FixPlus(FixMinus(FixMinus(Im(S0), Im(S8)), FixMinus(Re(S4), Re(S12))), FixPlus(FixTimes(FixMinus(S32, S33), -0.7071067811865475), FixTimes(FixMinus(S39, S46), 0.7071067811865476)))
  assign s114 = s147 + s148;
  // FixPlus(FixTimes(FixPlus(FixMinus(S48, S49), FixMinus(S121, S122)), -0.3826834323650898), FixTimes(FixPlus(FixMinus(S55, S62), FixPlus(S123, S124)), 0.9238795325112867))
  assign s115 = s149 + s150;
  // FixPlus(FixMinus(Re(Input()), Re(Input())), FixMinus(FixTimes(FixMinus(S32, S33), 0.7071067811865476), FixTimes(FixMinus(S39, S46), -0.7071067811865475)))
  assign s116 = s151 + s152;
  // FixMinus(FixTimes(FixPlus(FixMinus(S48, S49), FixMinus(S121, S122)), 0.9238795325112867), FixTimes(FixPlus(FixMinus(S55, S62), FixPlus(S123, S124)), -0.3826834323650898))
  assign s117 = s153 - s154;
  // FixMinus(FixMinus(FixPlus(Im(S0), Im(S8)), FixPlus(Im(S4), Im(S12))), FixMinus(FixPlus(Re(S2), Re(S10)), FixPlus(Re(S6), Re(S14))))
  assign s118 = s155 - s156;
  // FixPlus(FixTimes(FixMinus(FixPlus(S48, S49), FixPlus(S56, S57)), -0.7071067811865475), FixTimes(FixMinus(FixMinus(S53, S61), FixMinus(S68, S76)), 0.7071067811865476))
  assign s119 = s157 + s158;
  // FixMinus(FixPlus(Re(Input()), Re(Input())), FixPlus(Re(Input()), Re(Input())))
  assign s120 = s159 - s160;
  // FixMinus(FixTimes(FixMinus(FixPlus(S48, S49), FixPlus(S56, S57)), 0.7071067811865476), FixTimes(FixMinus(FixMinus(S53, S61), FixMinus(S68, S76)), -0.7071067811865475))
  assign s121 = s161 - s162;
  // FixPlus(FixPlus(FixMinus(Im(S0), Im(S8)), FixMinus(Re(S4), Re(S12))), FixPlus(FixTimes(FixMinus(S32, S33), -0.7071067811865475), FixTimes(FixPlus(S39, S46), -0.7071067811865475)))
  assign s122 = s163 + s164;
  // FixPlus(FixTimes(FixPlus(FixMinus(S48, S49), FixMinus(S123, S128)), -0.9238795325112867), FixTimes(FixPlus(FixPlus(S55, S62), FixPlus(S123, S128)), 0.38268343236508984))
  assign s123 = s165 + s166;
  // FixPlus(FixMinus(Re(Input()), Re(Input())), FixMinus(FixTimes(FixMinus(S32, S33), -0.7071067811865475), FixTimes(FixPlus(S39, S46), -0.7071067811865475)))
  assign s124 = s151 + s167;
  // FixMinus(FixTimes(FixPlus(FixMinus(S48, S49), FixMinus(S123, S128)), 0.38268343236508984), FixTimes(FixPlus(FixPlus(S55, S62), FixPlus(S123, S128)), -0.9238795325112867))
  assign s125 = s168 - s169;
  // FixMinus(FixPlus(FixPlus(Im(S0), Im(S8)), FixPlus(Im(S4), Im(S12))), FixPlus(FixPlus(Im(S2), Im(S10)), FixPlus(Im(S6), Im(S14))))
  assign s126 = s141 - s142;
  // FixMinus(FixPlus(FixPlus(Re(S1), Re(S9)), FixPlus(Re(S5), Re(S13))), FixPlus(FixPlus(Re(S3), Re(S11)), FixPlus(Re(S7), Re(S15))))
  assign s127 = s145 - s146;
  // FixMinus(FixMinus(FixMinus(Im(S0), Im(S8)), FixMinus(Re(S4), Re(S12))), FixPlus(FixTimes(FixMinus(S32, S33), -0.7071067811865475), FixTimes(FixMinus(S39, S46), 0.7071067811865476)))
  assign s130 = s147 - s148;
  // FixPlus(FixTimes(FixMinus(FixMinus(S48, S49), FixMinus(S121, S122)), -0.9238795325112867), FixTimes(FixMinus(FixMinus(S55, S62), FixPlus(S123, S124)), -0.3826834323650898))
  assign s131 = s172 + s173;
  // FixMinus(FixMinus(Re(Input()), Re(Input())), FixMinus(FixTimes(FixMinus(S32, S33), 0.7071067811865476), FixTimes(FixMinus(S39, S46), -0.7071067811865475)))
  assign s132 = s151 - s152;
  // FixMinus(FixTimes(FixMinus(FixMinus(S48, S49), FixMinus(S121, S122)), -0.3826834323650898), FixTimes(FixMinus(FixMinus(S55, S62), FixPlus(S123, S124)), -0.9238795325112867))
  assign s133 = s174 - s175;
  // FixPlus(FixMinus(FixPlus(Im(S0), Im(S8)), FixPlus(Im(S4), Im(S12))), FixMinus(FixPlus(Re(S2), Re(S10)), FixPlus(Re(S6), Re(S14))))
  assign s134 = s155 + s156;
  // FixPlus(FixTimes(FixMinus(FixPlus(S48, S49), FixPlus(S56, S57)), -0.7071067811865475), FixTimes(FixPlus(FixMinus(S53, S61), FixMinus(S68, S76)), -0.7071067811865475))
  assign s135 = s157 + s176;
  // FixMinus(FixTimes(FixMinus(FixPlus(S48, S49), FixPlus(S56, S57)), -0.7071067811865475), FixTimes(FixPlus(FixMinus(S53, S61), FixMinus(S68, S76)), -0.7071067811865475))
  assign s136 = s157 - s176;
  // FixMinus(FixPlus(FixMinus(Im(S0), Im(S8)), FixMinus(Re(S4), Re(S12))), FixPlus(FixTimes(FixMinus(S32, S33), -0.7071067811865475), FixTimes(FixPlus(S39, S46), -0.7071067811865475)))
  assign s137 = s163 - s164;
  // FixPlus(FixTimes(FixMinus(FixMinus(S48, S49), FixMinus(S123, S128)), -0.3826834323650898), FixTimes(FixMinus(FixPlus(S55, S62), FixPlus(S123, S128)), -0.9238795325112867))
  assign s138 = s177 + s178;
  // FixMinus(FixMinus(Re(Input()), Re(Input())), FixMinus(FixTimes(FixMinus(S32, S33), -0.7071067811865475), FixTimes(FixPlus(S39, S46), -0.7071067811865475)))
  assign s139 = s151 - s167;
  // FixMinus(FixTimes(FixMinus(FixMinus(S48, S49), FixMinus(S123, S128)), -0.9238795325112867), FixTimes(FixMinus(FixPlus(S55, S62), FixPlus(S123, S128)), -0.3826834323650898))
  assign s140 = s179 - s180;
  // FixPlus(FixPlus(Re(Input()), Re(Input())), FixPlus(Re(Input()), Re(Input())))
  assign s170 = s199 + s200;
  // FixPlus(FixPlus(Re(Input()), Re(Input())), FixPlus(Re(Input()), Re(Input())))
  assign s171 = s210 + s211;
  // FixPlus(FixPlus(Im(Input()), Im(Input())), FixPlus(Im(Input()), Im(Input())))
  assign s181 = s221 + s222;
  // FixPlus(FixPlus(Im(Input()), Im(Input())), FixPlus(Im(Input()), Im(Input())))
  assign s182 = s223 + s224;
  // FixPlus(FixPlus(Im(Input()), Im(Input())), FixPlus(Im(Input()), Im(Input())))
  assign s183 = s225 + s226;
  // FixPlus(FixPlus(Im(Input()), Im(Input())), FixPlus(Im(Input()), Im(Input())))
  assign s184 = s227 + s228;
  // FixPlus(FixPlus(Re(Input()), Re(Input())), FixPlus(Re(Input()), Re(Input())))
  assign s185 = s229 + s230;
  // FixPlus(FixPlus(Re(Input()), Re(Input())), FixPlus(Re(Input()), Re(Input())))
  assign s186 = s231 + s232;
  // FixMinus(FixMinus(Im(Input()), Im(Input())), FixMinus(Re(Input()), Re(Input())))
  assign s187 = s233 - s234;
  // FixPlus(FixTimes(FixMinus(Re(S2), Re(S10)), -0.7071067811865475), FixTimes(FixMinus(FixMinus(S34, S35), FixMinus(S40, S41)), 0.7071067811865476))
  assign s188 = s235 + s236;
  // FixMinus(Re(Input()), Re(Input()))
  assign s191 = s239 - s240;
  // FixMinus(FixTimes(FixMinus(Re(S2), Re(S10)), 0.7071067811865476), FixTimes(FixMinus(FixMinus(S34, S35), FixMinus(S40, S41)), -0.7071067811865475))
  assign s192 = s241 - s242;
  // FixMinus(FixPlus(Im(Input()), Im(Input())), FixPlus(Im(Input()), Im(Input())))
  assign s195 = s221 - s222;
  // FixMinus(FixPlus(Re(Input()), Re(Input())), FixPlus(Re(Input()), Re(Input())))
  assign s196 = s210 - s211;
  // FixPlus(FixMinus(Im(Input()), Im(Input())), FixMinus(Re(Input()), Re(Input())))
  assign s203 = s233 + s234;
  // FixPlus(FixTimes(FixMinus(Re(S2), Re(S10)), -0.7071067811865475), FixTimes(FixPlus(FixMinus(S34, S35), FixMinus(S40, S41)), -0.7071067811865475))
  assign s204 = s235 + s251;
  // FixMinus(FixTimes(FixMinus(Re(S2), Re(S10)), -0.7071067811865475), FixTimes(FixPlus(FixMinus(S34, S35), FixMinus(S40, S41)), -0.7071067811865475))
  assign s207 = s235 - s251;
  // FixPlus(Re(Input()), Re(Input()))
  assign s247 = s285 + s286;
  // FixPlus(Re(Input()), Re(Input()))
  assign s248 = s293 + s294;
  // FixPlus(Re(Input()), Re(Input()))
  assign s256 = s302 + s303;
  // FixPlus(Re(Input()), Re(Input()))
  assign s257 = s304 + s305;
  // FixPlus(Im(Input()), Im(Input()))
  assign s267 = s315 + s316;
  // FixPlus(Im(Input()), Im(Input()))
  assign s268 = s317 + s318;
  // FixPlus(Im(Input()), Im(Input()))
  assign s269 = s319 + s320;
  // FixPlus(Im(Input()), Im(Input()))
  assign s270 = s321 + s322;
  // FixPlus(Im(Input()), Im(Input()))
  assign s273 = s325 + s326;
  // FixPlus(Im(Input()), Im(Input()))
  assign s274 = s327 + s328;
  // FixMinus(Im(Input()), Im(Input()))
  assign s279 = s315 - s316;
  // FixMinus(Re(Input()), Re(Input()))
  assign s280 = s293 - s294;
  // FixTimes(FixPlus(FixMinus(Re(S1), Re(S9)), FixMinus(FixTimes(S70, S109), FixTimes(S107, S110))), -0.3826834323650898)
  assign s283 = s335[29:14];
  // FixTimes(FixPlus(FixMinus(FixMinus(S50, S51), FixMinus(S56, S57)), FixPlus(FixTimes(S70, S110), FixTimes(S107, S109))), 0.9238795325112867)
  assign s284 = s336[29:14];
  // Re(Input())
  assign s285 = s337[15:0];
  // Re(Input())
  assign s286 = s338[15:0];
  // FixTimes(FixPlus(FixMinus(Re(S1), Re(S9)), FixMinus(FixTimes(S70, S109), FixTimes(S107, S110))), 0.9238795325112867)
  assign s289 = s341[29:14];
  // FixTimes(FixPlus(FixMinus(FixMinus(S50, S51), FixMinus(S56, S57)), FixPlus(FixTimes(S70, S110), FixTimes(S107, S109))), -0.3826834323650898)
  assign s290 = s342[29:14];
  // FixTimes(FixMinus(FixPlus(Re(S1), Re(S9)), FixPlus(Re(S5), Re(S13))), -0.7071067811865475)
  assign s291 = s343[29:14];
  // FixTimes(FixMinus(FixMinus(FixPlus(S50, S51), FixPlus(S58, S59)), FixMinus(FixPlus(S64, S65), FixPlus(S72, S73))), 0.7071067811865476)
  assign s292 = s344[29:14];
  // Re(Input())
  assign s293 = s345[15:0];
  // Re(Input())
  assign s294 = s346[15:0];
  // FixTimes(FixMinus(FixPlus(Re(S1), Re(S9)), FixPlus(Re(S5), Re(S13))), 0.7071067811865476)
  assign s295 = s347[29:14];
  // FixTimes(FixMinus(FixMinus(FixPlus(S50, S51), FixPlus(S58, S59)), FixMinus(FixPlus(S64, S65), FixPlus(S72, S73))), -0.7071067811865475)
  assign s296 = s348[29:14];
  // FixTimes(FixPlus(FixMinus(Re(S1), Re(S9)), FixMinus(FixTimes(S70, S110), FixTimes(S108, S110))), -0.9238795325112867)
  assign s298 = s350[29:14];
  // FixTimes(FixPlus(FixPlus(FixMinus(S50, S51), FixMinus(S56, S57)), FixPlus(FixTimes(S70, S110), FixTimes(S108, S110))), 0.38268343236508984)
  assign s299 = s351[29:14];
  // FixTimes(FixPlus(FixMinus(Re(S1), Re(S9)), FixMinus(FixTimes(S70, S110), FixTimes(S108, S110))), 0.38268343236508984)
  assign s300 = s352[29:14];
  // FixTimes(FixPlus(FixPlus(FixMinus(S50, S51), FixMinus(S56, S57)), FixPlus(FixTimes(S70, S110), FixTimes(S108, S110))), -0.9238795325112867)
  assign s301 = s353[29:14];
  // FixTimes(FixMinus(FixMinus(Re(S1), Re(S9)), FixMinus(FixTimes(S70, S109), FixTimes(S107, S110))), -0.9238795325112867)
  assign s306 = s358[29:14];
  // FixTimes(FixMinus(FixMinus(FixMinus(S50, S51), FixMinus(S56, S57)), FixPlus(FixTimes(S70, S110), FixTimes(S107, S109))), -0.3826834323650898)
  assign s307 = s359[29:14];
  // FixTimes(FixMinus(FixMinus(Re(S1), Re(S9)), FixMinus(FixTimes(S70, S109), FixTimes(S107, S110))), -0.3826834323650898)
  assign s308 = s360[29:14];
  // FixTimes(FixMinus(FixMinus(FixMinus(S50, S51), FixMinus(S56, S57)), FixPlus(FixTimes(S70, S110), FixTimes(S107, S109))), -0.9238795325112867)
  assign s309 = s361[29:14];
  // FixTimes(FixPlus(FixMinus(FixPlus(S50, S51), FixPlus(S58, S59)), FixMinus(FixPlus(S64, S65), FixPlus(S72, S73))), -0.7071067811865475)
  assign s310 = s362[29:14];
  // FixTimes(FixMinus(FixMinus(Re(S1), Re(S9)), FixMinus(FixTimes(S70, S110), FixTimes(S108, S110))), -0.3826834323650898)
  assign s311 = s363[29:14];
  // FixTimes(FixMinus(FixPlus(FixMinus(S50, S51), FixMinus(S56, S57)), FixPlus(FixTimes(S70, S110), FixTimes(S108, S110))), -0.9238795325112867)
  assign s312 = s364[29:14];
  // FixTimes(FixMinus(FixMinus(Re(S1), Re(S9)), FixMinus(FixTimes(S70, S110), FixTimes(S108, S110))), -0.9238795325112867)
  assign s313 = s365[29:14];
  // FixTimes(FixMinus(FixPlus(FixMinus(S50, S51), FixMinus(S56, S57)), FixPlus(FixTimes(S70, S110), FixTimes(S108, S110))), -0.3826834323650898)
  assign s314 = s366[29:14];
  // Im(Input())
  assign s315 = s337[31:16];
  // Im(Input())
  assign s316 = s338[31:16];
  // Im(Input())
  assign s317 = s345[31:16];
  // Im(Input())
  assign s318 = s346[31:16];
  // Im(Input())
  assign s321 = s369[31:16];
  // Im(Input())
  assign s322 = s370[31:16];
  // Im(Input())
  assign s327 = s375[31:16];
  // Im(Input())
  assign s328 = s376[31:16];
  assign s335 = $signed(s383) * $signed(16'd59267);
  assign s336 = $signed(s384) * $signed(16'd15136);
  assign s341 = $signed(s383) * $signed(16'd15136);
  assign s342 = $signed(s384) * $signed(16'd59267);
  assign s343 = $signed(s389) * $signed(16'd53951);
  assign s344 = $signed(s390) * $signed(16'd11585);
  assign s347 = $signed(s389) * $signed(16'd11585);
  assign s348 = $signed(s390) * $signed(16'd53951);
  assign s350 = $signed(s394) * $signed(16'd50400);
  assign s351 = $signed(s395) * $signed(16'd6269);
  assign s352 = $signed(s394) * $signed(16'd6269);
  assign s353 = $signed(s395) * $signed(16'd50400);
  assign s358 = $signed(s400) * $signed(16'd50400);
  assign s359 = $signed(s401) * $signed(16'd59267);
  assign s360 = $signed(s400) * $signed(16'd59267);
  assign s361 = $signed(s401) * $signed(16'd50400);
  assign s362 = $signed(s402) * $signed(16'd53951);
  assign s363 = $signed(s403) * $signed(16'd59267);
  assign s364 = $signed(s404) * $signed(16'd50400);
  assign s365 = $signed(s403) * $signed(16'd50400);
  assign s366 = $signed(s404) * $signed(16'd59267);
  // FixTimes(FixMinus(Re(Input()), Re(Input())), -0.7071067811865475)
  assign s381 = s419[29:14];
  // FixTimes(FixMinus(FixMinus(Im(S2), Im(S10)), FixMinus(Re(S6), Re(S14))), 0.7071067811865476)
  assign s382 = s420[29:14];
  // FixTimes(FixMinus(Re(Input()), Re(Input())), 0.7071067811865476)
  assign s387 = s425[29:14];
  // FixTimes(FixMinus(FixMinus(Im(S2), Im(S10)), FixMinus(Re(S6), Re(S14))), -0.7071067811865475)
  assign s388 = s426[29:14];
  // FixTimes(FixPlus(FixMinus(Im(S2), Im(S10)), FixMinus(Re(S6), Re(S14))), -0.7071067811865475)
  assign s393 = s431[29:14];
  // FixPlus(Re(Input()), Re(Input()))
  assign s415 = s453 + s454;
  // FixPlus(Re(Input()), Re(Input()))
  assign s416 = s455 + s456;
  assign s419 = $signed(s459) * $signed(16'd53951);
  assign s420 = $signed(s460) * $signed(16'd11585);
  // FixPlus(FixMinus(Re(Input()), Re(Input())), FixMinus(FixTimes(FixMinus(S64, S65), 0.7071067811865476), FixTimes(FixMinus(S71, S78), -0.7071067811865475)))
  assign s421 = s461 + s462;
  // FixPlus(FixMinus(FixMinus(Im(S1), Im(S9)), FixMinus(Re(S5), Re(S13))), FixPlus(FixTimes(FixMinus(S64, S65), -0.7071067811865475), FixTimes(FixMinus(S71, S78), 0.7071067811865476)))
  assign s422 = s463 + s464;
  assign s425 = $signed(s459) * $signed(16'd11585);
  assign s426 = $signed(s460) * $signed(16'd53951);
  // FixMinus(FixPlus(Re(Input()), Re(Input())), FixPlus(Re(Input()), Re(Input())))
  assign s427 = s377 - s378;
  // FixMinus(FixMinus(FixPlus(Im(S1), Im(S9)), FixPlus(Im(S5), Im(S13))), FixMinus(FixPlus(Re(S3), Re(S11)), FixPlus(Re(S7), Re(S15))))
  assign s428 = s467 - s468;
  assign s431 = $signed(s471) * $signed(16'd53951);
  // FixPlus(FixMinus(Re(Input()), Re(Input())), FixMinus(FixTimes(FixMinus(S64, S65), -0.7071067811865475), FixTimes(FixPlus(S71, S78), -0.7071067811865475)))
  assign s432 = s461 + s472;
  // FixPlus(FixPlus(FixMinus(Im(S1), Im(S9)), FixMinus(Re(S5), Re(S13))), FixPlus(FixTimes(FixMinus(S64, S65), -0.7071067811865475), FixTimes(FixPlus(S71, S78), -0.7071067811865475)))
  assign s433 = s473 + s474;
  // Re(Input())
  assign s434 = s475[15:0];
  // Re(Input())
  assign s435 = s476[15:0];
  // FixMinus(FixMinus(Re(Input()), Re(Input())), FixMinus(FixTimes(FixMinus(S64, S65), 0.7071067811865476), FixTimes(FixMinus(S71, S78), -0.7071067811865475)))
  assign s438 = s461 - s462;
  // FixMinus(FixMinus(FixMinus(Im(S1), Im(S9)), FixMinus(Re(S5), Re(S13))), FixPlus(FixTimes(FixMinus(S64, S65), -0.7071067811865475), FixTimes(FixMinus(S71, S78), 0.7071067811865476)))
  assign s439 = s463 - s464;
  // FixPlus(FixMinus(FixPlus(Im(S1), Im(S9)), FixPlus(Im(S5), Im(S13))), FixMinus(FixPlus(Re(S3), Re(S11)), FixPlus(Re(S7), Re(S15))))
  assign s440 = s467 + s468;
  // FixMinus(FixMinus(Re(Input()), Re(Input())), FixMinus(FixTimes(FixMinus(S64, S65), -0.7071067811865475), FixTimes(FixPlus(S71, S78), -0.7071067811865475)))
  assign s441 = s461 - s472;
  // FixMinus(FixPlus(FixMinus(Im(S1), Im(S9)), FixMinus(Re(S5), Re(S13))), FixPlus(FixTimes(FixMinus(S64, S65), -0.7071067811865475), FixTimes(FixPlus(S71, S78), -0.7071067811865475)))
  assign s442 = s473 - s474;
  // FixPlus(Im(Input()), Im(Input()))
  assign s447 = s483 + s484;
  // FixPlus(Im(Input()), Im(Input()))
  assign s448 = s485 + s486;
  // Re(Input())
  assign s453 = s491[15:0];
  // Re(Input())
  assign s454 = s492[15:0];
  // FixPlus(Re(Input()), Re(Input()))
  assign s457 = s495 + s496;
  // FixPlus(Re(Input()), Re(Input()))
  assign s458 = s497 + s498;
  // Re(Input())
  assign s477 = s517[15:0];
  // Re(Input())
  assign s478 = s518[15:0];
  // Im(Input())
  assign s479 = s515[31:16];
  // Im(Input())
  assign s480 = s516[31:16];
  // Im(Input())
  assign s483 = s519[31:16];
  // Im(Input())
  assign s484 = s520[31:16];
  // Im(Input())
  assign s485 = s521[31:16];
  // Im(Input())
  assign s486 = s522[31:16];
  // Re(Input())
  assign s493 = s521[15:0];
  // Re(Input())
  assign s494 = s522[15:0];
  // FixMinus(Re(Input()), Re(Input()))
  assign s499 = s434 - s435;
  // FixMinus(FixMinus(Im(Input()), Im(Input())), FixMinus(Re(Input()), Re(Input())))
  assign s500 = s531 - s532;
  // FixMinus(Re(Input()), Re(Input()))
  assign s501 = s453 - s454;
  // FixMinus(FixTimes(FixMinus(Re(S3), Re(S11)), 0.7071067811865476), FixTimes(FixMinus(FixMinus(S66, S67), FixMinus(S72, S73)), -0.7071067811865475))
  assign s502 = s533 - s534;
  // FixMinus(FixMinus(Im(Input()), Im(Input())), FixMinus(Re(Input()), Re(Input())))
  assign s503 = s535 - s536;
  // FixPlus(FixTimes(FixMinus(Re(S3), Re(S11)), -0.7071067811865475), FixTimes(FixMinus(FixMinus(S66, S67), FixMinus(S72, S73)), 0.7071067811865476))
  assign s504 = s537 + s538;
  // FixMinus(FixPlus(Im(Input()), Im(Input())), FixPlus(Im(Input()), Im(Input())))
  assign s507 = s409 - s410;
  // FixMinus(FixPlus(Re(Input()), Re(Input())), FixPlus(Re(Input()), Re(Input())))
  assign s508 = s417 - s418;
  // FixPlus(FixMinus(Im(Input()), Im(Input())), FixMinus(Re(Input()), Re(Input())))
  assign s511 = s531 + s532;
  // FixMinus(FixTimes(FixMinus(Re(S3), Re(S11)), -0.7071067811865475), FixTimes(FixPlus(FixMinus(S66, S67), FixMinus(S72, S73)), -0.7071067811865475))
  assign s512 = s537 - s543;
  // FixPlus(FixMinus(Im(Input()), Im(Input())), FixMinus(Re(Input()), Re(Input())))
  assign s513 = s535 + s536;
  // FixPlus(FixTimes(FixMinus(Re(S3), Re(S11)), -0.7071067811865475), FixTimes(FixPlus(FixMinus(S66, S67), FixMinus(S72, S73)), -0.7071067811865475))
  assign s514 = s537 + s543;
  // FixMinus(Im(Input()), Im(Input()))
  assign s560 = s479 - s480;
  // FixMinus(Re(Input()), Re(Input()))
  assign s561 = s477 - s478;
  // FixMinus(Im(Input()), Im(Input()))
  assign s564 = s483 - s484;
  // FixMinus(Re(Input()), Re(Input()))
  assign s565 = s493 - s494;
  // Re(Input())
  assign s585 = s610[15:0];
  // Re(Input())
  assign s586 = s611[15:0];
  // Im(Input())
  assign s606 = i3[31:16];
  // Im(Input())
  assign s607 = i11[31:16];
  // Re(Input())
  assign s612 = i7[15:0];
  // Re(Input())
  assign s613 = i15[15:0];
  // FixTimes(FixMinus(Re(Input()), Re(Input())), 0.7071067811865476)
  assign s614 = s619[29:14];
  // FixTimes(FixMinus(FixMinus(Im(S3), Im(S11)), FixMinus(Re(S7), Re(S15))), -0.7071067811865475)
  assign s615 = s620[29:14];
  // FixTimes(FixMinus(Re(Input()), Re(Input())), -0.7071067811865475)
  assign s616 = s621[29:14];
  // FixTimes(FixMinus(FixMinus(Im(S3), Im(S11)), FixMinus(Re(S7), Re(S15))), 0.7071067811865476)
  assign s617 = s622[29:14];
  // FixTimes(FixPlus(FixMinus(Im(S3), Im(S11)), FixMinus(Re(S7), Re(S15))), -0.7071067811865475)
  assign s618 = s623[29:14];
  assign s619 = $signed(s624) * $signed(16'd11585);
  assign s620 = $signed(s625) * $signed(16'd53951);
  assign s621 = $signed(s624) * $signed(16'd53951);
  assign s622 = $signed(s625) * $signed(16'd11585);
  assign s623 = $signed(s626) * $signed(16'd53951);
  // FixMinus(Re(Input()), Re(Input()))
  assign s627 = s585 - s586;
  // FixMinus(FixMinus(Im(Input()), Im(Input())), FixMinus(Re(Input()), Re(Input())))
  assign s628 = s630 - s631;
  // FixPlus(FixMinus(Im(Input()), Im(Input())), FixMinus(Re(Input()), Re(Input())))
  assign s629 = s630 + s631;
  // FixMinus(Im(Input()), Im(Input()))
  assign s632 = s606 - s607;
  // FixMinus(Re(Input()), Re(Input()))
  assign s633 = s612 - s613;
  always @(posedge clk)
    begin
      s17 <= s48;
      s18 <= s49;
      s19 <= s50;
      s20 <= s51;
      s21 <= s52;
      s22 <= s53;
      s23 <= s54;
      s24 <= s55;
      s25 <= s56;
      s26 <= s57;
      s27 <= s58;
      s28 <= s59;
      s29 <= s60;
      s30 <= s61;
      s31 <= s62;
      s32 <= s63;
      s33 <= s64;
      s34 <= s65;
      s35 <= s66;
      s36 <= s67;
      s37 <= s68;
      s38 <= s69;
      s39 <= s70;
      s40 <= s71;
      s41 <= s72;
      s42 <= s73;
      s43 <= s74;
      s44 <= s75;
      s45 <= s76;
      s46 <= s77;
      s47 <= s78;
      s79 <= s110;
      s80 <= s111;
      s81 <= s112;
      s82 <= s113;
      s83 <= s114;
      s84 <= s115;
      s85 <= s116;
      s86 <= s117;
      s87 <= s118;
      s88 <= s119;
      s89 <= s120;
      s90 <= s121;
      s91 <= s122;
      s92 <= s123;
      s93 <= s124;
      s94 <= s125;
      s95 <= s126;
      s96 <= s127;
      s97 <= s128;
      s98 <= s129;
      s99 <= s130;
      s100 <= s131;
      s101 <= s132;
      s102 <= s133;
      s103 <= s134;
      s104 <= s135;
      s105 <= s136;
      s106 <= s137;
      s107 <= s138;
      s108 <= s139;
      s109 <= s140;
      s128 <= s170;
      s129 <= s171;
      s141 <= s181;
      s142 <= s182;
      s143 <= s183;
      s144 <= s184;
      s145 <= s185;
      s146 <= s186;
      s147 <= s187;
      s148 <= s188;
      s149 <= s189;
      s150 <= s190;
      s151 <= s191;
      s152 <= s192;
      s153 <= s193;
      s154 <= s194;
      s155 <= s195;
      s156 <= s196;
      s157 <= s197;
      s158 <= s198;
      s159 <= s199;
      s160 <= s200;
      s161 <= s201;
      s162 <= s202;
      s163 <= s203;
      s164 <= s204;
      s165 <= s205;
      s166 <= s206;
      s167 <= s207;
      s168 <= s208;
      s169 <= s209;
      s172 <= s212;
      s173 <= s213;
      s174 <= s214;
      s175 <= s215;
      s176 <= s216;
      s177 <= s217;
      s178 <= s218;
      s179 <= s219;
      s180 <= s220;
      s189 <= s237;
      s190 <= s238;
      s193 <= s243;
      s194 <= s244;
      s197 <= s245;
      s198 <= s246;
      s199 <= s247;
      s200 <= s248;
      s201 <= s249;
      s202 <= s250;
      s205 <= s252;
      s206 <= s253;
      s208 <= s254;
      s209 <= s255;
      s210 <= s256;
      s211 <= s257;
      s212 <= s258;
      s213 <= s259;
      s214 <= s260;
      s215 <= s261;
      s216 <= s262;
      s217 <= s263;
      s218 <= s264;
      s219 <= s265;
      s220 <= s266;
      s221 <= s267;
      s222 <= s268;
      s223 <= s269;
      s224 <= s270;
      s225 <= s271;
      s226 <= s272;
      s227 <= s273;
      s228 <= s274;
      s229 <= s275;
      s230 <= s276;
      s231 <= s277;
      s232 <= s278;
      s233 <= s279;
      s234 <= s280;
      s235 <= s281;
      s236 <= s282;
      s237 <= s283;
      s238 <= s284;
      s239 <= s285;
      s240 <= s286;
      s241 <= s287;
      s242 <= s288;
      s243 <= s289;
      s244 <= s290;
      s245 <= s291;
      s246 <= s292;
      s249 <= s295;
      s250 <= s296;
      s251 <= s297;
      s252 <= s298;
      s253 <= s299;
      s254 <= s300;
      s255 <= s301;
      s258 <= s306;
      s259 <= s307;
      s260 <= s308;
      s261 <= s309;
      s262 <= s310;
      s263 <= s311;
      s264 <= s312;
      s265 <= s313;
      s266 <= s314;
      s271 <= s323;
      s272 <= s324;
      s275 <= s329;
      s276 <= s330;
      s277 <= s331;
      s278 <= s332;
      s281 <= s333;
      s282 <= s334;
      s287 <= s339;
      s288 <= s340;
      s297 <= s349;
      s302 <= s354;
      s303 <= s355;
      s304 <= s356;
      s305 <= s357;
      s319 <= s367;
      s320 <= s368;
      s323 <= s371;
      s324 <= s372;
      s325 <= s373;
      s326 <= s374;
      s329 <= s377;
      s330 <= s378;
      s331 <= s379;
      s332 <= s380;
      s333 <= s381;
      s334 <= s382;
      s337 <= s385;
      s338 <= s386;
      s339 <= s387;
      s340 <= s388;
      s345 <= s391;
      s346 <= s392;
      s349 <= s393;
      s354 <= s396;
      s355 <= s397;
      s356 <= s398;
      s357 <= s399;
      s367 <= s405;
      s368 <= s406;
      s369 <= s407;
      s370 <= s408;
      s371 <= s409;
      s372 <= s410;
      s373 <= s411;
      s374 <= s412;
      s375 <= s413;
      s376 <= s414;
      s377 <= s415;
      s378 <= s416;
      s379 <= s417;
      s380 <= s418;
      s383 <= s421;
      s384 <= s422;
      s385 <= s423;
      s386 <= s424;
      s389 <= s427;
      s390 <= s428;
      s391 <= s429;
      s392 <= s430;
      s394 <= s432;
      s395 <= s433;
      s396 <= s434;
      s397 <= s435;
      s398 <= s436;
      s399 <= s437;
      s400 <= s438;
      s401 <= s439;
      s402 <= s440;
      s403 <= s441;
      s404 <= s442;
      s405 <= s443;
      s406 <= s444;
      s407 <= s445;
      s408 <= s446;
      s409 <= s447;
      s410 <= s448;
      s411 <= s449;
      s412 <= s450;
      s413 <= s451;
      s414 <= s452;
      s417 <= s457;
      s418 <= s458;
      s423 <= s465;
      s424 <= s466;
      s429 <= s469;
      s430 <= s470;
      s436 <= s477;
      s437 <= s478;
      s443 <= s479;
      s444 <= s480;
      s445 <= s481;
      s446 <= s482;
      s449 <= s487;
      s450 <= s488;
      s451 <= s489;
      s452 <= s490;
      s455 <= s493;
      s456 <= s494;
      s459 <= s499;
      s460 <= s500;
      s461 <= s501;
      s462 <= s502;
      s463 <= s503;
      s464 <= s504;
      s465 <= s505;
      s466 <= s506;
      s467 <= s507;
      s468 <= s508;
      s469 <= s509;
      s470 <= s510;
      s471 <= s511;
      s472 <= s512;
      s473 <= s513;
      s474 <= s514;
      s475 <= s515;
      s476 <= s516;
      s481 <= s517;
      s482 <= s518;
      s487 <= s523;
      s488 <= s524;
      s489 <= s525;
      s490 <= s526;
      s491 <= s519;
      s492 <= s520;
      s495 <= s527;
      s496 <= s528;
      s497 <= s529;
      s498 <= s530;
      s505 <= s539;
      s506 <= s540;
      s509 <= s541;
      s510 <= s542;
      s515 <= s544;
      s516 <= s545;
      s517 <= s546;
      s518 <= s547;
      s519 <= s548;
      s520 <= s549;
      s521 <= s550;
      s522 <= s551;
      s523 <= s552;
      s524 <= s553;
      s525 <= s554;
      s526 <= s555;
      s527 <= s556;
      s528 <= s557;
      s529 <= s558;
      s530 <= s559;
      s531 <= s560;
      s532 <= s561;
      s533 <= s562;
      s534 <= s563;
      s535 <= s564;
      s536 <= s565;
      s537 <= s566;
      s538 <= s567;
      s539 <= s568;
      s540 <= s569;
      s541 <= s570;
      s542 <= s571;
      s543 <= s572;
      s544 <= s573;
      s545 <= s574;
      s546 <= s575;
      s547 <= s576;
      s548 <= s577;
      s549 <= s578;
      s550 <= s579;
      s551 <= s580;
      s552 <= s581;
      s553 <= s582;
      s554 <= s583;
      s555 <= s584;
      s556 <= s585;
      s557 <= s586;
      s558 <= s587;
      s559 <= s588;
      s562 <= s589;
      s563 <= s590;
      s566 <= s591;
      s567 <= s592;
      s568 <= s593;
      s569 <= s594;
      s570 <= s595;
      s571 <= s596;
      s572 <= s597;
      s573 <= s598;
      s574 <= s599;
      s575 <= s600;
      s576 <= s601;
      s577 <= s602;
      s578 <= s603;
      s579 <= s604;
      s580 <= s605;
      s581 <= s606;
      s582 <= s607;
      s583 <= s608;
      s584 <= s609;
      s587 <= s612;
      s588 <= s613;
      s589 <= s614;
      s590 <= s615;
      s591 <= s616;
      s592 <= s617;
      s593 <= i0;
      s594 <= i8;
      s595 <= i4;
      s596 <= i12;
      s597 <= s618;
      s598 <= i2;
      s599 <= i10;
      s600 <= i6;
      s601 <= i14;
      s602 <= i1;
      s603 <= i9;
      s604 <= i5;
      s605 <= i13;
      s608 <= i7;
      s609 <= i15;
      s610 <= i3;
      s611 <= i11;
      s624 <= s627;
      s625 <= s628;
      s626 <= s629;
      s630 <= s632;
      s631 <= s633;
    end
endmodule
